magic
tech gf180mcuD
magscale 1 10
timestamp 1712602796
<< metal1 >>
rect 346770 325054 346782 325106
rect 346834 325103 346846 325106
rect 347106 325103 347118 325106
rect 346834 325057 347118 325103
rect 346834 325054 346846 325057
rect 347106 325054 347118 325057
rect 347170 325054 347182 325106
rect 352370 267150 352382 267202
rect 352434 267199 352446 267202
rect 354274 267199 354286 267202
rect 352434 267153 354286 267199
rect 352434 267150 352446 267153
rect 354274 267150 354286 267153
rect 354338 267150 354350 267202
rect 338706 241502 338718 241554
rect 338770 241551 338782 241554
rect 340386 241551 340398 241554
rect 338770 241505 340398 241551
rect 338770 241502 338782 241505
rect 340386 241502 340398 241505
rect 340450 241502 340462 241554
rect 300178 160638 300190 160690
rect 300242 160687 300254 160690
rect 301298 160687 301310 160690
rect 300242 160641 301310 160687
rect 300242 160638 300254 160641
rect 301298 160638 301310 160641
rect 301362 160638 301374 160690
<< via1 >>
rect 346782 325054 346834 325106
rect 347118 325054 347170 325106
rect 352382 267150 352434 267202
rect 354286 267150 354338 267202
rect 338718 241502 338770 241554
rect 340398 241502 340450 241554
rect 300190 160638 300242 160690
rect 301310 160638 301362 160690
<< metal2 >>
rect 11032 595672 11256 597000
rect 11004 595560 11256 595672
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 33096 595560 33348 595672
rect 55160 595560 55412 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 99288 595560 99540 595672
rect 121352 595560 121604 595672
rect 4172 502516 4228 502526
rect 4172 469588 4228 502460
rect 4172 469522 4228 469532
rect 4508 388948 4564 388958
rect 4508 333396 4564 388892
rect 4508 333330 4564 333340
rect 11004 301588 11060 595560
rect 33292 590548 33348 595560
rect 55356 590660 55412 595560
rect 55356 590594 55412 590604
rect 33292 590482 33348 590492
rect 77308 583828 77364 595560
rect 99484 590772 99540 595560
rect 121548 590884 121604 595560
rect 121548 590818 121604 590828
rect 143388 595560 143640 595672
rect 165452 595560 165704 595672
rect 187516 595560 187768 595672
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319900 595560 320152 595672
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 430220 595560 430472 595672
rect 452284 595560 452536 595672
rect 474348 595560 474600 595672
rect 496412 595560 496664 595672
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 518504 595560 518756 595672
rect 99484 590706 99540 590716
rect 77308 583762 77364 583772
rect 143388 582148 143444 595560
rect 153692 590772 153748 590782
rect 143388 582082 143444 582092
rect 152012 590660 152068 590670
rect 57932 573076 57988 573086
rect 56252 530740 56308 530750
rect 14252 488404 14308 488414
rect 14252 390628 14308 488348
rect 56252 390740 56308 530684
rect 57932 390964 57988 573020
rect 93212 460180 93268 460190
rect 66332 417620 66388 417630
rect 64092 417060 64148 417070
rect 64092 413896 64148 417004
rect 66332 413896 66388 417564
rect 88172 417620 88228 417630
rect 68572 417508 68628 417518
rect 68572 413896 68628 417452
rect 73052 417396 73108 417406
rect 70812 417284 70868 417294
rect 70812 413896 70868 417228
rect 73052 413896 73108 417340
rect 85036 417396 85092 417406
rect 75292 417172 75348 417182
rect 75292 413896 75348 417116
rect 79772 416948 79828 416958
rect 77532 416724 77588 416734
rect 77532 413896 77588 416668
rect 79772 413896 79828 416892
rect 82012 416836 82068 416846
rect 82012 413896 82068 416780
rect 84812 416724 84868 416734
rect 61852 413364 61908 413374
rect 61852 413298 61908 413308
rect 57932 390898 57988 390908
rect 59612 403732 59668 403742
rect 59612 390852 59668 403676
rect 59612 390786 59668 390796
rect 56252 390674 56308 390684
rect 14252 390562 14308 390572
rect 78428 388164 78484 388174
rect 40908 386484 40964 386494
rect 38444 383348 38500 383358
rect 24332 383124 24388 383134
rect 11004 301522 11060 301532
rect 14252 380212 14308 380222
rect 13244 224308 13300 224318
rect 4172 121492 4228 121502
rect 4172 50372 4228 121436
rect 4172 50306 4228 50316
rect 11564 5908 11620 5918
rect 11564 480 11620 5852
rect 11368 392 11620 480
rect 13244 480 13300 224252
rect 14252 192052 14308 380156
rect 22764 232932 22820 232942
rect 14252 191986 14308 191996
rect 18956 229348 19012 229358
rect 15372 4228 15428 4238
rect 15372 480 15428 4172
rect 17276 4228 17332 4238
rect 17276 480 17332 4172
rect 13244 392 13496 480
rect 11368 -960 11592 392
rect 13272 -960 13496 392
rect 15176 392 15428 480
rect 17080 392 17332 480
rect 18956 480 19012 229292
rect 21084 4228 21140 4238
rect 21084 480 21140 4172
rect 18956 392 19208 480
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 392 21140 480
rect 22764 480 22820 232876
rect 24332 149716 24388 383068
rect 38332 380436 38388 380446
rect 34412 379652 34468 379662
rect 34412 276724 34468 379596
rect 34412 276658 34468 276668
rect 38220 379540 38276 379550
rect 38220 238308 38276 379484
rect 38220 238242 38276 238252
rect 38332 238196 38388 380380
rect 38444 240772 38500 383292
rect 38444 240706 38500 240716
rect 38556 383236 38612 383246
rect 38556 238532 38612 383180
rect 38556 238466 38612 238476
rect 40236 292404 40292 292414
rect 38332 238130 38388 238140
rect 35196 236180 35252 236190
rect 34188 232708 34244 232718
rect 24332 149650 24388 149660
rect 24668 214228 24724 214238
rect 24668 480 24724 214172
rect 30380 212660 30436 212670
rect 27692 79156 27748 79166
rect 27692 50260 27748 79100
rect 27692 50194 27748 50204
rect 26796 4228 26852 4238
rect 26796 480 26852 4172
rect 30380 480 30436 212604
rect 32508 4228 32564 4238
rect 32508 480 32564 4172
rect 22764 392 23016 480
rect 24668 392 24920 480
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 392 26852 480
rect 26600 -960 26824 392
rect 28504 -960 28728 480
rect 30380 392 30632 480
rect 30408 -960 30632 392
rect 32312 392 32564 480
rect 34188 480 34244 232652
rect 35196 4676 35252 236124
rect 38556 232820 38612 232830
rect 37996 227780 38052 227790
rect 35196 4610 35252 4620
rect 36876 222740 36932 222750
rect 36876 4452 36932 222684
rect 36876 4386 36932 4396
rect 37996 480 38052 227724
rect 38444 217588 38500 217598
rect 38444 4116 38500 217532
rect 38556 4340 38612 232764
rect 39900 221060 39956 221070
rect 39788 212548 39844 212558
rect 39788 4564 39844 212492
rect 39788 4498 39844 4508
rect 38556 4274 38612 4284
rect 38444 4050 38500 4060
rect 39900 480 39956 221004
rect 40124 214340 40180 214350
rect 40012 212772 40068 212782
rect 40012 4900 40068 212716
rect 40124 5012 40180 214284
rect 40236 47012 40292 292348
rect 40908 255388 40964 386428
rect 69692 386148 69748 386158
rect 55580 380996 55636 381006
rect 49532 379092 49588 379102
rect 49532 319060 49588 379036
rect 55580 360920 55636 380940
rect 63196 363748 63252 363758
rect 59388 363076 59444 363086
rect 59388 360920 59444 363020
rect 63196 360920 63252 363692
rect 67004 362964 67060 362974
rect 67004 360920 67060 362908
rect 69692 362964 69748 386092
rect 74620 379428 74676 379438
rect 69692 362898 69748 362908
rect 70812 363860 70868 363870
rect 70812 360920 70868 363804
rect 74620 360920 74676 379372
rect 78428 360920 78484 388108
rect 84812 383908 84868 416668
rect 85036 384020 85092 417340
rect 86492 417172 86548 417182
rect 85260 417060 85316 417070
rect 85260 397572 85316 417004
rect 85260 397506 85316 397516
rect 86492 392308 86548 417116
rect 86716 416948 86772 416958
rect 86716 397348 86772 416892
rect 87276 409108 87332 409118
rect 87276 407428 87332 409052
rect 87276 407362 87332 407372
rect 88172 397572 88228 417564
rect 88172 397506 88228 397516
rect 91532 417508 91588 417518
rect 86716 397282 86772 397292
rect 91532 392420 91588 417452
rect 93212 409668 93268 460124
rect 93212 409602 93268 409612
rect 152012 409556 152068 590604
rect 152012 409490 152068 409500
rect 153692 395668 153748 590716
rect 153692 395602 153748 395612
rect 155372 590548 155428 590558
rect 155372 392644 155428 590492
rect 160412 446068 160468 446078
rect 160412 399028 160468 446012
rect 160412 398962 160468 398972
rect 165452 397908 165508 595560
rect 168812 590884 168868 590894
rect 168812 409444 168868 590828
rect 186396 590548 186452 590558
rect 173852 583828 173908 583838
rect 168812 409378 168868 409388
rect 170492 582148 170548 582158
rect 168028 407428 168084 407438
rect 168028 406644 168084 407372
rect 168084 406588 168196 406644
rect 168028 406578 168084 406588
rect 165452 397842 165508 397852
rect 168028 405748 168084 405758
rect 168028 404964 168084 405692
rect 155372 392578 155428 392588
rect 91532 392354 91588 392364
rect 86492 392242 86548 392252
rect 85036 383954 85092 383964
rect 85708 391636 85764 391646
rect 84812 383842 84868 383852
rect 82236 379876 82292 379886
rect 82236 360920 82292 379820
rect 85708 363076 85764 391580
rect 103292 386932 103348 386942
rect 96572 386820 96628 386830
rect 94892 386708 94948 386718
rect 93660 380100 93716 380110
rect 91532 379988 91588 379998
rect 85708 361284 85764 363020
rect 85708 361218 85764 361228
rect 86044 363972 86100 363982
rect 86044 360920 86100 363916
rect 89852 362964 89908 362974
rect 89852 360920 89908 362908
rect 91532 362964 91588 379932
rect 91532 362898 91588 362908
rect 93660 360920 93716 380044
rect 49532 318994 49588 319004
rect 51660 360220 51800 360276
rect 46284 293188 46340 293198
rect 46284 292404 46340 293132
rect 51660 293188 51716 360220
rect 51660 293122 51716 293132
rect 59052 293972 59108 293982
rect 46284 290920 46340 292348
rect 59052 290920 59108 293916
rect 87276 293188 87332 293198
rect 71820 292404 71876 292414
rect 71820 290920 71876 292348
rect 84588 292404 84644 292414
rect 84588 290920 84644 292348
rect 87276 290388 87332 293132
rect 87276 290322 87332 290332
rect 40684 255332 40964 255388
rect 40684 238420 40740 255332
rect 93212 250628 93268 250638
rect 40684 238354 40740 238364
rect 40908 248500 40964 248510
rect 40908 235172 40964 248444
rect 90188 241220 90244 241230
rect 41132 240772 41188 240782
rect 41132 240706 41188 240716
rect 66220 240772 66276 240782
rect 66220 240706 66276 240716
rect 71596 240772 71652 240782
rect 71596 240706 71652 240716
rect 80556 240660 80612 240670
rect 80556 240594 80612 240604
rect 90188 240660 90244 241164
rect 90188 240594 90244 240604
rect 60844 240548 60900 240558
rect 60844 240482 60900 240492
rect 57260 240436 57316 240446
rect 57260 240370 57316 240380
rect 53676 240324 53732 240334
rect 53676 240258 53732 240268
rect 46508 240212 46564 240222
rect 46508 240146 46564 240156
rect 85932 240212 85988 240222
rect 85932 240146 85988 240156
rect 55468 240100 55524 240110
rect 42924 238532 42980 240072
rect 42924 238466 42980 238476
rect 44716 238308 44772 240072
rect 44716 238242 44772 238252
rect 48300 238196 48356 240072
rect 48300 238130 48356 238140
rect 50092 237972 50148 240072
rect 51884 238420 51940 240072
rect 55468 240034 55524 240044
rect 51884 238354 51940 238364
rect 50092 237906 50148 237916
rect 41020 235172 41076 235182
rect 40908 235116 41020 235172
rect 41020 235106 41076 235116
rect 41020 234500 41076 234510
rect 40908 227892 40964 227902
rect 40684 224532 40740 224542
rect 40684 48244 40740 224476
rect 40684 48178 40740 48188
rect 40796 224420 40852 224430
rect 40796 48020 40852 224364
rect 40908 50148 40964 227836
rect 40908 50082 40964 50092
rect 41020 49588 41076 234444
rect 41132 234388 41188 234398
rect 41132 49700 41188 234332
rect 59052 233492 59108 240072
rect 62636 238532 62692 240072
rect 62636 238466 62692 238476
rect 64428 238532 64484 240072
rect 64428 238466 64484 238476
rect 68012 237636 68068 240072
rect 69804 238196 69860 240072
rect 69804 238130 69860 238140
rect 73388 237972 73444 240072
rect 73388 237906 73444 237916
rect 75180 237860 75236 240072
rect 76972 238084 77028 240072
rect 76972 238018 77028 238028
rect 75180 237794 75236 237804
rect 78764 237748 78820 240072
rect 82348 239876 82404 240072
rect 82348 239810 82404 239820
rect 84140 238420 84196 240072
rect 87724 238532 87780 240072
rect 87724 238466 87780 238476
rect 84140 238354 84196 238364
rect 89516 238308 89572 240072
rect 89516 238242 89572 238252
rect 78764 237682 78820 237692
rect 68012 237570 68068 237580
rect 59052 233426 59108 233436
rect 93212 229460 93268 250572
rect 93212 229394 93268 229404
rect 93324 246372 93380 246382
rect 93324 227668 93380 246316
rect 93436 242004 93492 242014
rect 93436 231028 93492 241948
rect 94892 238084 94948 386652
rect 95116 386596 95172 386606
rect 95116 238308 95172 386540
rect 95340 385476 95396 385486
rect 95340 238532 95396 385420
rect 95340 238466 95396 238476
rect 95564 383460 95620 383470
rect 95116 238242 95172 238252
rect 95564 238196 95620 383404
rect 95564 238130 95620 238140
rect 94892 238018 94948 238028
rect 96572 237748 96628 386764
rect 96572 237682 96628 237692
rect 96796 385140 96852 385150
rect 96796 237636 96852 385084
rect 99932 385028 99988 385038
rect 99932 238420 99988 384972
rect 99932 238354 99988 238364
rect 103292 237972 103348 386876
rect 103292 237906 103348 237916
rect 104972 385364 105028 385374
rect 104972 237860 105028 385308
rect 111692 382676 111748 382686
rect 108332 321748 108388 321758
rect 106652 320068 106708 320078
rect 106652 263396 106708 320012
rect 108332 267652 108388 321692
rect 108332 267586 108388 267596
rect 106652 263330 106708 263340
rect 111692 241108 111748 382620
rect 167132 382116 167188 382126
rect 118412 381892 118468 381902
rect 111692 241042 111748 241052
rect 113372 381780 113428 381790
rect 113372 239988 113428 381724
rect 116732 381556 116788 381566
rect 116732 241220 116788 381500
rect 116732 241154 116788 241164
rect 118412 240772 118468 381836
rect 118412 240706 118468 240716
rect 120092 381668 120148 381678
rect 113372 239922 113428 239932
rect 120092 239876 120148 381612
rect 121772 380324 121828 380334
rect 120204 378980 120260 378990
rect 120204 361396 120260 378924
rect 121772 363972 121828 380268
rect 121772 363906 121828 363916
rect 120204 361330 120260 361340
rect 152796 321860 152852 321870
rect 144284 290388 144340 290398
rect 144284 289828 144340 290332
rect 144284 285880 144340 289772
rect 152796 285880 152852 321804
rect 161308 294868 161364 294878
rect 161308 285880 161364 294812
rect 167132 240100 167188 382060
rect 167244 356356 167300 356366
rect 167244 321860 167300 356300
rect 168028 342916 168084 404908
rect 168028 342850 168084 342860
rect 168140 346276 168196 406588
rect 167244 321794 167300 321804
rect 168140 320068 168196 346220
rect 168140 320002 168196 320012
rect 168812 382004 168868 382014
rect 167132 240034 167188 240044
rect 167244 318276 167300 318286
rect 120092 239810 120148 239820
rect 104972 237794 105028 237804
rect 96796 237570 96852 237580
rect 93436 230962 93492 230972
rect 93324 227602 93380 227612
rect 154924 217700 154980 217710
rect 154924 209944 154980 217644
rect 167244 217700 167300 318220
rect 168812 240212 168868 381948
rect 169148 289940 169204 289950
rect 169036 286468 169092 286478
rect 168924 284788 168980 284798
rect 168924 273924 168980 284732
rect 169036 275940 169092 286412
rect 169148 284004 169204 289884
rect 169148 283938 169204 283948
rect 169260 288148 169316 288158
rect 169260 279972 169316 288092
rect 169260 279906 169316 279916
rect 169372 286580 169428 286590
rect 169372 277956 169428 286524
rect 169372 277890 169428 277900
rect 169036 275874 169092 275884
rect 170492 274596 170548 582092
rect 172172 397796 172228 397806
rect 170492 274530 170548 274540
rect 170604 382228 170660 382238
rect 168924 273858 168980 273868
rect 170604 240324 170660 382172
rect 172172 322756 172228 397740
rect 172172 322690 172228 322700
rect 172956 331716 173012 331726
rect 170604 240258 170660 240268
rect 168812 240146 168868 240156
rect 172956 224868 173012 331660
rect 173852 275716 173908 583772
rect 183036 578788 183092 578798
rect 180572 417284 180628 417294
rect 177212 416836 177268 416846
rect 177212 397684 177268 416780
rect 177212 397618 177268 397628
rect 175532 395780 175588 395790
rect 173964 392868 174020 392878
rect 173964 330932 174020 392812
rect 175532 332836 175588 395724
rect 177324 392756 177380 392766
rect 177212 357476 177268 357486
rect 176204 355236 176260 355246
rect 175532 332770 175588 332780
rect 176092 347396 176148 347406
rect 173964 330866 174020 330876
rect 173852 275650 173908 275660
rect 174412 330596 174468 330606
rect 174412 230020 174468 330540
rect 175980 328356 176036 328366
rect 174636 326116 174692 326126
rect 174412 229954 174468 229964
rect 174524 324996 174580 325006
rect 172956 224802 173012 224812
rect 174524 222964 174580 324940
rect 174524 222898 174580 222908
rect 174636 221284 174692 326060
rect 175532 301588 175588 301598
rect 175532 276836 175588 301532
rect 175532 276770 175588 276780
rect 175644 283108 175700 283118
rect 175644 272132 175700 283052
rect 175644 272066 175700 272076
rect 175980 233268 176036 328300
rect 175980 233202 176036 233212
rect 176092 231252 176148 347340
rect 176092 231186 176148 231196
rect 176204 231140 176260 355180
rect 176204 231074 176260 231084
rect 176316 349524 176372 349534
rect 176316 224644 176372 349468
rect 177212 294868 177268 357420
rect 177324 336868 177380 392700
rect 180572 384132 180628 417228
rect 180572 384066 180628 384076
rect 181356 352996 181412 353006
rect 177884 351876 177940 351886
rect 177324 336802 177380 336812
rect 177772 345156 177828 345166
rect 177212 294802 177268 294812
rect 177772 228116 177828 345100
rect 177884 233044 177940 351820
rect 179452 348516 179508 348526
rect 177884 232978 177940 232988
rect 177996 346276 178052 346286
rect 177772 228050 177828 228060
rect 176316 224578 176372 224588
rect 174636 221218 174692 221228
rect 177996 221172 178052 346220
rect 179340 340676 179396 340686
rect 179228 327236 179284 327246
rect 179228 234836 179284 327180
rect 179228 234770 179284 234780
rect 179340 231364 179396 340620
rect 179452 234724 179508 348460
rect 179676 344036 179732 344046
rect 179452 234658 179508 234668
rect 179564 339556 179620 339566
rect 179340 231298 179396 231308
rect 179564 224756 179620 339500
rect 179564 224690 179620 224700
rect 179676 222628 179732 343980
rect 181132 342916 181188 342926
rect 181020 335076 181076 335086
rect 181020 228228 181076 335020
rect 181132 229796 181188 342860
rect 181132 229730 181188 229740
rect 181244 338436 181300 338446
rect 181020 228162 181076 228172
rect 181244 222852 181300 338380
rect 181356 229684 181412 352940
rect 182700 341796 182756 341806
rect 181356 229618 181412 229628
rect 182588 323876 182644 323886
rect 181244 222786 181300 222796
rect 179676 222562 179732 222572
rect 177996 221106 178052 221116
rect 182588 219604 182644 323820
rect 182700 233156 182756 341740
rect 182924 336196 182980 336206
rect 182700 233090 182756 233100
rect 182812 329476 182868 329486
rect 182588 219538 182644 219548
rect 167244 217634 167300 217644
rect 182812 216020 182868 329420
rect 182924 219380 182980 336140
rect 183036 273476 183092 578732
rect 184716 575540 184772 575550
rect 184604 354116 184660 354126
rect 183036 273410 183092 273420
rect 184492 337316 184548 337326
rect 182924 219314 182980 219324
rect 184492 217700 184548 337260
rect 184604 228004 184660 354060
rect 184716 267876 184772 575484
rect 186284 566132 186340 566142
rect 186172 543620 186228 543630
rect 186060 529284 186116 529294
rect 185612 412020 185668 412030
rect 185612 385588 185668 411964
rect 186060 389060 186116 529228
rect 186060 388994 186116 389004
rect 186172 387268 186228 543564
rect 186284 407988 186340 566076
rect 186284 407922 186340 407932
rect 186396 404068 186452 590492
rect 187516 566132 187572 595560
rect 189756 588868 189812 588878
rect 189644 577108 189700 577118
rect 187516 566066 187572 566076
rect 189308 575428 189364 575438
rect 187964 557956 188020 557966
rect 186396 404002 186452 404012
rect 187292 507780 187348 507790
rect 186172 387202 186228 387212
rect 185612 385522 185668 385532
rect 185724 383572 185780 383582
rect 184716 267810 184772 267820
rect 185612 382340 185668 382350
rect 185612 240436 185668 382284
rect 185724 363860 185780 383516
rect 185724 363794 185780 363804
rect 185948 380548 186004 380558
rect 185948 363748 186004 380492
rect 185948 363682 186004 363692
rect 186396 332836 186452 332846
rect 185612 240370 185668 240380
rect 186284 322756 186340 322766
rect 186284 234948 186340 322700
rect 186284 234882 186340 234892
rect 184604 227938 184660 227948
rect 186396 217812 186452 332780
rect 186508 296548 186564 296558
rect 186508 284788 186564 296492
rect 187292 289940 187348 507724
rect 187292 289874 187348 289884
rect 187404 493444 187460 493454
rect 187404 288148 187460 493388
rect 187404 288082 187460 288092
rect 187516 486276 187572 486286
rect 186508 284722 186564 284732
rect 187068 287364 187124 287374
rect 187068 282100 187124 287308
rect 187516 286580 187572 486220
rect 187740 479108 187796 479118
rect 187516 286514 187572 286524
rect 187628 464772 187684 464782
rect 187628 283108 187684 464716
rect 187740 286468 187796 479052
rect 187740 286402 187796 286412
rect 187852 457604 187908 457614
rect 187628 283042 187684 283052
rect 187068 282034 187124 282044
rect 187852 280644 187908 457548
rect 187964 409332 188020 557900
rect 187964 409266 188020 409276
rect 188076 414596 188132 414606
rect 188076 289828 188132 414540
rect 189308 407428 189364 575372
rect 189532 572068 189588 572078
rect 189308 407362 189364 407372
rect 189420 570388 189476 570398
rect 189308 350756 189364 350766
rect 189196 333956 189252 333966
rect 188076 289044 188132 289772
rect 189084 321636 189140 321646
rect 188076 288978 188132 288988
rect 188972 289044 189028 289054
rect 188076 280644 188132 280654
rect 187852 280588 188076 280644
rect 188076 280578 188132 280588
rect 188076 252196 188132 252206
rect 187964 251076 188020 251086
rect 187964 218036 188020 251020
rect 187964 217970 188020 217980
rect 186396 217746 186452 217756
rect 184492 217634 184548 217644
rect 182812 215954 182868 215964
rect 188076 214788 188132 252140
rect 188972 240212 189028 288988
rect 188972 240146 189028 240156
rect 189084 217924 189140 321580
rect 189196 219492 189252 333900
rect 189308 229908 189364 350700
rect 189420 272356 189476 570332
rect 189420 272290 189476 272300
rect 189532 268996 189588 572012
rect 189644 271236 189700 577052
rect 189644 271170 189700 271180
rect 189756 270116 189812 588812
rect 209580 578788 209636 595560
rect 231644 591332 231700 595560
rect 231644 591266 231700 591276
rect 209580 578722 209636 578732
rect 253708 568708 253764 595560
rect 275772 570388 275828 595560
rect 297836 591220 297892 595560
rect 297836 591154 297892 591164
rect 319900 591108 319956 595560
rect 319900 591042 319956 591052
rect 341964 577108 342020 595560
rect 364028 590996 364084 595560
rect 364028 590930 364084 590940
rect 386092 590884 386148 595560
rect 386092 590818 386148 590828
rect 408268 588868 408324 595560
rect 430220 590772 430276 595560
rect 430220 590706 430276 590716
rect 452284 590212 452340 595560
rect 452284 590146 452340 590156
rect 408268 588802 408324 588812
rect 341964 577042 342020 577052
rect 474348 572068 474404 595560
rect 496412 590660 496468 595560
rect 496412 590594 496468 590604
rect 518700 590660 518756 595560
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 518700 590594 518756 590604
rect 529788 590660 529844 590670
rect 474348 572002 474404 572012
rect 275772 570322 275828 570332
rect 253708 568642 253764 568652
rect 529340 526820 529396 526830
rect 511868 410116 511924 410126
rect 192444 392868 192500 410088
rect 197596 395780 197652 410088
rect 197596 395714 197652 395724
rect 192444 392802 192500 392812
rect 202748 392756 202804 410088
rect 207900 408548 207956 410088
rect 207900 406756 207956 408492
rect 207900 406690 207956 406700
rect 210364 407428 210420 407438
rect 202748 392690 202804 392700
rect 207004 403284 207060 403294
rect 205100 389172 205156 389182
rect 202748 382564 202804 382574
rect 201404 382452 201460 382462
rect 201404 379988 201460 382396
rect 202748 379988 202804 382508
rect 204204 382564 204260 382574
rect 203084 382452 203140 382462
rect 203084 379988 203140 382396
rect 204204 379988 204260 382508
rect 204876 382452 204932 382462
rect 204876 379988 204932 382396
rect 205100 379988 205156 389116
rect 207004 384748 207060 403228
rect 208348 402388 208404 402398
rect 208348 396508 208404 402332
rect 208348 396452 208516 396508
rect 206892 384692 207060 384748
rect 206108 382564 206164 382574
rect 206108 379988 206164 382508
rect 206444 382452 206500 382462
rect 206444 379988 206500 382396
rect 200984 379932 201460 379988
rect 202328 379932 202804 379988
rect 203000 379932 203140 379988
rect 203672 379932 204260 379988
rect 204344 379932 204932 379988
rect 205016 379932 205156 379988
rect 205688 379932 206164 379988
rect 206360 379932 206500 379988
rect 206892 379988 206948 384692
rect 208124 382452 208180 382462
rect 208124 379988 208180 382396
rect 208460 379988 208516 396452
rect 210364 384748 210420 407372
rect 213052 406084 213108 410088
rect 213052 406018 213108 406028
rect 218204 406644 218260 410088
rect 218204 405860 218260 406588
rect 218204 405794 218260 405804
rect 211036 404068 211092 404078
rect 211036 384748 211092 404012
rect 211708 399140 211764 399150
rect 211708 396508 211764 399084
rect 219100 399028 219156 399038
rect 215068 397908 215124 397918
rect 215068 396508 215124 397852
rect 211708 396452 211876 396508
rect 215068 396452 215236 396508
rect 211596 394548 211652 394558
rect 211596 391076 211652 394492
rect 211596 391010 211652 391020
rect 210252 384692 210420 384748
rect 210924 384692 211092 384748
rect 209468 382564 209524 382574
rect 209468 379988 209524 382508
rect 209804 382452 209860 382462
rect 209804 379988 209860 382396
rect 206892 379932 207032 379988
rect 207704 379932 208180 379988
rect 208376 379932 208516 379988
rect 209048 379932 209524 379988
rect 209720 379932 209860 379988
rect 210252 379988 210308 384692
rect 210924 379988 210980 384692
rect 211820 379988 211876 396452
rect 213612 395892 213668 395902
rect 210252 379932 210392 379988
rect 210924 379932 211064 379988
rect 211736 379932 211876 379988
rect 212268 392868 212324 392878
rect 212268 379988 212324 392812
rect 212940 392756 212996 392766
rect 212940 379988 212996 392700
rect 213612 379988 213668 395836
rect 214284 395780 214340 395790
rect 214284 379988 214340 395724
rect 215180 379988 215236 396452
rect 212268 379932 212408 379988
rect 212940 379932 213080 379988
rect 213612 379932 213752 379988
rect 214284 379932 214424 379988
rect 215096 379932 215236 379988
rect 215628 395668 215684 395678
rect 215628 379988 215684 395612
rect 216300 392644 216356 392654
rect 216300 379988 216356 392588
rect 216972 390964 217028 390974
rect 216972 379988 217028 390908
rect 217644 390740 217700 390750
rect 217644 379988 217700 390684
rect 218540 390628 218596 390638
rect 218540 379988 218596 390572
rect 219100 384748 219156 398972
rect 223356 398132 223412 410088
rect 228508 409892 228564 410088
rect 228508 406644 228564 409836
rect 233660 407428 233716 410088
rect 238812 407540 238868 410088
rect 243964 407652 244020 410088
rect 243964 407586 244020 407596
rect 238812 407474 238868 407484
rect 233660 407362 233716 407372
rect 249116 407092 249172 410088
rect 254268 407204 254324 410088
rect 254268 407138 254324 407148
rect 259420 408100 259476 410088
rect 249116 407026 249172 407036
rect 228508 406578 228564 406588
rect 259420 406644 259476 408044
rect 263788 410060 264600 410116
rect 268940 410060 269752 410116
rect 274652 410060 274904 410116
rect 280056 410060 280532 410116
rect 263788 407764 263844 410060
rect 259420 406578 259476 406588
rect 260428 406644 260484 406654
rect 252700 406420 252756 406430
rect 252028 405860 252084 405870
rect 251356 405748 251412 405758
rect 250012 400708 250068 400718
rect 223356 398066 223412 398076
rect 248668 399028 248724 399038
rect 248668 396508 248724 398972
rect 248668 396452 248836 396508
rect 215628 379932 215768 379988
rect 216300 379932 216440 379988
rect 216972 379932 217112 379988
rect 217644 379932 217784 379988
rect 218456 379932 218596 379988
rect 218988 384692 219156 384748
rect 219660 390852 219716 390862
rect 218988 379988 219044 384692
rect 219660 379988 219716 390796
rect 240828 386932 240884 386942
rect 232764 386484 232820 386494
rect 228732 383348 228788 383358
rect 223468 383124 223524 383134
rect 222572 380212 222628 380222
rect 222628 380156 222740 380212
rect 222572 380146 222628 380156
rect 222684 379988 222740 380156
rect 223468 379988 223524 383068
rect 226492 382116 226548 382126
rect 226492 381444 226548 382060
rect 226492 381378 226548 381388
rect 226716 382116 226772 382126
rect 226716 379988 226772 382060
rect 218988 379932 219128 379988
rect 219660 379932 219800 379988
rect 222684 379932 223160 379988
rect 223468 379932 223832 379988
rect 226520 379932 226772 379988
rect 228732 379988 228788 383292
rect 229292 383236 229348 383246
rect 229348 383180 229460 383236
rect 229292 383170 229348 383180
rect 229404 379988 229460 383180
rect 230636 381444 230692 381454
rect 230692 381388 230804 381444
rect 230636 381378 230692 381388
rect 230748 379988 230804 381388
rect 231868 380436 231924 380446
rect 231924 380380 232036 380436
rect 231868 380370 231924 380380
rect 231980 379988 232036 380380
rect 228732 379932 229208 379988
rect 229404 379932 229880 379988
rect 230748 379932 231224 379988
rect 231896 379932 232036 379988
rect 232764 379988 232820 386428
rect 237468 385252 237524 385262
rect 235228 382340 235284 382350
rect 235284 382284 235396 382340
rect 235228 382274 235284 382284
rect 233548 382228 233604 382238
rect 233548 379988 233604 382172
rect 233996 381780 234052 381790
rect 234052 381724 234164 381780
rect 233996 381714 234052 381724
rect 234108 379988 234164 381724
rect 235340 379988 235396 382284
rect 232764 379932 233240 379988
rect 233548 379932 233912 379988
rect 234108 379932 234584 379988
rect 235256 379932 235396 379988
rect 236124 381444 236180 381454
rect 236124 379988 236180 381388
rect 236908 380660 236964 380670
rect 236908 379988 236964 380604
rect 237468 379988 237524 385196
rect 238812 385140 238868 385150
rect 238588 381892 238644 381902
rect 238644 381836 238756 381892
rect 238588 381826 238644 381836
rect 238700 379988 238756 381836
rect 236124 379932 236600 379988
rect 236908 379932 237272 379988
rect 237468 379932 237944 379988
rect 238616 379932 238756 379988
rect 238812 379988 238868 385084
rect 239372 383460 239428 383470
rect 239428 383404 239540 383460
rect 239372 383394 239428 383404
rect 239484 379988 239540 383404
rect 240268 382676 240324 382686
rect 240268 379988 240324 382620
rect 240828 379988 240884 386876
rect 242844 386820 242900 386830
rect 242172 386708 242228 386718
rect 242060 385364 242116 385374
rect 242060 379988 242116 385308
rect 238812 379932 239288 379988
rect 239484 379932 239960 379988
rect 240268 379932 240632 379988
rect 240828 379932 241304 379988
rect 241976 379932 242116 379988
rect 242172 379988 242228 386652
rect 242844 379988 242900 386764
rect 247100 386596 247156 386606
rect 246204 385476 246260 385486
rect 245420 385028 245476 385038
rect 244076 381668 244132 381678
rect 244132 381612 244244 381668
rect 244076 381602 244132 381612
rect 243740 381556 243796 381566
rect 243740 379988 243796 381500
rect 244188 379988 244244 381612
rect 245420 379988 245476 384972
rect 242172 379932 242648 379988
rect 242844 379932 243320 379988
rect 243740 379932 243992 379988
rect 244188 379932 244664 379988
rect 245336 379932 245476 379988
rect 245532 382004 245588 382014
rect 245532 379988 245588 381948
rect 246204 379988 246260 385420
rect 247100 379988 247156 386540
rect 248556 385812 248612 385822
rect 248556 379988 248612 385756
rect 248780 379988 248836 396452
rect 250012 384748 250068 400652
rect 249900 384692 250068 384748
rect 250572 390628 250628 390638
rect 249788 382004 249844 382014
rect 249788 379988 249844 381948
rect 245532 379932 246008 379988
rect 246204 379932 246680 379988
rect 247100 379932 247352 379988
rect 248024 379932 248612 379988
rect 248696 379932 248836 379988
rect 249368 379932 249844 379988
rect 249900 379988 249956 384692
rect 250572 379988 250628 390572
rect 251356 384748 251412 405692
rect 252028 404068 252084 405804
rect 252028 404002 252084 404012
rect 251244 384692 251412 384748
rect 252476 385924 252532 385934
rect 251244 379988 251300 384692
rect 252476 379988 252532 385868
rect 252700 384748 252756 406364
rect 259420 405972 259476 405982
rect 257852 404852 257908 404862
rect 249900 379932 250040 379988
rect 250572 379932 250712 379988
rect 251244 379932 251384 379988
rect 252056 379932 252532 379988
rect 252588 384692 252756 384748
rect 253260 390740 253316 390750
rect 252588 379988 252644 384692
rect 253260 379988 253316 390684
rect 256620 385700 256676 385710
rect 255052 383012 255108 383022
rect 254716 382340 254772 382350
rect 254604 382284 254716 382340
rect 254604 379988 254660 382284
rect 254716 382274 254772 382284
rect 255052 379988 255108 382956
rect 256060 382228 256116 382238
rect 255948 382172 256060 382228
rect 255948 379988 256004 382172
rect 256060 382162 256116 382172
rect 256620 379988 256676 385644
rect 257852 383012 257908 404796
rect 257852 382946 257908 382956
rect 257964 387380 258020 387390
rect 256956 382788 257012 382798
rect 256956 379988 257012 382732
rect 257964 379988 258020 387324
rect 259420 384748 259476 405916
rect 259308 384692 259476 384748
rect 260316 387492 260372 387502
rect 258636 382452 258692 382462
rect 258636 379988 258692 382396
rect 259196 382004 259252 382014
rect 259196 379988 259252 381948
rect 252588 379932 252728 379988
rect 253260 379932 253400 379988
rect 254072 379932 254660 379988
rect 254744 379932 255108 379988
rect 255416 379932 256004 379988
rect 256088 379932 256676 379988
rect 256760 379932 257012 379988
rect 257432 379932 258020 379988
rect 258104 379932 258692 379988
rect 258776 379932 259252 379988
rect 259308 379988 259364 384692
rect 260316 379988 260372 387436
rect 260428 380884 260484 406588
rect 261212 405860 261268 405870
rect 261212 382340 261268 405804
rect 262780 404740 262836 404750
rect 262108 399140 262164 399150
rect 262108 396508 262164 399084
rect 262108 396452 262276 396508
rect 261212 382274 261268 382284
rect 261324 382676 261380 382686
rect 260428 380818 260484 380828
rect 261324 379988 261380 382620
rect 261996 382340 262052 382350
rect 261996 379988 262052 382284
rect 262220 379988 262276 396452
rect 262780 384748 262836 404684
rect 263452 399252 263508 399262
rect 263452 384748 263508 399196
rect 259308 379932 259448 379988
rect 260120 379932 260372 379988
rect 260792 379932 261380 379988
rect 261464 379932 262052 379988
rect 262136 379932 262276 379988
rect 262668 384692 262836 384748
rect 263340 384692 263508 384748
rect 262668 379988 262724 384692
rect 263340 379988 263396 384692
rect 263788 380772 263844 407708
rect 268156 408660 268212 408670
rect 266812 404628 266868 404638
rect 264124 402948 264180 402958
rect 264124 384748 264180 402892
rect 265468 399812 265524 399822
rect 264796 399364 264852 399374
rect 264796 384748 264852 399308
rect 265468 396508 265524 399756
rect 265468 396452 265636 396508
rect 263788 380706 263844 380716
rect 264012 384692 264180 384748
rect 264684 384692 264852 384748
rect 264012 379988 264068 384692
rect 264684 379988 264740 384692
rect 265580 379988 265636 396452
rect 266812 384748 266868 404572
rect 267484 402500 267540 402510
rect 267484 384748 267540 402444
rect 268156 384748 268212 408604
rect 268940 407876 268996 410060
rect 266700 384692 266868 384748
rect 267372 384692 267540 384748
rect 268044 384692 268212 384748
rect 268828 400820 268884 400830
rect 268828 384748 268884 400764
rect 268940 386036 268996 407820
rect 274652 407988 274708 410060
rect 280476 409444 280532 410060
rect 268940 385970 268996 385980
rect 270172 401380 270228 401390
rect 270172 384748 270228 401324
rect 274204 401268 274260 401278
rect 271516 401044 271572 401054
rect 268828 384692 268996 384748
rect 266588 382004 266644 382014
rect 266588 379988 266644 381948
rect 262668 379932 262808 379988
rect 263340 379932 263480 379988
rect 264012 379932 264152 379988
rect 264684 379932 264824 379988
rect 265496 379932 265636 379988
rect 266168 379932 266644 379988
rect 266700 379988 266756 384692
rect 267372 379988 267428 384692
rect 268044 379988 268100 384692
rect 268940 379988 268996 384692
rect 270060 384692 270228 384748
rect 270732 396340 270788 396350
rect 269948 384244 270004 384254
rect 269948 379988 270004 384188
rect 266700 379932 266840 379988
rect 267372 379932 267512 379988
rect 268044 379932 268184 379988
rect 268856 379932 268996 379988
rect 269528 379932 270004 379988
rect 270060 379988 270116 384692
rect 270732 379988 270788 396284
rect 271516 384748 271572 400988
rect 272860 400932 272916 400942
rect 271404 384692 271572 384748
rect 272300 396228 272356 396238
rect 271404 379988 271460 384692
rect 272300 379988 272356 396172
rect 272860 384748 272916 400876
rect 270060 379932 270200 379988
rect 270732 379932 270872 379988
rect 271404 379932 271544 379988
rect 272216 379932 272356 379988
rect 272748 384692 272916 384748
rect 273420 396004 273476 396014
rect 272748 379988 272804 384692
rect 273420 379988 273476 395948
rect 274204 384748 274260 401212
rect 274092 384692 274260 384748
rect 274652 385028 274708 407932
rect 280252 408436 280308 408446
rect 279580 402724 279636 402734
rect 278236 402612 278292 402622
rect 275548 401156 275604 401166
rect 275548 396508 275604 401100
rect 275548 396452 275716 396508
rect 274092 379988 274148 384692
rect 274652 380660 274708 384972
rect 274652 380594 274708 380604
rect 274764 395892 274820 395902
rect 274764 379988 274820 395836
rect 275660 379988 275716 396452
rect 272748 379932 272888 379988
rect 273420 379932 273560 379988
rect 274092 379932 274232 379988
rect 274764 379932 274904 379988
rect 275576 379932 275716 379988
rect 276108 395780 276164 395790
rect 276108 379988 276164 395724
rect 277452 395668 277508 395678
rect 276780 394548 276836 394558
rect 276780 379988 276836 394492
rect 277452 379988 277508 395612
rect 278236 384748 278292 402556
rect 279580 384748 279636 402668
rect 280252 384748 280308 408380
rect 280476 406644 280532 409388
rect 283948 409556 284004 409566
rect 280476 406578 280532 406588
rect 282268 409108 282324 409118
rect 280924 402836 280980 402846
rect 280924 384748 280980 402780
rect 282268 396508 282324 409052
rect 283612 406308 283668 406318
rect 282268 396452 282436 396508
rect 278124 384692 278292 384748
rect 279468 384692 279636 384748
rect 280140 384692 280308 384748
rect 280812 384692 280980 384748
rect 278124 379988 278180 384692
rect 279356 382116 279412 382126
rect 279356 379988 279412 382060
rect 276108 379932 276248 379988
rect 276780 379932 276920 379988
rect 277452 379932 277592 379988
rect 278124 379932 278264 379988
rect 278936 379932 279412 379988
rect 279468 379988 279524 384692
rect 280140 379988 280196 384692
rect 280812 379988 280868 384692
rect 281708 382004 281764 382014
rect 281708 379988 281764 381948
rect 282380 379988 282436 396452
rect 283388 386036 283444 386046
rect 283388 379988 283444 385980
rect 283612 384748 283668 406252
rect 279468 379932 279608 379988
rect 280140 379932 280280 379988
rect 280812 379932 280952 379988
rect 281624 379932 281764 379988
rect 282296 379932 282436 379988
rect 282968 379932 283444 379988
rect 283500 384692 283668 384748
rect 283500 379988 283556 384692
rect 283948 384468 284004 409500
rect 285180 409556 285236 410088
rect 285180 409490 285236 409500
rect 289772 410060 290360 410116
rect 295512 410060 295652 410116
rect 305816 410088 306628 410116
rect 310968 410088 311668 410116
rect 289772 409220 289828 410060
rect 286300 406196 286356 406206
rect 284732 404292 284788 404302
rect 284284 399476 284340 399486
rect 284284 384748 284340 399420
rect 283948 384402 284004 384412
rect 284172 384692 284340 384748
rect 284172 379988 284228 384692
rect 284732 382116 284788 404236
rect 286300 384748 286356 406140
rect 288316 399700 288372 399710
rect 286188 384692 286356 384748
rect 286860 390852 286916 390862
rect 284732 382050 284788 382060
rect 285516 382900 285572 382910
rect 285516 379988 285572 382844
rect 286076 382564 286132 382574
rect 286076 379988 286132 382508
rect 283500 379932 283640 379988
rect 284172 379932 284312 379988
rect 284984 379932 285572 379988
rect 285656 379932 286132 379988
rect 286188 379988 286244 384692
rect 286860 379988 286916 390796
rect 288316 384748 288372 399644
rect 288204 384692 288372 384748
rect 288092 382004 288148 382014
rect 288092 379988 288148 381948
rect 286188 379932 286328 379988
rect 286860 379932 287000 379988
rect 287672 379932 288148 379988
rect 288204 379988 288260 384692
rect 289772 384580 289828 409164
rect 295596 408996 295652 410060
rect 295596 406644 295652 408940
rect 295596 406578 295652 406588
rect 298172 409220 298228 409230
rect 297052 397012 297108 397022
rect 294924 392868 294980 392878
rect 293580 392644 293636 392654
rect 291564 387716 291620 387726
rect 289772 384514 289828 384524
rect 290220 387604 290276 387614
rect 289548 382788 289604 382798
rect 289548 379988 289604 382732
rect 290220 379988 290276 387548
rect 290556 382004 290612 382014
rect 290556 379988 290612 381948
rect 291564 379988 291620 387660
rect 292236 382116 292292 382126
rect 292236 379988 292292 382060
rect 293468 382004 293524 382014
rect 292908 380212 292964 380222
rect 292908 379988 292964 380156
rect 293468 379988 293524 381948
rect 288204 379932 288344 379988
rect 289016 379932 289604 379988
rect 289688 379932 290276 379988
rect 290360 379932 290612 379988
rect 291032 379932 291620 379988
rect 291704 379932 292292 379988
rect 292376 379932 292964 379988
rect 293048 379932 293524 379988
rect 293580 379988 293636 392588
rect 294252 390964 294308 390974
rect 294252 379988 294308 390908
rect 294924 379988 294980 392812
rect 295820 391188 295876 391198
rect 295820 379988 295876 391132
rect 296828 387828 296884 387838
rect 296828 379988 296884 387772
rect 297052 384748 297108 396956
rect 293580 379932 293720 379988
rect 294252 379932 294392 379988
rect 294924 379932 295064 379988
rect 295736 379932 295876 379988
rect 296408 379932 296884 379988
rect 296940 384692 297108 384748
rect 298060 387940 298116 387950
rect 296940 379988 296996 384692
rect 298060 379988 298116 387884
rect 298172 382676 298228 409164
rect 300636 408100 300692 410088
rect 305788 410060 306628 410088
rect 305788 409668 305844 410060
rect 305788 409602 305844 409612
rect 300636 408034 300692 408044
rect 300412 401716 300468 401726
rect 299740 399924 299796 399934
rect 299068 396900 299124 396910
rect 299068 396508 299124 396844
rect 299068 396452 299236 396508
rect 298172 382610 298228 382620
rect 298284 394772 298340 394782
rect 296940 379932 297080 379988
rect 297752 379932 298116 379988
rect 298284 379988 298340 394716
rect 299180 379988 299236 396452
rect 299740 384748 299796 399868
rect 300412 384748 300468 401660
rect 303772 398244 303828 398254
rect 302540 396116 302596 396126
rect 298284 379932 298424 379988
rect 299096 379932 299236 379988
rect 299628 384692 299796 384748
rect 300300 384692 300468 384748
rect 301644 394660 301700 394670
rect 299628 379988 299684 384692
rect 300300 379988 300356 384692
rect 301532 382788 301588 382798
rect 301532 379988 301588 382732
rect 299628 379932 299768 379988
rect 300300 379932 300440 379988
rect 301112 379932 301588 379988
rect 301644 379988 301700 394604
rect 302540 379988 302596 396060
rect 303772 384748 303828 398188
rect 305004 394996 305060 395006
rect 303660 384692 303828 384748
rect 304332 394100 304388 394110
rect 303548 382676 303604 382686
rect 303548 379988 303604 382620
rect 301644 379932 301784 379988
rect 302456 379932 302596 379988
rect 303128 379932 303604 379988
rect 303660 379988 303716 384692
rect 304332 379988 304388 394044
rect 305004 379988 305060 394940
rect 305900 394884 305956 394894
rect 305900 379988 305956 394828
rect 306572 380660 306628 410060
rect 310940 410060 311668 410088
rect 310940 409780 310996 410060
rect 310940 409714 310996 409724
rect 307132 408324 307188 408334
rect 307132 384748 307188 408268
rect 308252 404180 308308 404190
rect 307020 384692 307188 384748
rect 307692 394324 307748 394334
rect 306572 380594 306628 380604
rect 306908 382116 306964 382126
rect 306908 379988 306964 382060
rect 303660 379932 303800 379988
rect 304332 379932 304472 379988
rect 305004 379932 305144 379988
rect 305816 379932 305956 379988
rect 306488 379932 306964 379988
rect 307020 379988 307076 384692
rect 307692 379988 307748 394268
rect 308252 382900 308308 404124
rect 310492 397796 310548 397806
rect 309820 396676 309876 396686
rect 308252 382834 308308 382844
rect 308364 393876 308420 393886
rect 308364 379988 308420 393820
rect 309260 391300 309316 391310
rect 309260 379988 309316 391244
rect 309820 384748 309876 396620
rect 310492 384748 310548 397740
rect 307020 379932 307160 379988
rect 307692 379932 307832 379988
rect 308364 379932 308504 379988
rect 309176 379932 309316 379988
rect 309708 384692 309876 384748
rect 310380 384692 310548 384748
rect 311052 391412 311108 391422
rect 309708 379988 309764 384692
rect 310380 379988 310436 384692
rect 311052 379988 311108 391356
rect 311612 380772 311668 410060
rect 316092 396508 316148 410088
rect 315868 396452 316148 396508
rect 313740 390516 313796 390526
rect 313068 382900 313124 382910
rect 311612 380706 311668 380716
rect 312396 382004 312452 382014
rect 312396 379988 312452 381948
rect 313068 379988 313124 382844
rect 313628 382004 313684 382014
rect 313628 379988 313684 381948
rect 309708 379932 309848 379988
rect 310380 379932 310520 379988
rect 311052 379932 311192 379988
rect 311864 379932 312452 379988
rect 312536 379932 313124 379988
rect 313208 379932 313684 379988
rect 313740 379988 313796 390460
rect 315868 384804 315924 396452
rect 320908 389844 320964 389854
rect 320908 388948 320964 389788
rect 321244 389844 321300 410088
rect 324604 397572 324660 397582
rect 323932 397460 323988 397470
rect 321244 389778 321300 389788
rect 321804 391076 321860 391086
rect 320908 388882 320964 388892
rect 318444 388164 318500 388174
rect 315868 384356 315924 384748
rect 315868 384290 315924 384300
rect 316092 386148 316148 386158
rect 315084 382004 315140 382014
rect 315084 379988 315140 381948
rect 315196 380996 315252 381006
rect 315252 380940 315364 380996
rect 315196 380930 315252 380940
rect 315308 379988 315364 380940
rect 315868 380548 315924 380558
rect 315924 380492 316036 380548
rect 315868 380482 315924 380492
rect 315980 379988 316036 380492
rect 313740 379932 313880 379988
rect 314552 379932 315140 379988
rect 315224 379932 315364 379988
rect 315896 379932 316036 379988
rect 316092 379988 316148 386092
rect 316652 383572 316708 383582
rect 316708 383516 316820 383572
rect 316652 383506 316708 383516
rect 316764 379988 316820 383516
rect 318444 379988 318500 388108
rect 320012 383012 320068 383022
rect 320012 382116 320068 382956
rect 320012 382050 320068 382060
rect 319340 380324 319396 380334
rect 319396 380268 319508 380324
rect 319340 380258 319396 380268
rect 319452 379988 319508 380268
rect 320908 380100 320964 380110
rect 320572 379988 320628 379998
rect 316092 379932 316568 379988
rect 316764 379932 317240 379988
rect 318444 379932 318584 379988
rect 319452 379932 319928 379988
rect 320908 379988 320964 380044
rect 321804 379988 321860 391020
rect 322700 385588 322756 385598
rect 322700 379988 322756 385532
rect 323932 384748 323988 397404
rect 324604 384748 324660 397516
rect 326396 396508 326452 410088
rect 329308 397684 329364 397694
rect 325948 396452 326452 396508
rect 328636 397348 328692 397358
rect 323820 384692 323988 384748
rect 324492 384692 324660 384748
rect 325164 392420 325220 392430
rect 320908 379932 321272 379988
rect 321804 379932 321944 379988
rect 322616 379932 322756 379988
rect 322924 382004 322980 382014
rect 322924 379988 322980 381948
rect 323820 379988 323876 384692
rect 324492 379988 324548 384692
rect 325164 379988 325220 392364
rect 325836 384916 325892 384926
rect 325836 384804 325892 384860
rect 325948 384804 326004 396452
rect 325836 384748 326004 384804
rect 327180 392308 327236 392318
rect 325836 380548 325892 384748
rect 325948 384132 326004 384142
rect 326004 384076 326116 384132
rect 325948 384066 326004 384076
rect 325836 380482 325892 380492
rect 326060 379988 326116 384076
rect 322924 379932 323288 379988
rect 323820 379932 323960 379988
rect 324492 379932 324632 379988
rect 325164 379932 325304 379988
rect 325976 379932 326116 379988
rect 326284 384020 326340 384030
rect 326284 379988 326340 383964
rect 327180 379988 327236 392252
rect 328636 384748 328692 397292
rect 329308 396508 329364 397628
rect 329308 396452 329476 396508
rect 328524 384692 328692 384748
rect 327628 383908 327684 383918
rect 327628 379988 327684 383852
rect 328524 379988 328580 384692
rect 329420 379988 329476 396452
rect 331548 381332 331604 410088
rect 336700 383908 336756 410088
rect 336700 383842 336756 383852
rect 341180 409332 341236 409342
rect 331548 381266 331604 381276
rect 339388 383124 339444 383134
rect 326284 379932 326648 379988
rect 327180 379932 327320 379988
rect 327628 379932 327992 379988
rect 328524 379932 328664 379988
rect 329336 379932 329476 379988
rect 320572 379922 320628 379932
rect 319228 379876 319284 379886
rect 319228 379810 319284 379820
rect 200844 379764 200900 379774
rect 202188 379764 202244 379774
rect 200312 379708 200844 379764
rect 201656 379708 202188 379764
rect 200844 379698 200900 379708
rect 202188 379698 202244 379708
rect 220444 379652 220500 379662
rect 220444 379586 220500 379596
rect 222012 379540 222068 379550
rect 224028 379540 224084 379550
rect 227612 379540 227668 379550
rect 229068 379540 229124 379550
rect 222068 379484 222488 379540
rect 224084 379484 224504 379540
rect 227192 379484 227612 379540
rect 228536 379484 229068 379540
rect 222012 379474 222068 379484
rect 224028 379474 224084 379484
rect 227612 379474 227668 379484
rect 229068 379474 229124 379484
rect 230524 379540 230580 379550
rect 230524 379474 230580 379484
rect 235452 379540 235508 379550
rect 235508 379484 235928 379540
rect 235452 379474 235508 379484
rect 317884 379428 317940 379438
rect 317884 379362 317940 379372
rect 221116 379316 221172 379326
rect 221116 379250 221172 379260
rect 221788 379316 221844 379326
rect 221788 379250 221844 379260
rect 225148 379316 225204 379326
rect 225148 379250 225204 379260
rect 225820 379316 225876 379326
rect 225820 379250 225876 379260
rect 227836 379316 227892 379326
rect 227836 379250 227892 379260
rect 232540 379316 232596 379326
rect 232540 379250 232596 379260
rect 339388 344260 339444 383068
rect 340172 380212 340228 380222
rect 339388 344194 339444 344204
rect 339612 356356 339668 356366
rect 189756 270050 189812 270060
rect 339500 271236 339556 271246
rect 189532 268930 189588 268940
rect 339388 267764 339444 267774
rect 338716 241556 338772 241566
rect 338492 241554 338772 241556
rect 338492 241502 338718 241554
rect 338770 241502 338772 241554
rect 338492 241500 338772 241502
rect 194908 240212 194964 240222
rect 194908 240146 194964 240156
rect 189308 229842 189364 229852
rect 195804 224308 195860 240072
rect 196700 232932 196756 240072
rect 196700 232866 196756 232876
rect 195804 224242 195860 224252
rect 189196 219426 189252 219436
rect 189084 217858 189140 217868
rect 188076 214722 188132 214732
rect 197596 212660 197652 240072
rect 198492 227780 198548 240072
rect 199388 227892 199444 240072
rect 199388 227826 199444 227836
rect 198492 227714 198548 227724
rect 200284 224532 200340 240072
rect 200284 224466 200340 224476
rect 201180 217588 201236 240072
rect 201180 217522 201236 217532
rect 202076 212772 202132 240072
rect 202972 222740 203028 240072
rect 203868 229572 203924 240072
rect 203868 229506 203924 229516
rect 204764 224420 204820 240072
rect 205660 234500 205716 240072
rect 205660 234434 205716 234444
rect 206556 234388 206612 240072
rect 207452 234612 207508 240072
rect 208348 236964 208404 240072
rect 208348 236898 208404 236908
rect 207452 234546 207508 234556
rect 206556 234322 206612 234332
rect 209244 231588 209300 240072
rect 210140 231812 210196 240072
rect 210140 231746 210196 231756
rect 209244 231522 209300 231532
rect 211036 231476 211092 240072
rect 211932 231700 211988 240072
rect 211932 231634 211988 231644
rect 211036 231410 211092 231420
rect 212828 230916 212884 240072
rect 212828 230850 212884 230860
rect 213724 227780 213780 240072
rect 214620 227892 214676 240072
rect 215516 228340 215572 240072
rect 216412 228452 216468 240072
rect 216412 228386 216468 228396
rect 215516 228274 215572 228284
rect 214620 227826 214676 227836
rect 213724 227714 213780 227724
rect 217308 227556 217364 240072
rect 217308 227490 217364 227500
rect 204764 224354 204820 224364
rect 218204 224196 218260 240072
rect 219100 225092 219156 240072
rect 219100 225026 219156 225036
rect 219996 224308 220052 240072
rect 220892 224420 220948 240072
rect 221788 224532 221844 240072
rect 221788 224466 221844 224476
rect 220892 224354 220948 224364
rect 219996 224242 220052 224252
rect 218204 224130 218260 224140
rect 202972 222674 203028 222684
rect 222684 221508 222740 240072
rect 223580 234500 223636 240072
rect 223580 234434 223636 234444
rect 224476 221620 224532 240072
rect 224476 221554 224532 221564
rect 222684 221442 222740 221452
rect 225372 214228 225428 240072
rect 226268 236964 226324 240072
rect 226268 236898 226324 236908
rect 227164 221060 227220 240072
rect 228060 232820 228116 240072
rect 228060 232754 228116 232764
rect 227164 220994 227220 221004
rect 228956 215908 229012 240072
rect 228956 215842 229012 215852
rect 229852 214340 229908 240072
rect 230748 214452 230804 240072
rect 230748 214386 230804 214396
rect 229852 214274 229908 214284
rect 225372 214162 225428 214172
rect 202076 212706 202132 212716
rect 197596 212594 197652 212604
rect 231644 212548 231700 240072
rect 232540 225988 232596 240072
rect 233436 236964 233492 240072
rect 233436 236898 233492 236908
rect 234332 234276 234388 240072
rect 235228 237076 235284 240072
rect 236152 240044 236740 240100
rect 235228 237010 235284 237020
rect 236684 236964 236740 240044
rect 236684 236898 236740 236908
rect 237020 236964 237076 240072
rect 237020 236898 237076 236908
rect 234332 234210 234388 234220
rect 237916 232820 237972 240072
rect 238812 236964 238868 240072
rect 238812 236898 238868 236908
rect 239708 232932 239764 240072
rect 240604 236964 240660 240072
rect 240604 236898 240660 236908
rect 239708 232866 239764 232876
rect 237916 232754 237972 232764
rect 232540 225922 232596 225932
rect 241500 213332 241556 240072
rect 242396 237076 242452 240072
rect 243320 240044 243572 240100
rect 242396 237010 242452 237020
rect 243516 236964 243572 240044
rect 244188 238532 244244 240072
rect 244188 238466 244244 238476
rect 245084 238532 245140 240072
rect 245084 238466 245140 238476
rect 245980 237748 246036 240072
rect 246876 238308 246932 240072
rect 246876 238242 246932 238252
rect 247772 237860 247828 240072
rect 248668 237972 248724 240072
rect 249564 238084 249620 240072
rect 250460 238420 250516 240072
rect 250460 238354 250516 238364
rect 251356 238196 251412 240072
rect 252252 238532 252308 240072
rect 252252 238466 252308 238476
rect 251356 238130 251412 238140
rect 249564 238018 249620 238028
rect 248668 237906 248724 237916
rect 247772 237794 247828 237804
rect 245980 237682 246036 237692
rect 253148 237524 253204 240072
rect 253148 237458 253204 237468
rect 243516 236898 243572 236908
rect 254044 215012 254100 240072
rect 254044 214946 254100 214956
rect 254940 214340 254996 240072
rect 255836 215908 255892 240072
rect 255836 215842 255892 215852
rect 254940 214274 254996 214284
rect 241500 213266 241556 213276
rect 231644 212482 231700 212492
rect 256732 212436 256788 240072
rect 257628 214116 257684 240072
rect 258524 214452 258580 240072
rect 259420 216580 259476 240072
rect 259420 216514 259476 216524
rect 258524 214386 258580 214396
rect 257628 214050 257684 214060
rect 260316 212548 260372 240072
rect 260316 212482 260372 212492
rect 256732 212370 256788 212380
rect 261212 209972 261268 240072
rect 262108 216692 262164 240072
rect 262108 216626 262164 216636
rect 263004 210756 263060 240072
rect 263900 211540 263956 240072
rect 263900 211474 263956 211484
rect 263004 210690 263060 210700
rect 264796 210084 264852 240072
rect 265692 211652 265748 240072
rect 266616 240044 267092 240100
rect 267036 236964 267092 240044
rect 267484 237076 267540 240072
rect 268408 240044 268660 240100
rect 267484 237010 267540 237020
rect 267036 236898 267092 236908
rect 268604 236964 268660 240044
rect 268604 236898 268660 236908
rect 265692 211586 265748 211596
rect 264796 210018 264852 210028
rect 261212 209906 261268 209916
rect 269052 209636 269108 209646
rect 269052 209188 269108 209580
rect 269052 209122 269108 209132
rect 269276 145348 269332 240072
rect 269724 238532 269780 238542
rect 269612 237524 269668 237534
rect 269276 145282 269332 145292
rect 269388 227556 269444 227566
rect 41132 49634 41188 49644
rect 45612 50148 45668 50158
rect 161756 50148 161812 50158
rect 41020 49522 41076 49532
rect 40796 47954 40852 47964
rect 40236 46946 40292 46956
rect 45388 47012 45444 47022
rect 45388 5908 45444 46956
rect 45388 5842 45444 5852
rect 40124 4946 40180 4956
rect 40012 4834 40068 4844
rect 42028 4676 42084 4686
rect 41804 4228 41860 4238
rect 41804 480 41860 4172
rect 42028 4228 42084 4620
rect 42028 4162 42084 4172
rect 45612 480 45668 50092
rect 49868 49812 49924 49822
rect 49644 49700 49700 49710
rect 46956 47908 47012 47918
rect 46956 47124 47012 47852
rect 46956 47058 47012 47068
rect 47516 4340 47572 4350
rect 47516 480 47572 4284
rect 49644 4340 49700 49644
rect 49644 4274 49700 4284
rect 49420 4228 49476 4238
rect 49420 480 49476 4172
rect 49868 4228 49924 49756
rect 87500 49588 87556 49598
rect 49868 4162 49924 4172
rect 53228 48244 53284 48254
rect 53228 480 53284 48188
rect 77980 48132 78036 48142
rect 62748 46228 62804 46238
rect 60844 5012 60900 5022
rect 58940 4116 58996 4126
rect 55132 3444 55188 3454
rect 55132 480 55188 3388
rect 57148 3444 57204 3454
rect 57148 480 57204 3388
rect 58940 480 58996 4060
rect 60844 480 60900 4956
rect 62748 480 62804 46172
rect 68460 42868 68516 42878
rect 64652 4900 64708 4910
rect 64652 480 64708 4844
rect 66556 4788 66612 4798
rect 66556 480 66612 4732
rect 68460 480 68516 42812
rect 76076 4676 76132 4686
rect 72268 4564 72324 4574
rect 70364 4452 70420 4462
rect 70364 480 70420 4396
rect 72268 480 72324 4508
rect 74396 4116 74452 4126
rect 74396 480 74452 4060
rect 34188 392 34440 480
rect 32312 -960 32536 392
rect 34216 -960 34440 392
rect 36120 -960 36344 480
rect 37996 392 38248 480
rect 39900 392 40152 480
rect 41804 392 42056 480
rect 38024 -960 38248 392
rect 39928 -960 40152 392
rect 41832 -960 42056 392
rect 43736 -960 43960 480
rect 45612 392 45864 480
rect 47516 392 47768 480
rect 49420 392 49672 480
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 480
rect 53228 392 53480 480
rect 55132 392 55384 480
rect 53256 -960 53480 392
rect 55160 -960 55384 392
rect 57064 -960 57288 480
rect 58940 392 59192 480
rect 60844 392 61096 480
rect 62748 392 63000 480
rect 64652 392 64904 480
rect 66556 392 66808 480
rect 68460 392 68712 480
rect 70364 392 70616 480
rect 72268 392 72520 480
rect 58968 -960 59192 392
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 70392 -960 70616 392
rect 72296 -960 72520 392
rect 74200 392 74452 480
rect 76076 480 76132 4620
rect 77980 480 78036 48076
rect 81788 48020 81844 48030
rect 79884 41188 79940 41198
rect 79884 480 79940 41132
rect 81788 480 81844 47964
rect 85708 41300 85764 41310
rect 83692 37828 83748 37838
rect 83692 480 83748 37772
rect 85708 480 85764 41244
rect 87500 480 87556 49532
rect 95116 49588 95172 49598
rect 91308 41412 91364 41422
rect 89628 4116 89684 4126
rect 89628 480 89684 4060
rect 76076 392 76328 480
rect 77980 392 78232 480
rect 79884 392 80136 480
rect 81788 392 82040 480
rect 83692 392 83944 480
rect 74200 -960 74424 392
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 83720 -960 83944 392
rect 85624 -960 85848 480
rect 87500 392 87752 480
rect 87528 -960 87752 392
rect 89432 392 89684 480
rect 91308 480 91364 41356
rect 93212 4340 93268 4350
rect 93212 480 93268 4284
rect 95116 480 95172 49532
rect 97356 48692 97412 50120
rect 269388 50148 269444 227500
rect 156044 50036 156100 50046
rect 150332 49924 150388 49934
rect 144620 49812 144676 49822
rect 97356 47908 97412 48636
rect 97356 47842 97412 47852
rect 112252 49700 112308 49710
rect 106540 44660 106596 44670
rect 100828 44548 100884 44558
rect 97244 4900 97300 4910
rect 97244 480 97300 4844
rect 91308 392 91560 480
rect 93212 392 93464 480
rect 95116 392 95368 480
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 392 97300 480
rect 98924 4228 98980 4238
rect 98924 480 98980 4172
rect 100828 480 100884 44492
rect 102956 4228 103012 4238
rect 102956 480 103012 4172
rect 104860 4116 104916 4126
rect 104860 480 104916 4060
rect 98924 392 99176 480
rect 100828 392 101080 480
rect 97048 -960 97272 392
rect 98952 -960 99176 392
rect 100856 -960 101080 392
rect 102760 392 103012 480
rect 104664 392 104916 480
rect 106540 480 106596 44604
rect 108444 41524 108500 41534
rect 108444 480 108500 41468
rect 110796 4228 110852 4238
rect 110572 4172 110796 4228
rect 110572 480 110628 4172
rect 110796 4162 110852 4172
rect 106540 392 106792 480
rect 108444 392 108696 480
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 -960 108696 392
rect 110376 392 110628 480
rect 112252 480 112308 49644
rect 138908 48244 138964 48254
rect 133196 48132 133252 48142
rect 127484 48020 127540 48030
rect 121772 47908 121828 47918
rect 119868 43092 119924 43102
rect 114268 42980 114324 42990
rect 114268 480 114324 42924
rect 117964 41636 118020 41646
rect 116284 4340 116340 4350
rect 116284 480 116340 4284
rect 112252 392 112504 480
rect 110376 -960 110600 392
rect 112280 -960 112504 392
rect 114184 -960 114408 480
rect 116088 392 116340 480
rect 117964 480 118020 41580
rect 119868 480 119924 43036
rect 121772 480 121828 47852
rect 125580 46340 125636 46350
rect 123676 41748 123732 41758
rect 123676 480 123732 41692
rect 125580 480 125636 46284
rect 127484 480 127540 47964
rect 131292 46452 131348 46462
rect 129388 41972 129444 41982
rect 129388 480 129444 41916
rect 131292 480 131348 46396
rect 133196 480 133252 48076
rect 135324 4452 135380 4462
rect 135324 480 135380 4396
rect 137228 3444 137284 3454
rect 137228 480 137284 3388
rect 117964 392 118216 480
rect 119868 392 120120 480
rect 121772 392 122024 480
rect 123676 392 123928 480
rect 125580 392 125832 480
rect 127484 392 127736 480
rect 129388 392 129640 480
rect 131292 392 131544 480
rect 133196 392 133448 480
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 392
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 392 135380 480
rect 137032 392 137284 480
rect 138908 480 138964 48188
rect 142828 43204 142884 43214
rect 140812 38276 140868 38286
rect 140812 480 140868 38220
rect 142828 480 142884 43148
rect 144620 480 144676 49756
rect 146524 38164 146580 38174
rect 146524 480 146580 38108
rect 148652 3444 148708 3454
rect 148652 480 148708 3388
rect 138908 392 139160 480
rect 140812 392 141064 480
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144620 392 144872 480
rect 146524 392 146776 480
rect 144648 -960 144872 392
rect 146552 -960 146776 392
rect 148456 392 148708 480
rect 150332 480 150388 49868
rect 152236 44772 152292 44782
rect 152236 480 152292 44716
rect 154476 4116 154532 4126
rect 154364 4060 154476 4116
rect 154364 480 154420 4060
rect 154476 4050 154532 4060
rect 150332 392 150584 480
rect 152236 392 152488 480
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 392 154420 480
rect 156044 480 156100 49980
rect 158172 5908 158228 5918
rect 158172 480 158228 5852
rect 160076 4564 160132 4574
rect 160076 480 160132 4508
rect 156044 392 156296 480
rect 154168 -960 154392 392
rect 156072 -960 156296 392
rect 157976 392 158228 480
rect 159880 392 160132 480
rect 161756 480 161812 50092
rect 201740 48580 201796 48590
rect 196028 48356 196084 48366
rect 190316 45332 190372 45342
rect 184604 45220 184660 45230
rect 178892 45108 178948 45118
rect 173180 44996 173236 45006
rect 167468 44884 167524 44894
rect 163884 7588 163940 7598
rect 163884 480 163940 7532
rect 165788 4788 165844 4798
rect 165788 480 165844 4732
rect 161756 392 162008 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 392 163940 480
rect 165592 392 165844 480
rect 167468 480 167524 44828
rect 169372 29428 169428 29438
rect 169372 480 169428 29372
rect 171500 4676 171556 4686
rect 171500 480 171556 4620
rect 167468 392 167720 480
rect 169372 392 169624 480
rect 163688 -960 163912 392
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 392 171556 480
rect 173180 480 173236 44940
rect 175084 43428 175140 43438
rect 175084 480 175140 43372
rect 176988 43316 177044 43326
rect 176988 480 177044 43260
rect 178892 480 178948 45052
rect 180796 41076 180852 41086
rect 180796 480 180852 41020
rect 182700 37940 182756 37950
rect 182700 480 182756 37884
rect 184604 480 184660 45164
rect 188412 38052 188468 38062
rect 186508 31108 186564 31118
rect 186508 480 186564 31052
rect 188412 480 188468 37996
rect 190316 480 190372 45276
rect 192332 41860 192388 41870
rect 192220 12628 192276 12638
rect 192220 480 192276 12572
rect 192332 4900 192388 41804
rect 192332 4834 192388 4844
rect 194348 4900 194404 4910
rect 194348 480 194404 4844
rect 173180 392 173432 480
rect 175084 392 175336 480
rect 176988 392 177240 480
rect 178892 392 179144 480
rect 180796 392 181048 480
rect 182700 392 182952 480
rect 184604 392 184856 480
rect 186508 392 186760 480
rect 188412 392 188664 480
rect 190316 392 190568 480
rect 192220 392 192472 480
rect 171304 -960 171528 392
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 392
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 392 194404 480
rect 196028 480 196084 48300
rect 199948 46564 200004 46574
rect 197932 39508 197988 39518
rect 197932 480 197988 39452
rect 199948 480 200004 46508
rect 201740 480 201796 48524
rect 203644 48468 203700 48478
rect 203644 480 203700 48412
rect 212268 47796 212324 50120
rect 269388 50082 269444 50092
rect 269500 224196 269556 224206
rect 212268 47730 212324 47740
rect 269500 44884 269556 224140
rect 269500 44818 269556 44828
rect 207452 44436 207508 44446
rect 205772 5012 205828 5022
rect 205772 480 205828 4956
rect 196028 392 196280 480
rect 197932 392 198184 480
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 392 205828 480
rect 207452 480 207508 44380
rect 209356 31220 209412 31230
rect 209356 480 209412 31164
rect 269612 31220 269668 237468
rect 269724 48468 269780 238476
rect 269836 210868 269892 210878
rect 269836 207956 269892 210812
rect 269836 207890 269892 207900
rect 270172 147028 270228 240072
rect 270172 146962 270228 146972
rect 270508 238420 270564 238430
rect 269724 48402 269780 48412
rect 269612 31154 269668 31164
rect 270508 12628 270564 238364
rect 270844 228452 270900 228462
rect 270732 227780 270788 227790
rect 270620 225092 270676 225102
rect 270620 44996 270676 225036
rect 270732 48244 270788 227724
rect 270844 50036 270900 228396
rect 270844 49970 270900 49980
rect 270956 228340 271012 228350
rect 270956 49924 271012 228284
rect 271068 133588 271124 240072
rect 271292 231028 271348 231038
rect 271068 133522 271124 133532
rect 271180 227892 271236 227902
rect 270956 49858 271012 49868
rect 271180 49812 271236 227836
rect 271292 196420 271348 230972
rect 271292 196354 271348 196364
rect 271180 49746 271236 49756
rect 271292 145460 271348 145470
rect 270732 48178 270788 48188
rect 270620 44930 270676 44940
rect 271292 36820 271348 145404
rect 271964 106708 272020 240072
rect 272860 238308 272916 240072
rect 272860 238242 272916 238252
rect 273420 239876 273476 239886
rect 272300 235172 272356 235182
rect 272188 209524 272244 209534
rect 272188 180852 272244 209468
rect 272188 180786 272244 180796
rect 272300 153636 272356 235116
rect 272300 149548 272356 153580
rect 272188 149492 272356 149548
rect 272412 211316 272468 211326
rect 272188 131348 272244 149492
rect 272412 148820 272468 211260
rect 272524 209860 272580 209870
rect 272524 157556 272580 209804
rect 272748 209636 272804 209646
rect 272636 209524 272692 209534
rect 272636 166292 272692 209468
rect 272748 175028 272804 209580
rect 272860 209188 272916 209198
rect 272860 177940 272916 209132
rect 272860 177874 272916 177884
rect 272972 203140 273028 203150
rect 272748 174962 272804 174972
rect 272636 166226 272692 166236
rect 272524 157490 272580 157500
rect 272412 148754 272468 148764
rect 272188 131282 272244 131292
rect 272300 143668 272356 143678
rect 271964 106642 272020 106652
rect 272300 50260 272356 143612
rect 272412 140308 272468 140318
rect 272412 50372 272468 140252
rect 272972 99316 273028 203084
rect 273308 154420 273364 154430
rect 273084 154196 273140 154206
rect 273084 134260 273140 154140
rect 273084 134194 273140 134204
rect 273196 144564 273252 144574
rect 273196 128436 273252 144508
rect 273308 137172 273364 154364
rect 273308 137106 273364 137116
rect 273196 128370 273252 128380
rect 273420 105140 273476 239820
rect 273756 237636 273812 240072
rect 273756 237570 273812 237580
rect 273980 238084 274036 238094
rect 273756 234500 273812 234510
rect 273756 202468 273812 234444
rect 273756 202402 273812 202412
rect 273868 213332 273924 213342
rect 273420 105074 273476 105084
rect 272972 99250 273028 99260
rect 273084 91588 273140 91598
rect 272972 89908 273028 89918
rect 272972 73108 273028 89852
rect 273084 78932 273140 91532
rect 273084 78866 273140 78876
rect 272972 73042 273028 73052
rect 272412 50306 272468 50316
rect 272972 70196 273028 70206
rect 272300 50194 272356 50204
rect 272972 48132 273028 70140
rect 273196 67284 273252 67294
rect 273084 64372 273140 64382
rect 273084 50036 273140 64316
rect 273084 49970 273140 49980
rect 272972 48066 273028 48076
rect 273196 48020 273252 67228
rect 273756 58548 273812 58558
rect 273756 49924 273812 58492
rect 273756 49858 273812 49868
rect 273196 47954 273252 47964
rect 271292 36754 271348 36764
rect 270508 12562 270564 12572
rect 273868 4452 273924 213276
rect 273980 31108 274036 238028
rect 274092 237972 274148 237982
rect 274092 41076 274148 237916
rect 274652 105028 274708 240072
rect 274764 227668 274820 227678
rect 274764 200788 274820 227612
rect 274764 200722 274820 200732
rect 274652 104962 274708 104972
rect 274764 128548 274820 128558
rect 274764 81844 274820 128492
rect 275548 125188 275604 240072
rect 276332 239764 276388 239774
rect 275548 125122 275604 125132
rect 275660 238196 275716 238206
rect 274764 81778 274820 81788
rect 274876 107156 274932 107166
rect 274876 76020 274932 107100
rect 274876 75954 274932 75964
rect 274204 52724 274260 52734
rect 274204 49812 274260 52668
rect 274204 49746 274260 49756
rect 274092 41010 274148 41020
rect 275660 39508 275716 238140
rect 275884 224532 275940 224542
rect 275772 224308 275828 224318
rect 275772 45108 275828 224252
rect 275884 45332 275940 224476
rect 275884 45266 275940 45276
rect 275996 224420 276052 224430
rect 275996 45220 276052 224364
rect 275996 45154 276052 45164
rect 276108 221620 276164 221630
rect 275772 45042 275828 45052
rect 276108 44436 276164 221564
rect 276220 221508 276276 221518
rect 276220 48356 276276 221452
rect 276332 199892 276388 239708
rect 276332 199826 276388 199836
rect 276444 115108 276500 240072
rect 277340 131908 277396 240072
rect 277340 131842 277396 131852
rect 278012 238980 278068 238990
rect 276444 115042 276500 115052
rect 276220 48290 276276 48300
rect 276108 44370 276164 44380
rect 275660 39442 275716 39452
rect 273980 31042 274036 31052
rect 273868 4386 273924 4396
rect 211484 4116 211540 4126
rect 211484 480 211540 4060
rect 278012 4116 278068 238924
rect 278236 135268 278292 240072
rect 278236 135202 278292 135212
rect 278908 237748 278964 237758
rect 278908 7588 278964 237692
rect 279132 152292 279188 240072
rect 279132 152226 279188 152236
rect 279692 239652 279748 239662
rect 278908 7522 278964 7532
rect 279692 4788 279748 239596
rect 279916 237636 279972 237646
rect 279804 214116 279860 214126
rect 279804 103348 279860 214060
rect 279916 132020 279972 237580
rect 280028 152740 280084 240072
rect 280028 152674 280084 152684
rect 280588 237860 280644 237870
rect 279916 131954 279972 131964
rect 279804 103282 279860 103292
rect 280588 43428 280644 237804
rect 280924 236964 280980 240072
rect 280924 236898 280980 236908
rect 280700 234612 280756 234622
rect 280700 203140 280756 234556
rect 280700 203074 280756 203084
rect 281372 215012 281428 215022
rect 281372 103796 281428 214956
rect 281820 160244 281876 240072
rect 282716 237524 282772 240072
rect 282716 237458 282772 237468
rect 281820 160178 281876 160188
rect 283052 235060 283108 235070
rect 283052 233492 283108 235004
rect 281372 103730 281428 103740
rect 283052 90580 283108 233436
rect 283612 160356 283668 240072
rect 284508 160692 284564 240072
rect 284508 160626 284564 160636
rect 284732 237748 284788 237758
rect 283612 160290 283668 160300
rect 283052 90514 283108 90524
rect 280588 43362 280644 43372
rect 284732 5012 284788 237692
rect 284956 214228 285012 214238
rect 284844 212436 284900 212446
rect 284844 103684 284900 212380
rect 284844 103618 284900 103628
rect 284732 4946 284788 4956
rect 279692 4722 279748 4732
rect 284956 4228 285012 214172
rect 285404 152180 285460 240072
rect 285404 152114 285460 152124
rect 286300 149044 286356 240072
rect 287196 237636 287252 240072
rect 288120 240044 288260 240100
rect 287196 237570 287252 237580
rect 287980 239876 288036 239886
rect 287980 231868 288036 239820
rect 287980 231812 288148 231868
rect 286300 148978 286356 148988
rect 286412 219828 286468 219838
rect 286412 48244 286468 219772
rect 286412 48178 286468 48188
rect 286524 214788 286580 214798
rect 286524 45332 286580 214732
rect 286524 45266 286580 45276
rect 288092 4676 288148 231812
rect 288204 152628 288260 240044
rect 288428 236964 288484 236974
rect 288204 152562 288260 152572
rect 288316 216580 288372 216590
rect 288316 103572 288372 216524
rect 288428 155876 288484 236908
rect 288428 155810 288484 155820
rect 288988 150948 289044 240072
rect 289100 239316 289156 239326
rect 289100 238532 289156 239260
rect 289100 238466 289156 238476
rect 289772 218036 289828 218046
rect 288988 150882 289044 150892
rect 289660 216692 289716 216702
rect 288316 103506 288372 103516
rect 289660 103460 289716 216636
rect 289660 103394 289716 103404
rect 288204 61460 288260 61470
rect 288204 49700 288260 61404
rect 288204 49634 288260 49644
rect 288988 55636 289044 55646
rect 288988 49588 289044 55580
rect 288988 49522 289044 49532
rect 289772 33684 289828 217980
rect 289884 149156 289940 240072
rect 289884 149090 289940 149100
rect 289996 239316 290052 239326
rect 289772 33618 289828 33628
rect 289996 4900 290052 239260
rect 290780 236964 290836 240072
rect 290780 236898 290836 236908
rect 291564 238308 291620 238318
rect 290332 216356 290388 216366
rect 290108 216244 290164 216254
rect 290108 48580 290164 216188
rect 290108 48514 290164 48524
rect 290332 48468 290388 216300
rect 291452 214452 291508 214462
rect 290332 48402 290388 48412
rect 290556 213220 290612 213230
rect 290556 48356 290612 213164
rect 291452 103908 291508 214396
rect 291564 138628 291620 238252
rect 291676 155988 291732 240072
rect 291788 237524 291844 237534
rect 291788 160132 291844 237468
rect 291788 160066 291844 160076
rect 291676 155922 291732 155932
rect 292572 155652 292628 240072
rect 293244 237636 293300 237646
rect 292572 155586 292628 155596
rect 293132 215908 293188 215918
rect 291564 138562 291620 138572
rect 293132 104132 293188 215852
rect 293244 162148 293300 237580
rect 293244 162082 293300 162092
rect 293468 155540 293524 240072
rect 293468 155474 293524 155484
rect 294364 151060 294420 240072
rect 294924 236964 294980 236974
rect 294364 150994 294420 151004
rect 294812 214340 294868 214350
rect 293132 104066 293188 104076
rect 291452 103842 291508 103852
rect 294812 103236 294868 214284
rect 294924 155764 294980 236908
rect 294924 155698 294980 155708
rect 295036 212548 295092 212558
rect 295036 104020 295092 212492
rect 295260 152852 295316 240072
rect 295260 152786 295316 152796
rect 296156 150276 296212 240072
rect 296940 197428 296996 197438
rect 296940 157332 296996 197372
rect 296940 157266 296996 157276
rect 297052 155428 297108 240072
rect 297164 237412 297220 237422
rect 297164 158900 297220 237356
rect 297164 158834 297220 158844
rect 297276 237300 297332 237310
rect 297276 158788 297332 237244
rect 297276 158722 297332 158732
rect 297052 155362 297108 155372
rect 297948 150836 298004 240072
rect 298732 204148 298788 204158
rect 298620 200900 298676 200910
rect 298508 199220 298564 199230
rect 298396 195748 298452 195758
rect 298396 156996 298452 195692
rect 298508 157444 298564 199164
rect 298508 157378 298564 157388
rect 298620 157108 298676 200844
rect 298732 157556 298788 204092
rect 298844 159460 298900 240072
rect 298844 159394 298900 159404
rect 298956 237860 299012 237870
rect 298956 159012 299012 237804
rect 299740 159348 299796 240072
rect 300412 237972 300468 237982
rect 299740 159282 299796 159292
rect 299964 197764 300020 197774
rect 298956 158946 299012 158956
rect 298732 157490 298788 157500
rect 299964 157220 300020 197708
rect 300188 197316 300244 197326
rect 300076 196532 300132 196542
rect 300076 157780 300132 196476
rect 300188 160690 300244 197260
rect 300412 160804 300468 237916
rect 300412 160738 300468 160748
rect 300524 237524 300580 237534
rect 300188 160638 300190 160690
rect 300242 160638 300244 160690
rect 300188 160626 300244 160638
rect 300076 157714 300132 157724
rect 299964 157154 300020 157164
rect 298620 157042 298676 157052
rect 298396 156930 298452 156940
rect 297948 150770 298004 150780
rect 296156 150210 296212 150220
rect 300524 149604 300580 237468
rect 300636 159236 300692 240072
rect 301532 236964 301588 240072
rect 302428 237412 302484 240072
rect 303324 237860 303380 240072
rect 303324 237794 303380 237804
rect 302428 237346 302484 237356
rect 301532 236898 301588 236908
rect 304220 236964 304276 240072
rect 305116 237524 305172 240072
rect 305116 237458 305172 237468
rect 306012 237300 306068 240072
rect 306936 240044 307412 240100
rect 306012 237234 306068 237244
rect 304220 236898 304276 236908
rect 307356 236964 307412 240044
rect 307804 237972 307860 240072
rect 308728 240044 309092 240100
rect 307804 237906 307860 237916
rect 307356 236898 307412 236908
rect 309036 236964 309092 240044
rect 309036 236898 309092 236908
rect 309596 236964 309652 240072
rect 309596 236898 309652 236908
rect 302764 234948 302820 234958
rect 301644 217924 301700 217934
rect 300972 211652 301028 211662
rect 300636 159170 300692 159180
rect 300860 205828 300916 205838
rect 300860 156884 300916 205772
rect 300860 156818 300916 156828
rect 300524 149538 300580 149548
rect 300972 106932 301028 211596
rect 301196 211540 301252 211550
rect 301084 199108 301140 199118
rect 301084 157668 301140 199052
rect 301084 157602 301140 157612
rect 301196 107044 301252 211484
rect 301644 196952 301700 217868
rect 302764 196952 302820 234892
rect 307244 234836 307300 234846
rect 305004 222964 305060 222974
rect 303884 219604 303940 219614
rect 303884 196952 303940 219548
rect 305004 196952 305060 222908
rect 306124 221284 306180 221294
rect 306124 196952 306180 221228
rect 307244 196952 307300 234780
rect 308364 233268 308420 233278
rect 308364 196952 308420 233212
rect 309484 216020 309540 216030
rect 309484 196952 309540 215964
rect 310492 197988 310548 240072
rect 310492 197922 310548 197932
rect 310604 230020 310660 230030
rect 310604 196952 310660 229964
rect 311388 197876 311444 240072
rect 311388 197810 311444 197820
rect 311724 224868 311780 224878
rect 311724 196952 311780 224812
rect 312284 197540 312340 240072
rect 312284 197474 312340 197484
rect 312844 217812 312900 217822
rect 312844 196952 312900 217756
rect 313180 201124 313236 240072
rect 314076 237860 314132 240072
rect 314076 237794 314132 237804
rect 313180 201058 313236 201068
rect 313964 219492 314020 219502
rect 313964 196952 314020 219436
rect 314972 201012 315028 240072
rect 314972 200946 315028 200956
rect 315084 228228 315140 228238
rect 315084 196952 315140 228172
rect 315868 197652 315924 240072
rect 315868 197586 315924 197596
rect 316204 219380 316260 219390
rect 316204 196952 316260 219324
rect 316764 201236 316820 240072
rect 317660 236964 317716 240072
rect 317660 236898 317716 236908
rect 318444 222852 318500 222862
rect 316764 201170 316820 201180
rect 317324 217700 317380 217710
rect 317324 196952 317380 217644
rect 318444 196952 318500 222796
rect 318556 197204 318612 240072
rect 319452 198212 319508 240072
rect 320348 237972 320404 240072
rect 321244 238084 321300 240072
rect 321244 238018 321300 238028
rect 320348 237906 320404 237916
rect 321804 233156 321860 233166
rect 320684 231364 320740 231374
rect 319452 198146 319508 198156
rect 319564 224756 319620 224766
rect 318556 197138 318612 197148
rect 319564 196952 319620 224700
rect 320684 196952 320740 231308
rect 321804 196952 321860 233100
rect 322140 197316 322196 240072
rect 323064 240044 323876 240100
rect 322140 197250 322196 197260
rect 322924 229796 322980 229806
rect 322924 196952 322980 229740
rect 323820 196532 323876 240044
rect 323932 199332 323988 240072
rect 323932 199266 323988 199276
rect 324044 222628 324100 222638
rect 324044 196952 324100 222572
rect 324828 198100 324884 240072
rect 325276 240044 325752 240100
rect 324828 198034 324884 198044
rect 325164 228116 325220 228126
rect 325164 196952 325220 228060
rect 325276 197204 325332 240044
rect 325276 197138 325332 197148
rect 326284 221172 326340 221182
rect 326284 196952 326340 221116
rect 326620 205828 326676 240072
rect 326620 205762 326676 205772
rect 327404 231252 327460 231262
rect 327404 196952 327460 231196
rect 323820 196466 323876 196476
rect 327516 196532 327572 240072
rect 328412 199220 328468 240072
rect 328412 199154 328468 199164
rect 328524 234724 328580 234734
rect 328524 196952 328580 234668
rect 329308 204148 329364 240072
rect 329308 204082 329364 204092
rect 329644 224644 329700 224654
rect 329644 196952 329700 224588
rect 330204 197764 330260 240072
rect 330204 197698 330260 197708
rect 330764 229908 330820 229918
rect 330764 196952 330820 229852
rect 331100 199108 331156 240072
rect 331100 199042 331156 199052
rect 331884 233044 331940 233054
rect 331884 196952 331940 232988
rect 331996 197428 332052 240072
rect 332892 200900 332948 240072
rect 333816 240044 334292 240100
rect 334236 236964 334292 240044
rect 334236 236898 334292 236908
rect 334684 236964 334740 240072
rect 337372 238084 337428 238094
rect 334684 236898 334740 236908
rect 337148 237972 337204 237982
rect 335244 231140 335300 231150
rect 332892 200834 332948 200844
rect 333004 229684 333060 229694
rect 331996 197362 332052 197372
rect 333004 196952 333060 229628
rect 335132 229460 335188 229470
rect 334124 228004 334180 228014
rect 334124 196952 334180 227948
rect 335132 207508 335188 229404
rect 335132 207442 335188 207452
rect 335244 196952 335300 231084
rect 336924 214676 336980 214686
rect 336812 212660 336868 212670
rect 327516 196466 327572 196476
rect 336364 162484 336420 162494
rect 301308 160692 301364 160702
rect 301308 160690 301896 160692
rect 301308 160638 301310 160690
rect 301362 160638 301896 160690
rect 301308 160636 301896 160638
rect 301308 160626 301364 160636
rect 304332 160580 304388 160590
rect 304388 160524 305032 160580
rect 304332 160514 304388 160524
rect 302876 160468 302932 160478
rect 302932 160412 303464 160468
rect 302876 160402 302932 160412
rect 306572 157892 306628 160104
rect 306572 157826 306628 157836
rect 308140 156996 308196 160104
rect 308140 156930 308196 156940
rect 309708 156884 309764 160104
rect 311276 157780 311332 160104
rect 311276 157714 311332 157724
rect 312844 157444 312900 160104
rect 314412 157556 314468 160104
rect 314412 157490 314468 157500
rect 312844 157378 312900 157388
rect 315980 157220 316036 160104
rect 317548 157668 317604 160104
rect 317548 157602 317604 157612
rect 319116 157332 319172 160104
rect 319116 157266 319172 157276
rect 315980 157154 316036 157164
rect 320684 157108 320740 160104
rect 322252 157892 322308 160104
rect 322252 157826 322308 157836
rect 323820 157220 323876 160104
rect 323820 157154 323876 157164
rect 320684 157042 320740 157052
rect 309708 156818 309764 156828
rect 325388 156884 325444 160104
rect 326956 157556 327012 160104
rect 326956 157490 327012 157500
rect 328524 157444 328580 160104
rect 328524 157378 328580 157388
rect 330092 156996 330148 160104
rect 331660 157332 331716 160104
rect 333228 157780 333284 160104
rect 333228 157714 333284 157724
rect 334796 157668 334852 160104
rect 334796 157602 334852 157612
rect 331660 157266 331716 157276
rect 330092 156930 330148 156940
rect 325388 156818 325444 156828
rect 335916 154532 335972 154542
rect 334684 151396 334740 151406
rect 330092 151284 330148 151294
rect 323372 146244 323428 146254
rect 323372 122612 323428 146188
rect 323372 122546 323428 122556
rect 301196 106978 301252 106988
rect 300972 106866 301028 106876
rect 295036 103954 295092 103964
rect 294812 103170 294868 103180
rect 330092 84756 330148 151228
rect 331772 149716 331828 149726
rect 330876 145572 330932 145582
rect 330876 140308 330932 145516
rect 330876 140242 330932 140252
rect 331772 87668 331828 149660
rect 334684 143668 334740 151340
rect 334684 143602 334740 143612
rect 335132 122724 335188 122734
rect 335132 89908 335188 122668
rect 335916 122724 335972 154476
rect 336364 145460 336420 162428
rect 336364 145394 336420 145404
rect 335916 122658 335972 122668
rect 335132 89842 335188 89852
rect 331772 87602 331828 87612
rect 330092 84690 330148 84700
rect 327516 52948 327572 52958
rect 293580 48692 293636 50120
rect 293580 48626 293636 48636
rect 290556 48290 290612 48300
rect 300748 48244 300804 50120
rect 307916 48356 307972 50120
rect 315084 48468 315140 50120
rect 322252 48580 322308 50120
rect 327516 48692 327572 52892
rect 327516 48626 327572 48636
rect 322252 48514 322308 48524
rect 315084 48402 315140 48412
rect 307916 48290 307972 48300
rect 300748 48178 300804 48188
rect 289996 4834 290052 4844
rect 288092 4610 288148 4620
rect 336812 4340 336868 212604
rect 336924 48692 336980 214620
rect 337036 212772 337092 212782
rect 337036 74900 337092 212716
rect 337148 149492 337204 237916
rect 337148 149426 337204 149436
rect 337260 197988 337316 197998
rect 337260 142660 337316 197932
rect 337372 152404 337428 238028
rect 337596 237860 337652 237870
rect 337596 165508 337652 237804
rect 337596 165442 337652 165452
rect 337372 152338 337428 152348
rect 337260 142594 337316 142604
rect 337036 74834 337092 74844
rect 336924 48626 336980 48636
rect 338492 41300 338548 241500
rect 338716 241490 338772 241500
rect 338940 240548 338996 240558
rect 338604 240436 338660 240446
rect 338604 46340 338660 240380
rect 338604 46274 338660 46284
rect 338716 240324 338772 240334
rect 338716 42868 338772 240268
rect 338828 197876 338884 197886
rect 338828 137732 338884 197820
rect 338828 137666 338884 137676
rect 338940 43204 338996 240492
rect 339388 43316 339444 267708
rect 339500 46564 339556 271180
rect 339612 162820 339668 356300
rect 339724 350196 339780 350206
rect 339724 164164 339780 350140
rect 339724 164098 339780 164108
rect 339836 336084 339892 336094
rect 339612 162754 339668 162764
rect 339836 157108 339892 336028
rect 339948 277060 340004 277070
rect 339948 240212 340004 277004
rect 339948 240146 340004 240156
rect 340060 273924 340116 273934
rect 340060 238532 340116 273868
rect 340060 238466 340116 238476
rect 340172 177156 340228 380156
rect 341068 337316 341124 337326
rect 340284 246708 340340 246718
rect 340284 236292 340340 246652
rect 340956 245364 341012 245374
rect 340956 243348 341012 245308
rect 341068 243572 341124 337260
rect 341180 294308 341236 409276
rect 341852 383124 341908 410088
rect 345212 407316 345268 407326
rect 342748 407092 342804 407102
rect 342748 406756 342804 407036
rect 342748 406690 342804 406700
rect 343532 393204 343588 393214
rect 341852 383058 341908 383068
rect 343196 389060 343252 389070
rect 343084 365092 343140 365102
rect 341180 294242 341236 294252
rect 341852 356132 341908 356142
rect 341292 280532 341348 280542
rect 341292 267148 341348 280476
rect 341180 267092 341348 267148
rect 341180 250068 341236 267092
rect 341180 250002 341236 250012
rect 341292 250404 341348 250414
rect 341292 246932 341348 250348
rect 341292 246866 341348 246876
rect 341068 243516 341348 243572
rect 340956 243292 341124 243348
rect 340396 241556 340452 241566
rect 340396 241462 340452 241500
rect 340956 239540 341012 239550
rect 340508 237748 340564 237758
rect 340284 236226 340340 236236
rect 340396 237636 340452 237646
rect 340396 220108 340452 237580
rect 340172 177090 340228 177100
rect 340284 220052 340452 220108
rect 340284 186564 340340 220052
rect 340284 173068 340340 186508
rect 340508 189252 340564 237692
rect 340956 237636 341012 239484
rect 340956 237570 341012 237580
rect 341068 236404 341124 243292
rect 341068 236338 341124 236348
rect 341292 220108 341348 243516
rect 340508 173068 340564 189196
rect 339836 157042 339892 157052
rect 339948 173012 340340 173068
rect 340396 173012 340564 173068
rect 341068 220052 341348 220108
rect 339948 154532 340004 173012
rect 339948 154466 340004 154476
rect 340396 153524 340452 173012
rect 341068 156884 341124 220052
rect 341852 162708 341908 356076
rect 341852 162642 341908 162652
rect 341964 352548 342020 352558
rect 341964 161140 342020 352492
rect 342972 340900 343028 340910
rect 342636 299012 342692 299022
rect 342524 277284 342580 277294
rect 342412 268772 342468 268782
rect 341964 161074 342020 161084
rect 342076 256228 342132 256238
rect 341068 156818 341124 156828
rect 340396 151396 340452 153468
rect 340396 151330 340452 151340
rect 342076 151172 342132 256172
rect 342188 248276 342244 248286
rect 342188 237748 342244 248220
rect 342188 237682 342244 237692
rect 342188 201124 342244 201134
rect 342188 163828 342244 201068
rect 342188 163762 342244 163772
rect 342300 198212 342356 198222
rect 342300 162260 342356 198156
rect 342300 162194 342356 162204
rect 342300 157220 342356 157230
rect 342300 156884 342356 157164
rect 342300 156818 342356 156828
rect 342076 151106 342132 151116
rect 342412 150724 342468 268716
rect 342524 248500 342580 277228
rect 342524 248434 342580 248444
rect 342412 150658 342468 150668
rect 342524 247828 342580 247838
rect 342524 95732 342580 247772
rect 342524 95666 342580 95676
rect 342636 48468 342692 298956
rect 342748 263844 342804 263854
rect 342748 239764 342804 263788
rect 342748 239698 342804 239708
rect 342860 249508 342916 249518
rect 342860 236068 342916 249452
rect 342860 236002 342916 236012
rect 342972 157332 343028 340844
rect 343084 268772 343140 365036
rect 343196 291396 343252 389004
rect 343308 387268 343364 387278
rect 343308 292516 343364 387212
rect 343420 379764 343476 379774
rect 343420 293188 343476 379708
rect 343532 372260 343588 393148
rect 345212 385812 345268 407260
rect 345212 385746 345268 385756
rect 345548 384468 345604 384478
rect 343532 372194 343588 372204
rect 345436 381332 345492 381342
rect 345324 365988 345380 365998
rect 345212 357924 345268 357934
rect 343980 342692 344036 342702
rect 343868 341796 343924 341806
rect 343644 340004 343700 340014
rect 343420 293122 343476 293132
rect 343532 339108 343588 339118
rect 343308 292450 343364 292460
rect 343196 291330 343252 291340
rect 343084 268706 343140 268716
rect 343196 272804 343252 272814
rect 343196 237972 343252 272748
rect 343308 271012 343364 271022
rect 343308 239316 343364 270956
rect 343420 267428 343476 267438
rect 343420 239876 343476 267372
rect 343532 250404 343588 339052
rect 343644 264628 343700 339948
rect 343644 264562 343700 264572
rect 343532 250338 343588 250348
rect 343420 239810 343476 239820
rect 343308 239250 343364 239260
rect 343196 237906 343252 237916
rect 343532 238756 343588 238766
rect 342972 157266 343028 157276
rect 342748 157108 342804 157118
rect 342748 150388 342804 157052
rect 342748 150322 342804 150332
rect 342636 48402 342692 48412
rect 339500 46498 339556 46508
rect 339388 43250 339444 43260
rect 338940 43138 338996 43148
rect 338716 42802 338772 42812
rect 338492 41234 338548 41244
rect 343532 41188 343588 238700
rect 343756 238644 343812 238654
rect 343644 209972 343700 209982
rect 343644 107380 343700 209916
rect 343644 107314 343700 107324
rect 343756 41412 343812 238588
rect 343868 157780 343924 341740
rect 343868 157714 343924 157724
rect 343980 157668 344036 342636
rect 344092 273700 344148 273710
rect 344092 238980 344148 273644
rect 344092 238914 344148 238924
rect 344428 254884 344484 254894
rect 344428 238644 344484 254828
rect 344540 252644 344596 252654
rect 344540 245140 344596 252588
rect 344540 245074 344596 245084
rect 344652 245252 344708 245262
rect 344652 240324 344708 245196
rect 344652 240258 344708 240268
rect 344428 238578 344484 238588
rect 344316 208404 344372 208414
rect 343980 157602 344036 157612
rect 344204 177268 344260 177278
rect 344204 157556 344260 177212
rect 344204 157490 344260 157500
rect 344316 156996 344372 208348
rect 344316 156930 344372 156940
rect 345100 195860 345156 195870
rect 345100 149268 345156 195804
rect 345100 149202 345156 149212
rect 345212 147588 345268 357868
rect 345324 163716 345380 365932
rect 345436 358596 345492 381276
rect 345436 358530 345492 358540
rect 345324 163650 345380 163660
rect 345436 348964 345492 348974
rect 345436 158676 345492 348908
rect 345548 309092 345604 384412
rect 345772 383908 345828 383918
rect 345772 366212 345828 383852
rect 345772 366146 345828 366156
rect 346892 380660 346948 380670
rect 346892 329308 346948 380604
rect 347004 377524 347060 410088
rect 348572 410004 348628 410014
rect 348572 382900 348628 409948
rect 351260 409444 351316 409454
rect 351148 409332 351204 409342
rect 348684 407988 348740 407998
rect 348684 385924 348740 407932
rect 350588 407876 350644 407886
rect 350364 407764 350420 407774
rect 348684 385858 348740 385868
rect 350252 404404 350308 404414
rect 348572 382834 348628 382844
rect 350252 382452 350308 404348
rect 350364 387492 350420 407708
rect 350364 387426 350420 387436
rect 350476 400036 350532 400046
rect 350252 382386 350308 382396
rect 350364 384580 350420 384590
rect 347004 377458 347060 377468
rect 348572 370468 348628 370478
rect 346780 329252 346948 329308
rect 347004 359716 347060 359726
rect 347004 329308 347060 359660
rect 347004 329252 347284 329308
rect 346780 328356 346836 329252
rect 346780 325106 346836 328300
rect 347228 325332 347284 329252
rect 346780 325054 346782 325106
rect 346834 325054 346836 325106
rect 346780 325042 346836 325054
rect 347004 325276 347284 325332
rect 345548 309026 345604 309036
rect 346108 314916 346164 314926
rect 345548 299124 345604 299134
rect 345548 257012 345604 299068
rect 345996 283892 346052 283902
rect 345884 282212 345940 282222
rect 345772 262388 345828 262398
rect 345548 256946 345604 256956
rect 345660 258692 345716 258702
rect 345436 158610 345492 158620
rect 345548 197540 345604 197550
rect 345212 147522 345268 147532
rect 345548 139412 345604 197484
rect 345660 154532 345716 258636
rect 345660 154466 345716 154476
rect 345772 150500 345828 262332
rect 345884 154308 345940 282156
rect 345884 154242 345940 154252
rect 345772 150434 345828 150444
rect 345548 139346 345604 139356
rect 345996 48244 346052 283836
rect 346108 157892 346164 314860
rect 346892 308644 346948 308654
rect 346444 285348 346500 285358
rect 346220 255780 346276 255790
rect 346220 240212 346276 255724
rect 346220 240146 346276 240156
rect 346332 248500 346388 248510
rect 346332 161028 346388 248444
rect 346444 246820 346500 285292
rect 346668 276388 346724 276398
rect 346444 246754 346500 246764
rect 346556 250404 346612 250414
rect 346332 160962 346388 160972
rect 346108 157826 346164 157836
rect 346556 157444 346612 250348
rect 346668 229348 346724 276332
rect 346668 229282 346724 229292
rect 346556 157378 346612 157388
rect 346892 50260 346948 308588
rect 347004 147700 347060 325276
rect 347004 147634 347060 147644
rect 347116 325106 347172 325118
rect 347116 325054 347118 325106
rect 347170 325054 347172 325106
rect 347116 116788 347172 325054
rect 347228 280532 347284 280542
rect 347228 159572 347284 280476
rect 348012 273028 348068 273038
rect 348012 267148 348068 272972
rect 347788 267092 348068 267148
rect 347788 245252 347844 267092
rect 347788 245186 347844 245196
rect 347900 262948 347956 262958
rect 347900 240548 347956 262892
rect 348012 253988 348068 253998
rect 348012 241556 348068 253932
rect 348012 241490 348068 241500
rect 347900 240482 347956 240492
rect 347228 159506 347284 159516
rect 347340 197652 347396 197662
rect 347340 148708 347396 197596
rect 348572 165060 348628 370412
rect 350252 364196 350308 364206
rect 348572 164994 348628 165004
rect 348684 362404 348740 362414
rect 348684 162036 348740 362348
rect 348796 354340 348852 354350
rect 348796 164276 348852 354284
rect 349020 346276 349076 346286
rect 348796 164210 348852 164220
rect 348908 345380 348964 345390
rect 348908 162932 348964 345324
rect 349020 165172 349076 346220
rect 349580 270116 349636 270126
rect 349468 260260 349524 260270
rect 349356 246932 349412 246942
rect 349244 244916 349300 244926
rect 349020 165106 349076 165116
rect 349132 238644 349188 238654
rect 348908 162866 348964 162876
rect 348684 161970 348740 161980
rect 347340 148642 347396 148652
rect 347116 116722 347172 116732
rect 349132 102228 349188 238588
rect 349244 162484 349300 244860
rect 349244 162418 349300 162428
rect 349132 102162 349188 102172
rect 349356 101444 349412 246876
rect 349468 240436 349524 260204
rect 349580 252644 349636 270060
rect 349580 252578 349636 252588
rect 349468 240370 349524 240380
rect 350252 164500 350308 364140
rect 350364 312564 350420 384524
rect 350476 382788 350532 399980
rect 350588 387380 350644 407820
rect 351148 407092 351204 409276
rect 351148 406644 351204 407036
rect 351260 406756 351316 409388
rect 351260 406690 351316 406700
rect 351148 406578 351204 406588
rect 352044 406644 352100 406654
rect 350588 387314 350644 387324
rect 351820 389844 351876 389854
rect 350476 382722 350532 382732
rect 350588 383124 350644 383134
rect 350588 370692 350644 383068
rect 350588 370626 350644 370636
rect 350812 381444 350868 381454
rect 350364 312498 350420 312508
rect 350476 358820 350532 358830
rect 350252 164434 350308 164444
rect 350364 247940 350420 247950
rect 349356 101378 349412 101388
rect 346892 50194 346948 50204
rect 350364 50148 350420 247884
rect 350476 164388 350532 358764
rect 350476 164322 350532 164332
rect 350588 355236 350644 355246
rect 350588 162596 350644 355180
rect 350700 348068 350756 348078
rect 350700 164612 350756 348012
rect 350812 248276 350868 381388
rect 350924 380772 350980 380782
rect 350924 334404 350980 380716
rect 351820 346500 351876 389788
rect 351820 346434 351876 346444
rect 351932 370692 351988 370702
rect 350924 334338 350980 334348
rect 351260 284452 351316 284462
rect 351260 278964 351316 284396
rect 350812 248210 350868 248220
rect 350924 252084 350980 252094
rect 350700 164546 350756 164556
rect 350588 162530 350644 162540
rect 350812 151172 350868 151182
rect 350812 149716 350868 151116
rect 350812 146132 350868 149660
rect 350812 146066 350868 146076
rect 350924 110180 350980 252028
rect 350924 110114 350980 110124
rect 351036 249508 351092 249518
rect 351036 104356 351092 249452
rect 351260 236516 351316 278908
rect 351260 236450 351316 236460
rect 351372 264740 351428 264750
rect 351372 234612 351428 264684
rect 351372 234546 351428 234556
rect 351484 264628 351540 264638
rect 351484 208404 351540 264572
rect 351820 261268 351876 261278
rect 351820 257012 351876 261212
rect 351820 256946 351876 256956
rect 351820 245252 351876 245262
rect 351820 239540 351876 245196
rect 351820 239474 351876 239484
rect 351484 208338 351540 208348
rect 351148 200788 351204 200798
rect 351148 171332 351204 200732
rect 351148 170436 351204 171276
rect 351148 170370 351204 170380
rect 351260 196420 351316 196430
rect 351260 195300 351316 196364
rect 351260 167748 351316 195244
rect 351260 167682 351316 167692
rect 351932 154420 351988 370636
rect 352044 261828 352100 406588
rect 352156 382788 352212 410088
rect 355516 408100 355572 408110
rect 353724 407652 353780 407662
rect 352716 407204 352772 407214
rect 352156 381444 352212 382732
rect 352156 381378 352212 381388
rect 352268 406756 352324 406766
rect 352156 380548 352212 380558
rect 352156 352548 352212 380492
rect 352156 352482 352212 352492
rect 352268 268772 352324 406700
rect 352604 404964 352660 404974
rect 352604 388836 352660 404908
rect 352380 384804 352436 384814
rect 352380 340452 352436 384748
rect 352380 340386 352436 340396
rect 352492 377524 352548 377534
rect 352380 312564 352436 312574
rect 352380 310212 352436 312508
rect 352380 310146 352436 310156
rect 352380 309092 352436 309102
rect 352380 304164 352436 309036
rect 352380 304098 352436 304108
rect 352268 268706 352324 268716
rect 352380 267202 352436 267214
rect 352380 267150 352382 267202
rect 352434 267150 352436 267202
rect 352380 267148 352436 267150
rect 352044 261762 352100 261772
rect 352156 267092 352436 267148
rect 352156 233492 352212 267092
rect 352156 233426 352212 233436
rect 352380 257012 352436 257022
rect 352380 255780 352436 256956
rect 352044 225540 352100 225550
rect 352044 181412 352100 225484
rect 352044 181346 352100 181356
rect 352156 219492 352212 219502
rect 352156 179788 352212 219436
rect 352044 179732 352212 179788
rect 352268 207396 352324 207406
rect 352044 178500 352100 179732
rect 352044 163940 352100 178444
rect 352268 173684 352324 207340
rect 352380 198212 352436 255724
rect 352380 198146 352436 198156
rect 352492 179788 352548 377468
rect 352268 173124 352324 173628
rect 352268 173058 352324 173068
rect 352380 179732 352548 179788
rect 352380 172900 352436 179732
rect 352044 163874 352100 163884
rect 352268 172844 352436 172900
rect 351932 154354 351988 154364
rect 352268 153076 352324 172844
rect 352380 171332 352436 171342
rect 352380 165396 352436 171276
rect 352604 168028 352660 388780
rect 352716 245252 352772 407148
rect 353612 404516 353668 404526
rect 353612 382228 353668 404460
rect 353724 385700 353780 407596
rect 355180 407540 355236 407550
rect 353724 385634 353780 385644
rect 353836 399588 353892 399598
rect 353836 382564 353892 399532
rect 354844 397460 354900 397470
rect 354732 394212 354788 394222
rect 354060 393988 354116 393998
rect 354060 382676 354116 393932
rect 354732 387940 354788 394156
rect 354844 390964 354900 397404
rect 354956 397348 355012 397358
rect 354956 391188 355012 397292
rect 355068 397124 355124 397134
rect 355068 394212 355124 397068
rect 355068 394146 355124 394156
rect 355180 393988 355236 407484
rect 355404 406532 355460 406542
rect 355292 403060 355348 403070
rect 355292 398132 355348 403004
rect 355292 398066 355348 398076
rect 355404 397908 355460 406476
rect 354956 391122 355012 391132
rect 355068 393932 355236 393988
rect 355292 397852 355460 397908
rect 354844 390898 354900 390908
rect 355068 390740 355124 393932
rect 355180 393764 355236 393774
rect 355180 392644 355236 393708
rect 355180 392578 355236 392588
rect 355068 390674 355124 390684
rect 354732 387874 354788 387884
rect 354060 382610 354116 382620
rect 353836 382498 353892 382508
rect 355292 382340 355348 397852
rect 355404 397236 355460 397246
rect 355404 387828 355460 397180
rect 355516 390628 355572 408044
rect 357308 404964 357364 410088
rect 362460 407316 362516 410088
rect 367612 408212 367668 410088
rect 367612 408146 367668 408156
rect 372764 408100 372820 410088
rect 372764 408034 372820 408044
rect 377916 407988 377972 410088
rect 379596 408660 379652 408670
rect 379596 408212 379652 408604
rect 379596 408146 379652 408156
rect 377916 407922 377972 407932
rect 383068 407540 383124 410088
rect 383068 407474 383124 407484
rect 383292 407540 383348 407550
rect 362460 407250 362516 407260
rect 357308 404898 357364 404908
rect 383292 399812 383348 407484
rect 388220 404852 388276 410088
rect 393372 407652 393428 410088
rect 398524 407876 398580 410088
rect 398524 407810 398580 407820
rect 399756 407876 399812 407886
rect 393372 407586 393428 407596
rect 397292 407652 397348 407662
rect 388220 404786 388276 404796
rect 383292 399746 383348 399756
rect 371980 397460 372036 397470
rect 361228 396788 361284 396798
rect 361228 395220 361284 396732
rect 361228 395154 361284 395164
rect 358204 395108 358260 395118
rect 358204 394996 358260 395052
rect 365148 395108 365204 395118
rect 365148 394996 365204 395052
rect 371980 394996 372036 397404
rect 386428 397348 386484 397358
rect 379820 395108 379876 395118
rect 379820 394996 379876 395052
rect 358204 394940 358904 394996
rect 365148 394940 365848 394996
rect 371980 394940 372792 394996
rect 379736 394940 379876 394996
rect 386428 394996 386484 397292
rect 393148 397236 393204 397246
rect 393148 394996 393204 397180
rect 397292 396340 397348 407596
rect 399756 404740 399812 407820
rect 403676 407428 403732 410088
rect 408828 407764 408884 410088
rect 408828 407698 408884 407708
rect 403676 407362 403732 407372
rect 403900 407428 403956 407438
rect 399756 404674 399812 404684
rect 403900 402948 403956 407372
rect 413980 406532 414036 410088
rect 419132 407876 419188 410088
rect 419132 407810 419188 407820
rect 413980 406466 414036 406476
rect 419356 407764 419412 407774
rect 403900 402882 403956 402892
rect 414092 399924 414148 399934
rect 414092 397460 414148 399868
rect 414092 397394 414148 397404
rect 406812 397124 406868 397134
rect 397292 396274 397348 396284
rect 400204 397012 400260 397022
rect 400204 394996 400260 396956
rect 403116 396564 403172 396574
rect 386428 394940 386680 394996
rect 393148 394940 393624 394996
rect 400204 394940 400568 394996
rect 403116 394772 403172 396508
rect 406812 394996 406868 397068
rect 413756 396564 413812 396574
rect 413756 394996 413812 396508
rect 419356 396228 419412 407708
rect 424284 407428 424340 410088
rect 429436 407540 429492 410088
rect 430108 408436 430164 408446
rect 430108 408100 430164 408380
rect 430108 408034 430164 408044
rect 429436 407474 429492 407484
rect 424284 407362 424340 407372
rect 424956 407428 425012 407438
rect 421596 401716 421652 401726
rect 421596 397348 421652 401660
rect 424956 399700 425012 407372
rect 434588 404628 434644 410088
rect 439740 408212 439796 410088
rect 439740 408146 439796 408156
rect 444892 407876 444948 410088
rect 444892 407810 444948 407820
rect 450044 407652 450100 410088
rect 455196 407764 455252 410088
rect 455196 407698 455252 407708
rect 450044 407586 450100 407596
rect 434588 404562 434644 404572
rect 445116 407540 445172 407550
rect 424956 399634 425012 399644
rect 442092 400036 442148 400046
rect 421596 397282 421652 397292
rect 427644 397460 427700 397470
rect 419356 396162 419412 396172
rect 420700 396900 420756 396910
rect 420700 394996 420756 396844
rect 427644 394996 427700 397404
rect 435148 397348 435204 397358
rect 429212 396900 429268 396910
rect 406812 394940 407512 394996
rect 413756 394940 414456 394996
rect 420700 394940 421400 394996
rect 427644 394940 428344 394996
rect 403116 394706 403172 394716
rect 429212 394660 429268 396844
rect 435148 394996 435204 397292
rect 442092 394996 442148 399980
rect 445116 399476 445172 407484
rect 445116 399410 445172 399420
rect 448588 396900 448644 396910
rect 448588 394996 448644 396844
rect 455308 396564 455364 396574
rect 455308 394996 455364 396508
rect 460348 396004 460404 410088
rect 460348 395938 460404 395948
rect 464492 406644 464548 406654
rect 464492 395892 464548 406588
rect 465500 406644 465556 410088
rect 465500 406578 465556 406588
rect 464492 395826 464548 395836
rect 466172 406084 466228 406094
rect 466172 395892 466228 406028
rect 466172 395826 466228 395836
rect 469196 398244 469252 398254
rect 469196 394996 469252 398188
rect 470652 395780 470708 410088
rect 472892 406644 472948 406654
rect 472892 403060 472948 406588
rect 472892 402994 472948 403004
rect 470652 395714 470708 395724
rect 475804 395668 475860 410088
rect 480956 404292 481012 410088
rect 486108 408100 486164 410088
rect 486108 408034 486164 408044
rect 490588 410060 491288 410116
rect 490588 406756 490644 410060
rect 496412 407652 496468 410088
rect 496412 407586 496468 407596
rect 501564 407540 501620 410088
rect 501564 407474 501620 407484
rect 504700 408324 504756 408334
rect 490588 406690 490644 406700
rect 480956 404226 481012 404236
rect 475804 395602 475860 395612
rect 497644 401604 497700 401614
rect 497644 394996 497700 401548
rect 504700 396508 504756 408268
rect 506716 399588 506772 410088
rect 511868 410050 511924 410060
rect 517020 407428 517076 410088
rect 522172 407540 522228 410088
rect 522172 407474 522228 407484
rect 527324 407540 527380 410088
rect 527324 407474 527380 407484
rect 517020 407362 517076 407372
rect 529340 402836 529396 526764
rect 529340 402770 529396 402780
rect 529452 489188 529508 489198
rect 529452 401380 529508 489132
rect 529564 479892 529620 479902
rect 529564 402500 529620 479836
rect 529564 402434 529620 402444
rect 529676 470484 529732 470494
rect 529452 401314 529508 401324
rect 506716 399522 506772 399532
rect 529676 399364 529732 470428
rect 529788 409332 529844 590604
rect 540540 575540 540596 595560
rect 562604 590548 562660 595560
rect 562604 590482 562660 590492
rect 584668 590212 584724 595560
rect 584668 590146 584724 590156
rect 540540 575474 540596 575484
rect 537628 546308 537684 546318
rect 532588 541604 532644 541614
rect 530908 513380 530964 513390
rect 529788 409266 529844 409276
rect 529900 465668 529956 465678
rect 529676 399298 529732 399308
rect 529900 399252 529956 465612
rect 529900 399186 529956 399196
rect 530012 460852 530068 460862
rect 530012 399140 530068 460796
rect 530012 399074 530068 399084
rect 530124 414596 530180 414606
rect 530124 399028 530180 414540
rect 530124 398962 530180 398972
rect 518028 396788 518084 396798
rect 504700 396452 504868 396508
rect 504812 394996 504868 396452
rect 435148 394940 435288 394996
rect 442092 394940 442232 394996
rect 448588 394940 449176 394996
rect 455308 394940 456120 394996
rect 469196 394940 470008 394996
rect 483858 394940 483868 394996
rect 483924 394940 483934 394996
rect 497644 394940 497784 394996
rect 504728 394940 504868 394996
rect 518028 394996 518084 396732
rect 518028 394940 518616 394996
rect 525522 394940 525532 394996
rect 525588 394940 525598 394996
rect 490812 394884 490868 394894
rect 490812 394818 490868 394828
rect 476924 394772 476980 394782
rect 476924 394706 476980 394716
rect 511644 394772 511700 394782
rect 511644 394706 511700 394716
rect 429212 394594 429268 394604
rect 463036 394660 463092 394670
rect 463036 394594 463092 394604
rect 530908 394548 530964 513324
rect 531020 452228 531076 452238
rect 531020 405972 531076 452172
rect 531244 424004 531300 424014
rect 531020 405906 531076 405916
rect 531132 419300 531188 419310
rect 531132 400708 531188 419244
rect 531244 405748 531300 423948
rect 531244 405682 531300 405692
rect 532588 404180 532644 541548
rect 534268 536900 534324 536910
rect 532700 456932 532756 456942
rect 532700 409220 532756 456876
rect 532700 409154 532756 409164
rect 532812 447524 532868 447534
rect 532812 404404 532868 447468
rect 532924 438116 532980 438126
rect 532924 404516 532980 438060
rect 533036 433412 533092 433422
rect 533036 405860 533092 433356
rect 534268 406308 534324 536844
rect 534380 532196 534436 532206
rect 534380 409108 534436 532140
rect 535948 522788 536004 522798
rect 534380 409042 534436 409052
rect 534492 503972 534548 503982
rect 534268 406242 534324 406252
rect 533036 405794 533092 405804
rect 532924 404450 532980 404460
rect 532812 404338 532868 404348
rect 532588 404114 532644 404124
rect 534492 401268 534548 503916
rect 534492 401202 534548 401212
rect 534604 494564 534660 494574
rect 534604 401044 534660 494508
rect 534604 400978 534660 400988
rect 534716 485156 534772 485166
rect 534716 400820 534772 485100
rect 535948 402724 536004 522732
rect 535948 402658 536004 402668
rect 536060 518084 536116 518094
rect 536060 402612 536116 518028
rect 536060 402546 536116 402556
rect 536172 508676 536228 508686
rect 536172 401156 536228 508620
rect 536172 401090 536228 401100
rect 536284 499268 536340 499278
rect 536284 400932 536340 499212
rect 537628 406196 537684 546252
rect 545132 482916 545188 482926
rect 537628 406130 537684 406140
rect 540092 456484 540148 456494
rect 540092 402388 540148 456428
rect 545132 409892 545188 482860
rect 587132 443268 587188 443278
rect 545132 409826 545188 409836
rect 560252 410004 560308 410014
rect 540092 402322 540148 402332
rect 536284 400866 536340 400876
rect 534716 400754 534772 400764
rect 531132 400642 531188 400652
rect 539308 397796 539364 397806
rect 531804 396676 531860 396686
rect 531804 394996 531860 396620
rect 539308 394996 539364 397740
rect 546252 396900 546308 396910
rect 546252 394996 546308 396844
rect 553196 396676 553252 396686
rect 553196 394996 553252 396620
rect 560252 396508 560308 409948
rect 587132 406644 587188 443212
rect 587132 406578 587188 406588
rect 583884 404068 583940 404078
rect 583772 403284 583828 403294
rect 574028 396900 574084 396910
rect 567084 396564 567140 396574
rect 560252 396452 560420 396508
rect 560364 394996 560420 396452
rect 531804 394940 532504 394996
rect 539308 394940 539448 394996
rect 546252 394940 546392 394996
rect 553196 394940 553336 394996
rect 560280 394940 560420 394996
rect 567084 394996 567140 396508
rect 574028 394996 574084 396844
rect 580972 396788 581028 396798
rect 580972 394996 581028 396732
rect 582988 395892 583044 395902
rect 567084 394940 567224 394996
rect 574028 394940 574168 394996
rect 580972 394940 581112 394996
rect 582988 394884 583044 395836
rect 582988 394818 583044 394828
rect 583660 394884 583716 394894
rect 530908 394482 530964 394492
rect 355516 390562 355572 390572
rect 355404 387762 355460 387772
rect 355292 382274 355348 382284
rect 353612 382162 353668 382172
rect 353612 366884 353668 366894
rect 353500 310212 353556 310222
rect 352716 245186 352772 245196
rect 352828 272132 352884 272142
rect 352828 238644 352884 272076
rect 352828 238578 352884 238588
rect 353500 236852 353556 310156
rect 353500 236786 353556 236796
rect 352716 213444 352772 213454
rect 352716 175812 352772 213388
rect 352716 175746 352772 175756
rect 353500 173908 353556 173918
rect 352380 165330 352436 165340
rect 352492 167972 352660 168028
rect 352716 171108 352772 171118
rect 352492 162372 352548 167972
rect 352604 162372 352660 162382
rect 352492 162316 352604 162372
rect 352604 162306 352660 162316
rect 352604 154420 352660 154430
rect 352604 153748 352660 154364
rect 352604 153682 352660 153692
rect 352268 149548 352324 153020
rect 352268 149492 352436 149548
rect 352380 145572 352436 149492
rect 352380 145506 352436 145516
rect 351036 104290 351092 104300
rect 351148 58772 351204 58782
rect 351148 57204 351204 58716
rect 352716 58772 352772 171052
rect 353500 165620 353556 173852
rect 353500 165554 353556 165564
rect 353612 156212 353668 366828
rect 355404 361508 355460 361518
rect 353612 156146 353668 156156
rect 353724 353444 353780 353454
rect 353724 147252 353780 353388
rect 355292 351652 355348 351662
rect 353836 349860 353892 349870
rect 353836 161028 353892 349804
rect 354508 338212 354564 338222
rect 354060 317044 354116 317054
rect 353948 298116 354004 298126
rect 353948 272132 354004 298060
rect 353948 272066 354004 272076
rect 353836 160962 353892 160972
rect 353948 252084 354004 252094
rect 353724 147186 353780 147196
rect 353948 99092 354004 252028
rect 354060 234500 354116 316988
rect 354396 284788 354452 284798
rect 354284 273924 354340 273934
rect 354284 267202 354340 273868
rect 354284 267150 354286 267202
rect 354338 267150 354340 267202
rect 354060 234164 354116 234444
rect 354060 234098 354116 234108
rect 354172 238644 354228 238654
rect 354060 183316 354116 183326
rect 354060 159572 354116 183260
rect 354172 173908 354228 238588
rect 354172 173842 354228 173852
rect 354172 173684 354228 173694
rect 354172 165284 354228 173628
rect 354172 165218 354228 165228
rect 354284 164052 354340 267150
rect 354284 163986 354340 163996
rect 354060 159506 354116 159516
rect 354396 107268 354452 284732
rect 354508 177268 354564 338156
rect 354620 287364 354676 287374
rect 354620 234388 354676 287308
rect 355068 279412 355124 279422
rect 355068 238308 355124 279356
rect 355068 238242 355124 238252
rect 354620 234322 354676 234332
rect 354620 234164 354676 234174
rect 354620 231868 354676 234108
rect 354620 231812 354788 231868
rect 354508 177202 354564 177212
rect 354732 166292 354788 231812
rect 354732 166226 354788 166236
rect 355180 183428 355236 183438
rect 354396 107202 354452 107212
rect 353948 99026 354004 99036
rect 352716 58706 352772 58716
rect 351148 52948 351204 57148
rect 351148 52882 351204 52892
rect 350364 50082 350420 50092
rect 345996 48178 346052 48188
rect 355180 45220 355236 183372
rect 355292 147140 355348 351596
rect 355404 161252 355460 361452
rect 355404 161186 355460 161196
rect 355516 238308 355572 238318
rect 355516 155316 355572 238252
rect 486444 165620 486500 165630
rect 422716 165396 422772 165406
rect 365820 165172 365876 165182
rect 365820 165106 365876 165116
rect 358204 165004 358904 165060
rect 372092 165004 372792 165060
rect 379736 165004 379876 165060
rect 358204 162932 358260 165004
rect 358204 162866 358260 162876
rect 372092 162484 372148 165004
rect 379820 164612 379876 165004
rect 379820 164546 379876 164556
rect 386540 165004 386680 165060
rect 393484 165004 393624 165060
rect 399868 165004 400568 165060
rect 407372 165004 407512 165060
rect 414316 165004 414456 165060
rect 421260 165004 421400 165060
rect 372092 162418 372148 162428
rect 386540 158676 386596 165004
rect 393484 161028 393540 165004
rect 399868 164164 399924 165004
rect 399868 164098 399924 164108
rect 407372 161308 407428 165004
rect 407372 161252 407540 161308
rect 393484 160962 393540 160972
rect 386540 158610 386596 158620
rect 355516 155250 355572 155260
rect 366268 155316 366324 155326
rect 355292 147074 355348 147084
rect 366268 145908 366324 155260
rect 407484 147140 407540 161252
rect 414316 161140 414372 165004
rect 414316 161074 414372 161084
rect 420812 164724 420868 164734
rect 420812 154308 420868 164668
rect 421260 161308 421316 165004
rect 421820 163940 421876 163950
rect 421260 161252 421428 161308
rect 420812 154242 420868 154252
rect 421372 147252 421428 161252
rect 421820 153972 421876 163884
rect 421820 149548 421876 153916
rect 422492 156996 422548 157006
rect 422492 154308 422548 156940
rect 421820 149492 422324 149548
rect 421372 147186 421428 147196
rect 407484 147074 407540 147084
rect 366268 93492 366324 145852
rect 401884 147028 401940 147038
rect 400316 145348 400372 145358
rect 386092 107380 386148 107390
rect 376572 104132 376628 104142
rect 372988 103796 373044 103806
rect 372988 99988 373044 103740
rect 374668 103236 374724 103246
rect 374668 99988 374724 103180
rect 376572 99988 376628 104076
rect 383964 104020 384020 104030
rect 381388 103908 381444 103918
rect 378028 103684 378084 103694
rect 378028 99988 378084 103628
rect 379708 103348 379764 103358
rect 379708 99988 379764 103292
rect 381388 99988 381444 103852
rect 383180 103572 383236 103582
rect 383180 99988 383236 103516
rect 372988 99932 373688 99988
rect 374668 99932 375256 99988
rect 376572 99932 376824 99988
rect 378028 99932 378392 99988
rect 379708 99932 379960 99988
rect 381388 99932 381528 99988
rect 383096 99932 383236 99988
rect 383964 99988 384020 103964
rect 386092 99988 386148 107324
rect 390796 107044 390852 107054
rect 387100 103460 387156 103470
rect 387100 99988 387156 103404
rect 389228 103236 389284 103246
rect 389228 99988 389284 103180
rect 390796 99988 390852 106988
rect 393932 106932 393988 106942
rect 392364 103348 392420 103358
rect 392364 99988 392420 103292
rect 393932 99988 393988 106876
rect 395500 106820 395556 106830
rect 395500 99988 395556 106764
rect 396508 104132 396564 104142
rect 396508 99988 396564 104076
rect 398188 104132 398244 104142
rect 398188 99988 398244 104076
rect 400316 102508 400372 145292
rect 401884 102508 401940 146972
rect 421820 144676 421876 144686
rect 421708 144564 421764 144574
rect 406588 138628 406644 138638
rect 403452 133588 403508 133598
rect 403452 102508 403508 133532
rect 406588 114268 406644 138572
rect 415996 135268 416052 135278
rect 408156 132020 408212 132030
rect 406588 114212 406756 114268
rect 400204 102452 400372 102508
rect 401772 102452 401940 102508
rect 403340 102452 403508 102508
rect 404908 106708 404964 106718
rect 400204 99988 400260 102452
rect 401772 99988 401828 102452
rect 403340 99988 403396 102452
rect 404908 99988 404964 106652
rect 406588 105028 406644 105038
rect 406588 102564 406644 104972
rect 406588 102498 406644 102508
rect 406700 99988 406756 114212
rect 408156 102508 408212 131964
rect 414428 131908 414484 131918
rect 411292 125188 411348 125198
rect 383964 99932 384664 99988
rect 386092 99932 386232 99988
rect 387100 99932 387800 99988
rect 389228 99932 389368 99988
rect 390796 99932 390936 99988
rect 392364 99932 392504 99988
rect 393932 99932 394072 99988
rect 395500 99932 395640 99988
rect 396508 99932 397208 99988
rect 398188 99932 398776 99988
rect 400204 99932 400344 99988
rect 401772 99932 401912 99988
rect 403340 99932 403480 99988
rect 404908 99932 405048 99988
rect 406616 99932 406756 99988
rect 408044 102452 408212 102508
rect 408940 102564 408996 102574
rect 411292 102508 411348 125132
rect 412860 115108 412916 115118
rect 412860 102508 412916 115052
rect 414428 102508 414484 131852
rect 415996 102508 416052 135212
rect 408044 99988 408100 102452
rect 408940 99988 408996 102508
rect 411180 102452 411348 102508
rect 412748 102452 412916 102508
rect 414316 102452 414484 102508
rect 415884 102452 416052 102508
rect 411180 99988 411236 102452
rect 412748 99988 412804 102452
rect 414316 99988 414372 102452
rect 415884 99988 415940 102452
rect 408044 99932 408184 99988
rect 408940 99932 409752 99988
rect 411180 99932 411320 99988
rect 412748 99932 412888 99988
rect 414316 99932 414456 99988
rect 415884 99932 416024 99988
rect 366268 91476 366324 93436
rect 366268 91410 366324 91420
rect 420028 81620 420084 81630
rect 367836 58324 367892 58334
rect 367836 57204 367892 58268
rect 367836 53284 367892 57148
rect 367836 53228 368004 53284
rect 367948 51044 368004 53228
rect 367948 50978 368004 50988
rect 419356 52164 419412 52174
rect 419356 49812 419412 52108
rect 419356 49746 419412 49756
rect 420028 48132 420084 81564
rect 420028 48066 420084 48076
rect 420140 77364 420196 77374
rect 420140 48020 420196 77308
rect 421708 77364 421764 144508
rect 421820 82292 421876 144620
rect 421932 122612 421988 122622
rect 421932 87220 421988 122556
rect 421932 87154 421988 87164
rect 421820 82226 421876 82236
rect 421708 77298 421764 77308
rect 420252 72436 420308 72446
rect 420252 50036 420308 72380
rect 422268 72436 422324 149492
rect 422268 72370 422324 72380
rect 421932 68852 421988 68862
rect 421932 67508 421988 68796
rect 420252 49970 420308 49980
rect 420364 62580 420420 62590
rect 420364 49924 420420 62524
rect 420364 49858 420420 49868
rect 421708 57652 421764 57662
rect 421708 49588 421764 57596
rect 421932 49700 421988 67452
rect 422492 52724 422548 154252
rect 422716 154196 422772 165340
rect 466172 165396 466228 165406
rect 422716 57652 422772 154140
rect 422940 165284 422996 165294
rect 422940 154084 422996 165228
rect 427644 165004 428344 165060
rect 435148 165004 435288 165060
rect 441868 165004 442232 165060
rect 448588 165004 449176 165060
rect 455980 165004 456120 165060
rect 462364 165004 463064 165060
rect 422940 62580 422996 154028
rect 423164 164948 423220 164958
rect 423164 154420 423220 164892
rect 427644 164276 427700 165004
rect 427644 164210 427700 164220
rect 435148 162596 435204 165004
rect 441868 162708 441924 165004
rect 448588 162820 448644 165004
rect 448588 162754 448644 162764
rect 441868 162642 441924 162652
rect 435148 162530 435204 162540
rect 455980 161308 456036 165004
rect 462364 164388 462420 165004
rect 462364 164322 462420 164332
rect 464940 164164 464996 164174
rect 463596 163940 463652 163950
rect 458220 162484 458276 162494
rect 457772 161364 457828 161374
rect 455980 161252 456148 161308
rect 423164 68852 423220 154364
rect 456092 147588 456148 161252
rect 456092 147522 456148 147532
rect 457772 137732 457828 161308
rect 458108 159908 458164 159918
rect 457884 159684 457940 159694
rect 457884 139188 457940 159628
rect 457996 158004 458052 158014
rect 457996 141092 458052 157948
rect 458108 146132 458164 159852
rect 458220 147700 458276 162428
rect 459452 154644 459508 154654
rect 458220 147634 458276 147644
rect 458556 148372 458612 148382
rect 458108 146066 458164 146076
rect 458556 142660 458612 148316
rect 458556 142594 458612 142604
rect 457996 141026 458052 141036
rect 459452 139412 459508 154588
rect 463596 154308 463652 163884
rect 463596 149912 463652 154252
rect 464940 154196 464996 164108
rect 466172 161308 466228 165340
rect 469308 165004 470008 165060
rect 476952 165004 477092 165060
rect 483896 165004 484036 165060
rect 469308 162484 469364 165004
rect 477036 162932 477092 165004
rect 477036 162866 477092 162876
rect 481068 164052 481124 164062
rect 469308 162418 469364 162428
rect 464940 149912 464996 154140
rect 466060 161252 466228 161308
rect 466060 154084 466116 161252
rect 479724 159908 479780 159918
rect 470316 157892 470372 157902
rect 466060 149828 466116 154028
rect 467628 154420 467684 154430
rect 467628 149912 467684 154364
rect 468972 153972 469028 153982
rect 468972 149912 469028 153916
rect 470316 153972 470372 157836
rect 473788 156996 473844 157006
rect 473004 154756 473060 154766
rect 470316 153906 470372 153916
rect 471660 153972 471716 153982
rect 470316 152964 470372 152974
rect 466060 149772 466312 149828
rect 470316 149716 470372 152908
rect 471660 151396 471716 153916
rect 471660 149912 471716 151340
rect 473004 149912 473060 154700
rect 473788 152964 473844 156940
rect 473788 152898 473844 152908
rect 474348 156324 474404 156334
rect 474348 149912 474404 156268
rect 475692 152964 475748 152974
rect 475692 149912 475748 152908
rect 478380 151284 478436 151294
rect 477036 149940 477092 149950
rect 478380 149912 478436 151228
rect 479724 149912 479780 159852
rect 481068 149912 481124 163996
rect 483980 161252 484036 165004
rect 483980 161186 484036 161196
rect 482412 158116 482468 158126
rect 482412 149912 482468 158060
rect 483756 154532 483812 154542
rect 483756 149912 483812 154476
rect 485100 152964 485156 152974
rect 485100 149912 485156 152908
rect 486444 149912 486500 165564
rect 557900 165508 557956 165518
rect 490700 165004 490840 165060
rect 497784 165004 497924 165060
rect 490700 162036 490756 165004
rect 490700 161970 490756 161980
rect 495852 163268 495908 163278
rect 487788 154532 487844 154542
rect 487788 149912 487844 154476
rect 488908 154532 488964 154542
rect 488908 149940 488964 154476
rect 490476 154532 490532 154542
rect 488908 149884 489160 149940
rect 490476 149912 490532 154476
rect 491820 154532 491876 154542
rect 491820 149912 491876 154476
rect 493164 154532 493220 154542
rect 493164 149912 493220 154476
rect 494732 153300 494788 153310
rect 494508 152964 494564 152974
rect 494508 149912 494564 152908
rect 477036 149874 477092 149884
rect 470316 149650 470372 149660
rect 494732 149716 494788 153244
rect 495852 149912 495908 163212
rect 497868 162932 497924 165004
rect 504028 165004 504728 165060
rect 511532 165004 511672 165060
rect 517916 165004 518616 165060
rect 525420 165004 525560 165060
rect 532364 165004 532504 165060
rect 539308 165004 539448 165060
rect 546392 165004 546532 165060
rect 553298 165004 553308 165060
rect 553364 165004 553374 165060
rect 504028 164500 504084 165004
rect 504028 164434 504084 164444
rect 497868 162866 497924 162876
rect 502796 162372 502852 162382
rect 497196 161700 497252 161710
rect 497196 149912 497252 161644
rect 502796 154532 502852 162316
rect 508732 160244 508788 160254
rect 502796 154466 502852 154476
rect 506604 154532 506660 154542
rect 500108 154084 500164 154094
rect 497308 153636 497364 153646
rect 497308 152740 497364 153580
rect 497308 152674 497364 152684
rect 498540 152964 498596 152974
rect 498540 149912 498596 152908
rect 499884 152964 499940 152974
rect 499884 149912 499940 152908
rect 494732 149650 494788 149660
rect 500108 149716 500164 154028
rect 501228 153860 501284 153870
rect 500668 153412 500724 153422
rect 500668 150948 500724 153356
rect 500668 150882 500724 150892
rect 501228 149912 501284 153804
rect 502572 153748 502628 153758
rect 502572 149912 502628 153692
rect 505260 153524 505316 153534
rect 503916 153076 503972 153086
rect 503916 149912 503972 153020
rect 505260 149912 505316 153468
rect 505596 152964 505652 152974
rect 505596 152628 505652 152908
rect 505596 152562 505652 152572
rect 506604 149912 506660 154476
rect 508732 154532 508788 160188
rect 510748 155988 510804 155998
rect 508732 154466 508788 154476
rect 510636 155876 510692 155886
rect 509292 153636 509348 153646
rect 507276 153524 507332 153534
rect 507276 150836 507332 153468
rect 507276 150770 507332 150780
rect 507948 152292 508004 152302
rect 507948 149912 508004 152236
rect 509292 149912 509348 153580
rect 510636 149912 510692 155820
rect 510748 153748 510804 155932
rect 510748 153682 510804 153692
rect 511532 150724 511588 165004
rect 517916 163716 517972 165004
rect 517916 163650 517972 163660
rect 520044 162148 520100 162158
rect 516012 160692 516068 160702
rect 514668 160356 514724 160366
rect 513324 160132 513380 160142
rect 511532 150658 511588 150668
rect 511980 154532 512036 154542
rect 511980 149912 512036 154476
rect 513324 149912 513380 160076
rect 514668 149912 514724 160300
rect 516012 149912 516068 160636
rect 518700 153300 518756 153310
rect 517356 152180 517412 152190
rect 517356 149912 517412 152124
rect 518700 149912 518756 153244
rect 520044 149912 520100 162092
rect 522508 159460 522564 159470
rect 522508 153860 522564 159404
rect 525420 156212 525476 165004
rect 532364 162932 532420 165004
rect 532364 162866 532420 162876
rect 539308 162932 539364 165004
rect 539308 162866 539364 162876
rect 546476 162932 546532 165004
rect 546476 162866 546532 162876
rect 557004 164724 557060 164734
rect 554652 162260 554708 162270
rect 540876 160580 540932 160590
rect 525420 156146 525476 156156
rect 532588 159348 532644 159358
rect 525420 155764 525476 155774
rect 522508 153794 522564 153804
rect 524076 154084 524132 154094
rect 522732 153412 522788 153422
rect 520828 153300 520884 153310
rect 520828 151060 520884 153244
rect 520828 150994 520884 151004
rect 521388 152964 521444 152974
rect 521388 149912 521444 152908
rect 522732 149912 522788 153356
rect 524076 149912 524132 154028
rect 524188 152964 524244 152974
rect 524188 150276 524244 152908
rect 524188 150210 524244 150220
rect 525420 149912 525476 155708
rect 528108 155652 528164 155662
rect 526764 153748 526820 153758
rect 526764 149912 526820 153692
rect 528108 149912 528164 155596
rect 529452 155540 529508 155550
rect 529452 149912 529508 155484
rect 532588 154532 532644 159292
rect 535948 159236 536004 159246
rect 532588 154466 532644 154476
rect 534828 155428 534884 155438
rect 530796 153300 530852 153310
rect 530796 149912 530852 153244
rect 533484 153076 533540 153086
rect 532140 152964 532196 152974
rect 532140 149912 532196 152908
rect 533484 149912 533540 153020
rect 534828 149912 534884 155372
rect 535948 154420 536004 159180
rect 539196 159124 539252 159134
rect 535948 154354 536004 154364
rect 538860 154532 538916 154542
rect 537516 153860 537572 153870
rect 536172 153524 536228 153534
rect 536172 149912 536228 153468
rect 537516 149912 537572 153804
rect 538860 149912 538916 154476
rect 539196 154308 539252 159068
rect 539196 154242 539252 154252
rect 540204 154420 540260 154430
rect 540204 149912 540260 154364
rect 540876 153748 540932 160524
rect 550956 160468 551012 160478
rect 544236 159012 544292 159022
rect 542892 158900 542948 158910
rect 540876 153682 540932 153692
rect 541548 154308 541604 154318
rect 541548 149912 541604 154252
rect 542892 149912 542948 158844
rect 544236 149912 544292 158956
rect 548268 158788 548324 158798
rect 545580 152068 545636 152078
rect 545580 149912 545636 152012
rect 548268 149912 548324 158732
rect 549612 153748 549668 153758
rect 549612 149912 549668 153692
rect 550956 149912 551012 160412
rect 554540 157780 554596 157790
rect 554428 150388 554484 150398
rect 500108 149650 500164 149660
rect 546924 149604 546980 149614
rect 546924 149538 546980 149548
rect 459452 139346 459508 139356
rect 457884 139122 457940 139132
rect 457772 137666 457828 137676
rect 554428 131012 554484 150332
rect 554540 140532 554596 157724
rect 554540 140466 554596 140476
rect 554428 130946 554484 130956
rect 554652 125972 554708 162204
rect 556892 161476 556948 161486
rect 555100 161364 555156 161374
rect 554988 158004 555044 158014
rect 554876 148708 554932 148718
rect 554652 125906 554708 125916
rect 554764 148372 554820 148382
rect 554764 112196 554820 148316
rect 554876 120260 554932 148652
rect 554876 120194 554932 120204
rect 554764 112130 554820 112140
rect 554988 108836 555044 157948
rect 555100 113204 555156 161308
rect 556332 159684 556388 159694
rect 555212 157668 555268 157678
rect 555212 141428 555268 157612
rect 556220 157332 556276 157342
rect 555212 141362 555268 141372
rect 556108 157220 556164 157230
rect 556108 132020 556164 157164
rect 556220 138292 556276 157276
rect 556220 138226 556276 138236
rect 556108 131954 556164 131964
rect 555100 113138 555156 113148
rect 556332 110068 556388 159628
rect 556780 157556 556836 157566
rect 556444 154644 556500 154654
rect 556444 114772 556500 154588
rect 556556 149828 556612 149838
rect 556556 121044 556612 149772
rect 556668 149268 556724 149278
rect 556668 124180 556724 149212
rect 556780 133588 556836 157500
rect 556780 133522 556836 133532
rect 556668 124114 556724 124124
rect 556556 120978 556612 120988
rect 556444 114706 556500 114716
rect 556332 110002 556388 110012
rect 554988 108770 555044 108780
rect 554316 104132 554372 104142
rect 458556 99988 458612 99998
rect 457660 98756 457716 98766
rect 449372 98420 449428 98430
rect 449372 97860 449428 98364
rect 449372 97794 449428 97804
rect 457660 92708 457716 98700
rect 457660 92642 457716 92652
rect 458444 97860 458500 97870
rect 458444 72212 458500 97804
rect 458444 72146 458500 72156
rect 423164 68786 423220 68796
rect 422940 62514 422996 62524
rect 422716 57586 422772 57596
rect 458556 54852 458612 99932
rect 554316 99988 554372 104076
rect 554316 99922 554372 99932
rect 556892 70868 556948 161420
rect 557004 75572 557060 164668
rect 557788 149492 557844 149502
rect 557788 127316 557844 149436
rect 557900 142996 557956 165452
rect 560280 165004 560756 165060
rect 567224 165004 567812 165060
rect 574168 165004 574532 165060
rect 581112 165004 581252 165060
rect 560700 162596 560756 165004
rect 567756 162820 567812 165004
rect 567756 162754 567812 162764
rect 574476 162708 574532 165004
rect 581196 164724 581252 165004
rect 581196 164658 581252 164668
rect 574476 162642 574532 162652
rect 560700 162530 560756 162540
rect 558348 159796 558404 159806
rect 558236 152404 558292 152414
rect 557900 142930 557956 142940
rect 558012 151172 558068 151182
rect 557788 127250 557844 127260
rect 558012 88116 558068 151116
rect 558012 88050 558068 88060
rect 558124 147924 558180 147934
rect 558124 86548 558180 147868
rect 558236 128884 558292 152348
rect 558236 128818 558292 128828
rect 558124 86482 558180 86492
rect 558348 78708 558404 159740
rect 583660 157892 583716 394828
rect 583772 377188 583828 403228
rect 583772 377122 583828 377132
rect 583660 157826 583716 157836
rect 559468 157444 559524 157454
rect 558460 152852 558516 152862
rect 558460 83412 558516 152796
rect 559468 135156 559524 157388
rect 559580 157108 559636 157118
rect 559580 136724 559636 157052
rect 583884 156996 583940 404012
rect 590604 394884 590660 394894
rect 584668 393204 584724 393214
rect 584668 162820 584724 393148
rect 590492 392868 590548 392878
rect 590492 324548 590548 392812
rect 590604 364196 590660 394828
rect 590604 364130 590660 364140
rect 590492 324482 590548 324492
rect 590492 284676 590548 284686
rect 590492 165396 590548 284620
rect 590492 165330 590548 165340
rect 590604 245028 590660 245038
rect 590604 164164 590660 244972
rect 590604 164098 590660 164108
rect 590828 205380 590884 205390
rect 590828 163940 590884 205324
rect 590828 163874 590884 163884
rect 584668 162754 584724 162764
rect 583884 156930 583940 156940
rect 559580 136658 559636 136668
rect 559468 135090 559524 135100
rect 558460 83346 558516 83356
rect 558348 78642 558404 78652
rect 557004 75506 557060 75516
rect 556892 70802 556948 70812
rect 590492 73220 590548 73230
rect 557788 69300 557844 69310
rect 458556 54786 458612 54796
rect 554428 56084 554484 56094
rect 422492 52658 422548 52668
rect 421932 49634 421988 49644
rect 421708 49522 421764 49532
rect 420140 47954 420196 47964
rect 355180 45154 355236 45164
rect 554428 45220 554484 56028
rect 557788 50372 557844 69244
rect 558348 66164 558404 66174
rect 558124 63028 558180 63038
rect 557788 50306 557844 50316
rect 557900 59892 557956 59902
rect 557900 50260 557956 59836
rect 557900 50194 557956 50204
rect 558012 58324 558068 58334
rect 558012 48356 558068 58268
rect 558124 48468 558180 62972
rect 558236 61460 558292 61470
rect 558236 50148 558292 61404
rect 558236 50082 558292 50092
rect 558124 48402 558180 48412
rect 558012 48290 558068 48300
rect 558348 48244 558404 66108
rect 558348 48178 558404 48188
rect 590492 45332 590548 73164
rect 590604 60004 590660 60014
rect 590604 48692 590660 59948
rect 590604 48626 590660 48636
rect 590492 45266 590548 45276
rect 554428 45154 554484 45164
rect 343756 41346 343812 41356
rect 343532 41122 343588 41132
rect 336812 4274 336868 4284
rect 580860 5012 580916 5022
rect 284956 4162 285012 4172
rect 278012 4050 278068 4060
rect 580860 480 580916 4956
rect 207452 392 207704 480
rect 209356 392 209608 480
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 392 211540 480
rect 211288 -960 211512 392
rect 213192 -960 213416 480
rect 215096 -960 215320 480
rect 217000 -960 217224 480
rect 218904 -960 219128 480
rect 220808 -960 221032 480
rect 222712 -960 222936 480
rect 224616 -960 224840 480
rect 226520 -960 226744 480
rect 228424 -960 228648 480
rect 230328 -960 230552 480
rect 232232 -960 232456 480
rect 234136 -960 234360 480
rect 236040 -960 236264 480
rect 237944 -960 238168 480
rect 239848 -960 240072 480
rect 241752 -960 241976 480
rect 243656 -960 243880 480
rect 245560 -960 245784 480
rect 247464 -960 247688 480
rect 249368 -960 249592 480
rect 251272 -960 251496 480
rect 253176 -960 253400 480
rect 255080 -960 255304 480
rect 256984 -960 257208 480
rect 258888 -960 259112 480
rect 260792 -960 261016 480
rect 262696 -960 262920 480
rect 264600 -960 264824 480
rect 266504 -960 266728 480
rect 268408 -960 268632 480
rect 270312 -960 270536 480
rect 272216 -960 272440 480
rect 274120 -960 274344 480
rect 276024 -960 276248 480
rect 277928 -960 278152 480
rect 279832 -960 280056 480
rect 281736 -960 281960 480
rect 283640 -960 283864 480
rect 285544 -960 285768 480
rect 287448 -960 287672 480
rect 289352 -960 289576 480
rect 291256 -960 291480 480
rect 293160 -960 293384 480
rect 295064 -960 295288 480
rect 296968 -960 297192 480
rect 298872 -960 299096 480
rect 300776 -960 301000 480
rect 302680 -960 302904 480
rect 304584 -960 304808 480
rect 306488 -960 306712 480
rect 308392 -960 308616 480
rect 310296 -960 310520 480
rect 312200 -960 312424 480
rect 314104 -960 314328 480
rect 316008 -960 316232 480
rect 317912 -960 318136 480
rect 319816 -960 320040 480
rect 321720 -960 321944 480
rect 323624 -960 323848 480
rect 325528 -960 325752 480
rect 327432 -960 327656 480
rect 329336 -960 329560 480
rect 331240 -960 331464 480
rect 333144 -960 333368 480
rect 335048 -960 335272 480
rect 336952 -960 337176 480
rect 338856 -960 339080 480
rect 340760 -960 340984 480
rect 342664 -960 342888 480
rect 344568 -960 344792 480
rect 346472 -960 346696 480
rect 348376 -960 348600 480
rect 350280 -960 350504 480
rect 352184 -960 352408 480
rect 354088 -960 354312 480
rect 355992 -960 356216 480
rect 357896 -960 358120 480
rect 359800 -960 360024 480
rect 361704 -960 361928 480
rect 363608 -960 363832 480
rect 365512 -960 365736 480
rect 367416 -960 367640 480
rect 369320 -960 369544 480
rect 371224 -960 371448 480
rect 373128 -960 373352 480
rect 375032 -960 375256 480
rect 376936 -960 377160 480
rect 378840 -960 379064 480
rect 380744 -960 380968 480
rect 382648 -960 382872 480
rect 384552 -960 384776 480
rect 386456 -960 386680 480
rect 388360 -960 388584 480
rect 390264 -960 390488 480
rect 392168 -960 392392 480
rect 394072 -960 394296 480
rect 395976 -960 396200 480
rect 397880 -960 398104 480
rect 399784 -960 400008 480
rect 401688 -960 401912 480
rect 403592 -960 403816 480
rect 405496 -960 405720 480
rect 407400 -960 407624 480
rect 409304 -960 409528 480
rect 411208 -960 411432 480
rect 413112 -960 413336 480
rect 415016 -960 415240 480
rect 416920 -960 417144 480
rect 418824 -960 419048 480
rect 420728 -960 420952 480
rect 422632 -960 422856 480
rect 424536 -960 424760 480
rect 426440 -960 426664 480
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432152 -960 432376 480
rect 434056 -960 434280 480
rect 435960 -960 436184 480
rect 437864 -960 438088 480
rect 439768 -960 439992 480
rect 441672 -960 441896 480
rect 443576 -960 443800 480
rect 445480 -960 445704 480
rect 447384 -960 447608 480
rect 449288 -960 449512 480
rect 451192 -960 451416 480
rect 453096 -960 453320 480
rect 455000 -960 455224 480
rect 456904 -960 457128 480
rect 458808 -960 459032 480
rect 460712 -960 460936 480
rect 462616 -960 462840 480
rect 464520 -960 464744 480
rect 466424 -960 466648 480
rect 468328 -960 468552 480
rect 470232 -960 470456 480
rect 472136 -960 472360 480
rect 474040 -960 474264 480
rect 475944 -960 476168 480
rect 477848 -960 478072 480
rect 479752 -960 479976 480
rect 481656 -960 481880 480
rect 483560 -960 483784 480
rect 485464 -960 485688 480
rect 487368 -960 487592 480
rect 489272 -960 489496 480
rect 491176 -960 491400 480
rect 493080 -960 493304 480
rect 494984 -960 495208 480
rect 496888 -960 497112 480
rect 498792 -960 499016 480
rect 500696 -960 500920 480
rect 502600 -960 502824 480
rect 504504 -960 504728 480
rect 506408 -960 506632 480
rect 508312 -960 508536 480
rect 510216 -960 510440 480
rect 512120 -960 512344 480
rect 514024 -960 514248 480
rect 515928 -960 516152 480
rect 517832 -960 518056 480
rect 519736 -960 519960 480
rect 521640 -960 521864 480
rect 523544 -960 523768 480
rect 525448 -960 525672 480
rect 527352 -960 527576 480
rect 529256 -960 529480 480
rect 531160 -960 531384 480
rect 533064 -960 533288 480
rect 534968 -960 535192 480
rect 536872 -960 537096 480
rect 538776 -960 539000 480
rect 540680 -960 540904 480
rect 542584 -960 542808 480
rect 544488 -960 544712 480
rect 546392 -960 546616 480
rect 548296 -960 548520 480
rect 550200 -960 550424 480
rect 552104 -960 552328 480
rect 554008 -960 554232 480
rect 555912 -960 556136 480
rect 557816 -960 558040 480
rect 559720 -960 559944 480
rect 561624 -960 561848 480
rect 563528 -960 563752 480
rect 565432 -960 565656 480
rect 567336 -960 567560 480
rect 569240 -960 569464 480
rect 571144 -960 571368 480
rect 573048 -960 573272 480
rect 574952 -960 575176 480
rect 576856 -960 577080 480
rect 578760 -960 578984 480
rect 580664 392 580916 480
rect 582540 4340 582596 4350
rect 582540 480 582596 4284
rect 584444 4228 584500 4238
rect 584444 480 584500 4172
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 4172 502460 4228 502516
rect 4172 469532 4228 469588
rect 4508 388892 4564 388948
rect 4508 333340 4564 333396
rect 55356 590604 55412 590660
rect 33292 590492 33348 590548
rect 121548 590828 121604 590884
rect 99484 590716 99540 590772
rect 77308 583772 77364 583828
rect 153692 590716 153748 590772
rect 143388 582092 143444 582148
rect 152012 590604 152068 590660
rect 57932 573020 57988 573076
rect 56252 530684 56308 530740
rect 14252 488348 14308 488404
rect 93212 460124 93268 460180
rect 66332 417564 66388 417620
rect 64092 417004 64148 417060
rect 88172 417564 88228 417620
rect 68572 417452 68628 417508
rect 73052 417340 73108 417396
rect 70812 417228 70868 417284
rect 85036 417340 85092 417396
rect 75292 417116 75348 417172
rect 79772 416892 79828 416948
rect 77532 416668 77588 416724
rect 82012 416780 82068 416836
rect 84812 416668 84868 416724
rect 61852 413308 61908 413364
rect 57932 390908 57988 390964
rect 59612 403676 59668 403732
rect 59612 390796 59668 390852
rect 56252 390684 56308 390740
rect 14252 390572 14308 390628
rect 78428 388108 78484 388164
rect 40908 386428 40964 386484
rect 38444 383292 38500 383348
rect 24332 383068 24388 383124
rect 11004 301532 11060 301588
rect 14252 380156 14308 380212
rect 13244 224252 13300 224308
rect 4172 121436 4228 121492
rect 4172 50316 4228 50372
rect 11564 5852 11620 5908
rect 22764 232876 22820 232932
rect 14252 191996 14308 192052
rect 18956 229292 19012 229348
rect 15372 4172 15428 4228
rect 17276 4172 17332 4228
rect 21084 4172 21140 4228
rect 38332 380380 38388 380436
rect 34412 379596 34468 379652
rect 34412 276668 34468 276724
rect 38220 379484 38276 379540
rect 38220 238252 38276 238308
rect 38444 240716 38500 240772
rect 38556 383180 38612 383236
rect 38556 238476 38612 238532
rect 40236 292348 40292 292404
rect 38332 238140 38388 238196
rect 35196 236124 35252 236180
rect 34188 232652 34244 232708
rect 24332 149660 24388 149716
rect 24668 214172 24724 214228
rect 30380 212604 30436 212660
rect 27692 79100 27748 79156
rect 27692 50204 27748 50260
rect 26796 4172 26852 4228
rect 32508 4172 32564 4228
rect 38556 232764 38612 232820
rect 37996 227724 38052 227780
rect 35196 4620 35252 4676
rect 36876 222684 36932 222740
rect 36876 4396 36932 4452
rect 38444 217532 38500 217588
rect 39900 221004 39956 221060
rect 39788 212492 39844 212548
rect 39788 4508 39844 4564
rect 38556 4284 38612 4340
rect 38444 4060 38500 4116
rect 40124 214284 40180 214340
rect 40012 212716 40068 212772
rect 69692 386092 69748 386148
rect 55580 380940 55636 380996
rect 49532 379036 49588 379092
rect 63196 363692 63252 363748
rect 59388 363020 59444 363076
rect 67004 362908 67060 362964
rect 74620 379372 74676 379428
rect 69692 362908 69748 362964
rect 70812 363804 70868 363860
rect 86492 417116 86548 417172
rect 85260 417004 85316 417060
rect 85260 397516 85316 397572
rect 86716 416892 86772 416948
rect 87276 409052 87332 409108
rect 87276 407372 87332 407428
rect 88172 397516 88228 397572
rect 91532 417452 91588 417508
rect 86716 397292 86772 397348
rect 93212 409612 93268 409668
rect 152012 409500 152068 409556
rect 153692 395612 153748 395668
rect 155372 590492 155428 590548
rect 160412 446012 160468 446068
rect 160412 398972 160468 399028
rect 168812 590828 168868 590884
rect 186396 590492 186452 590548
rect 173852 583772 173908 583828
rect 168812 409388 168868 409444
rect 170492 582092 170548 582148
rect 168028 407372 168084 407428
rect 168028 406588 168084 406644
rect 165452 397852 165508 397908
rect 168028 405692 168084 405748
rect 168028 404908 168084 404964
rect 155372 392588 155428 392644
rect 91532 392364 91588 392420
rect 86492 392252 86548 392308
rect 85036 383964 85092 384020
rect 85708 391580 85764 391636
rect 84812 383852 84868 383908
rect 82236 379820 82292 379876
rect 103292 386876 103348 386932
rect 96572 386764 96628 386820
rect 94892 386652 94948 386708
rect 93660 380044 93716 380100
rect 91532 379932 91588 379988
rect 85708 363020 85764 363076
rect 85708 361228 85764 361284
rect 86044 363916 86100 363972
rect 89852 362908 89908 362964
rect 91532 362908 91588 362964
rect 49532 319004 49588 319060
rect 46284 293132 46340 293188
rect 51660 293132 51716 293188
rect 59052 293916 59108 293972
rect 46284 292348 46340 292404
rect 87276 293132 87332 293188
rect 71820 292348 71876 292404
rect 84588 292348 84644 292404
rect 87276 290332 87332 290388
rect 93212 250572 93268 250628
rect 40684 238364 40740 238420
rect 40908 248444 40964 248500
rect 90188 241164 90244 241220
rect 41132 240716 41188 240772
rect 66220 240716 66276 240772
rect 71596 240716 71652 240772
rect 80556 240604 80612 240660
rect 90188 240604 90244 240660
rect 60844 240492 60900 240548
rect 57260 240380 57316 240436
rect 53676 240268 53732 240324
rect 46508 240156 46564 240212
rect 85932 240156 85988 240212
rect 42924 238476 42980 238532
rect 44716 238252 44772 238308
rect 48300 238140 48356 238196
rect 55468 240044 55524 240100
rect 51884 238364 51940 238420
rect 50092 237916 50148 237972
rect 41020 235116 41076 235172
rect 41020 234444 41076 234500
rect 40908 227836 40964 227892
rect 40684 224476 40740 224532
rect 40684 48188 40740 48244
rect 40796 224364 40852 224420
rect 40908 50092 40964 50148
rect 41132 234332 41188 234388
rect 62636 238476 62692 238532
rect 64428 238476 64484 238532
rect 69804 238140 69860 238196
rect 73388 237916 73444 237972
rect 76972 238028 77028 238084
rect 75180 237804 75236 237860
rect 82348 239820 82404 239876
rect 87724 238476 87780 238532
rect 84140 238364 84196 238420
rect 89516 238252 89572 238308
rect 78764 237692 78820 237748
rect 68012 237580 68068 237636
rect 59052 233436 59108 233492
rect 93212 229404 93268 229460
rect 93324 246316 93380 246372
rect 93436 241948 93492 242004
rect 95116 386540 95172 386596
rect 95340 385420 95396 385476
rect 95340 238476 95396 238532
rect 95564 383404 95620 383460
rect 95116 238252 95172 238308
rect 95564 238140 95620 238196
rect 94892 238028 94948 238084
rect 96572 237692 96628 237748
rect 96796 385084 96852 385140
rect 99932 384972 99988 385028
rect 99932 238364 99988 238420
rect 103292 237916 103348 237972
rect 104972 385308 105028 385364
rect 111692 382620 111748 382676
rect 108332 321692 108388 321748
rect 106652 320012 106708 320068
rect 108332 267596 108388 267652
rect 106652 263340 106708 263396
rect 167132 382060 167188 382116
rect 118412 381836 118468 381892
rect 111692 241052 111748 241108
rect 113372 381724 113428 381780
rect 116732 381500 116788 381556
rect 116732 241164 116788 241220
rect 118412 240716 118468 240772
rect 120092 381612 120148 381668
rect 113372 239932 113428 239988
rect 121772 380268 121828 380324
rect 120204 378924 120260 378980
rect 121772 363916 121828 363972
rect 120204 361340 120260 361396
rect 152796 321804 152852 321860
rect 144284 290332 144340 290388
rect 144284 289772 144340 289828
rect 161308 294812 161364 294868
rect 167244 356300 167300 356356
rect 168028 342860 168084 342916
rect 168140 346220 168196 346276
rect 167244 321804 167300 321860
rect 168140 320012 168196 320068
rect 168812 381948 168868 382004
rect 167132 240044 167188 240100
rect 167244 318220 167300 318276
rect 120092 239820 120148 239876
rect 104972 237804 105028 237860
rect 96796 237580 96852 237636
rect 93436 230972 93492 231028
rect 93324 227612 93380 227668
rect 154924 217644 154980 217700
rect 169148 289884 169204 289940
rect 169036 286412 169092 286468
rect 168924 284732 168980 284788
rect 169148 283948 169204 284004
rect 169260 288092 169316 288148
rect 169260 279916 169316 279972
rect 169372 286524 169428 286580
rect 169372 277900 169428 277956
rect 169036 275884 169092 275940
rect 172172 397740 172228 397796
rect 170492 274540 170548 274596
rect 170604 382172 170660 382228
rect 168924 273868 168980 273924
rect 172172 322700 172228 322756
rect 172956 331660 173012 331716
rect 170604 240268 170660 240324
rect 168812 240156 168868 240212
rect 183036 578732 183092 578788
rect 180572 417228 180628 417284
rect 177212 416780 177268 416836
rect 177212 397628 177268 397684
rect 175532 395724 175588 395780
rect 173964 392812 174020 392868
rect 177324 392700 177380 392756
rect 177212 357420 177268 357476
rect 176204 355180 176260 355236
rect 175532 332780 175588 332836
rect 176092 347340 176148 347396
rect 173964 330876 174020 330932
rect 173852 275660 173908 275716
rect 174412 330540 174468 330596
rect 175980 328300 176036 328356
rect 174636 326060 174692 326116
rect 174412 229964 174468 230020
rect 174524 324940 174580 324996
rect 172956 224812 173012 224868
rect 174524 222908 174580 222964
rect 175532 301532 175588 301588
rect 175532 276780 175588 276836
rect 175644 283052 175700 283108
rect 175644 272076 175700 272132
rect 175980 233212 176036 233268
rect 176092 231196 176148 231252
rect 176204 231084 176260 231140
rect 176316 349468 176372 349524
rect 180572 384076 180628 384132
rect 181356 352940 181412 352996
rect 177884 351820 177940 351876
rect 177324 336812 177380 336868
rect 177772 345100 177828 345156
rect 177212 294812 177268 294868
rect 179452 348460 179508 348516
rect 177884 232988 177940 233044
rect 177996 346220 178052 346276
rect 177772 228060 177828 228116
rect 176316 224588 176372 224644
rect 174636 221228 174692 221284
rect 179340 340620 179396 340676
rect 179228 327180 179284 327236
rect 179228 234780 179284 234836
rect 179676 343980 179732 344036
rect 179452 234668 179508 234724
rect 179564 339500 179620 339556
rect 179340 231308 179396 231364
rect 179564 224700 179620 224756
rect 181132 342860 181188 342916
rect 181020 335020 181076 335076
rect 181132 229740 181188 229796
rect 181244 338380 181300 338436
rect 181020 228172 181076 228228
rect 182700 341740 182756 341796
rect 181356 229628 181412 229684
rect 182588 323820 182644 323876
rect 181244 222796 181300 222852
rect 179676 222572 179732 222628
rect 177996 221116 178052 221172
rect 182924 336140 182980 336196
rect 182700 233100 182756 233156
rect 182812 329420 182868 329476
rect 182588 219548 182644 219604
rect 167244 217644 167300 217700
rect 184716 575484 184772 575540
rect 184604 354060 184660 354116
rect 183036 273420 183092 273476
rect 184492 337260 184548 337316
rect 182924 219324 182980 219380
rect 186284 566076 186340 566132
rect 186172 543564 186228 543620
rect 186060 529228 186116 529284
rect 185612 411964 185668 412020
rect 186060 389004 186116 389060
rect 186284 407932 186340 407988
rect 189756 588812 189812 588868
rect 189644 577052 189700 577108
rect 187516 566076 187572 566132
rect 189308 575372 189364 575428
rect 187964 557900 188020 557956
rect 186396 404012 186452 404068
rect 187292 507724 187348 507780
rect 186172 387212 186228 387268
rect 185612 385532 185668 385588
rect 185724 383516 185780 383572
rect 184716 267820 184772 267876
rect 185612 382284 185668 382340
rect 185724 363804 185780 363860
rect 185948 380492 186004 380548
rect 185948 363692 186004 363748
rect 186396 332780 186452 332836
rect 185612 240380 185668 240436
rect 186284 322700 186340 322756
rect 186284 234892 186340 234948
rect 184604 227948 184660 228004
rect 186508 296492 186564 296548
rect 187292 289884 187348 289940
rect 187404 493388 187460 493444
rect 187404 288092 187460 288148
rect 187516 486220 187572 486276
rect 186508 284732 186564 284788
rect 187068 287308 187124 287364
rect 187740 479052 187796 479108
rect 187516 286524 187572 286580
rect 187628 464716 187684 464772
rect 187740 286412 187796 286468
rect 187852 457548 187908 457604
rect 187628 283052 187684 283108
rect 187068 282044 187124 282100
rect 187964 409276 188020 409332
rect 188076 414540 188132 414596
rect 189532 572012 189588 572068
rect 189308 407372 189364 407428
rect 189420 570332 189476 570388
rect 189308 350700 189364 350756
rect 189196 333900 189252 333956
rect 188076 289772 188132 289828
rect 189084 321580 189140 321636
rect 188076 288988 188132 289044
rect 188972 288988 189028 289044
rect 188076 280588 188132 280644
rect 188076 252140 188132 252196
rect 187964 251020 188020 251076
rect 187964 217980 188020 218036
rect 186396 217756 186452 217812
rect 184492 217644 184548 217700
rect 182812 215964 182868 216020
rect 188972 240156 189028 240212
rect 189420 272300 189476 272356
rect 189644 271180 189700 271236
rect 231644 591276 231700 591332
rect 209580 578732 209636 578788
rect 297836 591164 297892 591220
rect 319900 591052 319956 591108
rect 364028 590940 364084 590996
rect 386092 590828 386148 590884
rect 430220 590716 430276 590772
rect 452284 590156 452340 590212
rect 408268 588812 408324 588868
rect 341964 577052 342020 577108
rect 496412 590604 496468 590660
rect 518700 590604 518756 590660
rect 529788 590604 529844 590660
rect 474348 572012 474404 572068
rect 275772 570332 275828 570388
rect 253708 568652 253764 568708
rect 529340 526764 529396 526820
rect 197596 395724 197652 395780
rect 192444 392812 192500 392868
rect 207900 408492 207956 408548
rect 207900 406700 207956 406756
rect 210364 407372 210420 407428
rect 202748 392700 202804 392756
rect 207004 403228 207060 403284
rect 205100 389116 205156 389172
rect 202748 382508 202804 382564
rect 201404 382396 201460 382452
rect 204204 382508 204260 382564
rect 203084 382396 203140 382452
rect 204876 382396 204932 382452
rect 208348 402332 208404 402388
rect 206108 382508 206164 382564
rect 206444 382396 206500 382452
rect 208124 382396 208180 382452
rect 213052 406028 213108 406084
rect 218204 406588 218260 406644
rect 218204 405804 218260 405860
rect 211036 404012 211092 404068
rect 211708 399084 211764 399140
rect 219100 398972 219156 399028
rect 215068 397852 215124 397908
rect 211596 394492 211652 394548
rect 211596 391020 211652 391076
rect 209468 382508 209524 382564
rect 209804 382396 209860 382452
rect 213612 395836 213668 395892
rect 212268 392812 212324 392868
rect 212940 392700 212996 392756
rect 214284 395724 214340 395780
rect 215628 395612 215684 395668
rect 216300 392588 216356 392644
rect 216972 390908 217028 390964
rect 217644 390684 217700 390740
rect 218540 390572 218596 390628
rect 228508 409836 228564 409892
rect 243964 407596 244020 407652
rect 238812 407484 238868 407540
rect 233660 407372 233716 407428
rect 254268 407148 254324 407204
rect 259420 408044 259476 408100
rect 249116 407036 249172 407092
rect 228508 406588 228564 406644
rect 263788 407708 263844 407764
rect 259420 406588 259476 406644
rect 260428 406588 260484 406644
rect 252700 406364 252756 406420
rect 252028 405804 252084 405860
rect 251356 405692 251412 405748
rect 250012 400652 250068 400708
rect 223356 398076 223412 398132
rect 248668 398972 248724 399028
rect 219660 390796 219716 390852
rect 240828 386876 240884 386932
rect 232764 386428 232820 386484
rect 228732 383292 228788 383348
rect 223468 383068 223524 383124
rect 222572 380156 222628 380212
rect 226492 382060 226548 382116
rect 226492 381388 226548 381444
rect 226716 382060 226772 382116
rect 229292 383180 229348 383236
rect 230636 381388 230692 381444
rect 231868 380380 231924 380436
rect 237468 385196 237524 385252
rect 235228 382284 235284 382340
rect 233548 382172 233604 382228
rect 233996 381724 234052 381780
rect 236124 381388 236180 381444
rect 236908 380604 236964 380660
rect 238812 385084 238868 385140
rect 238588 381836 238644 381892
rect 239372 383404 239428 383460
rect 240268 382620 240324 382676
rect 242844 386764 242900 386820
rect 242172 386652 242228 386708
rect 242060 385308 242116 385364
rect 247100 386540 247156 386596
rect 246204 385420 246260 385476
rect 245420 384972 245476 385028
rect 244076 381612 244132 381668
rect 243740 381500 243796 381556
rect 245532 381948 245588 382004
rect 248556 385756 248612 385812
rect 250572 390572 250628 390628
rect 249788 381948 249844 382004
rect 252028 404012 252084 404068
rect 252476 385868 252532 385924
rect 259420 405916 259476 405972
rect 257852 404796 257908 404852
rect 253260 390684 253316 390740
rect 256620 385644 256676 385700
rect 255052 382956 255108 383012
rect 254716 382284 254772 382340
rect 256060 382172 256116 382228
rect 257852 382956 257908 383012
rect 257964 387324 258020 387380
rect 256956 382732 257012 382788
rect 260316 387436 260372 387492
rect 258636 382396 258692 382452
rect 259196 381948 259252 382004
rect 261212 405804 261268 405860
rect 262780 404684 262836 404740
rect 262108 399084 262164 399140
rect 261212 382284 261268 382340
rect 261324 382620 261380 382676
rect 260428 380828 260484 380884
rect 261996 382284 262052 382340
rect 263452 399196 263508 399252
rect 268156 408604 268212 408660
rect 266812 404572 266868 404628
rect 264124 402892 264180 402948
rect 265468 399756 265524 399812
rect 264796 399308 264852 399364
rect 263788 380716 263844 380772
rect 267484 402444 267540 402500
rect 268940 407820 268996 407876
rect 268828 400764 268884 400820
rect 280476 409388 280532 409444
rect 274652 407932 274708 407988
rect 268940 385980 268996 386036
rect 270172 401324 270228 401380
rect 274204 401212 274260 401268
rect 271516 400988 271572 401044
rect 266588 381948 266644 382004
rect 270732 396284 270788 396340
rect 269948 384188 270004 384244
rect 272860 400876 272916 400932
rect 272300 396172 272356 396228
rect 273420 395948 273476 396004
rect 280252 408380 280308 408436
rect 279580 402668 279636 402724
rect 278236 402556 278292 402612
rect 275548 401100 275604 401156
rect 274652 384972 274708 385028
rect 274652 380604 274708 380660
rect 274764 395836 274820 395892
rect 276108 395724 276164 395780
rect 277452 395612 277508 395668
rect 276780 394492 276836 394548
rect 283948 409500 284004 409556
rect 280476 406588 280532 406644
rect 282268 409052 282324 409108
rect 280924 402780 280980 402836
rect 283612 406252 283668 406308
rect 279356 382060 279412 382116
rect 281708 381948 281764 382004
rect 283388 385980 283444 386036
rect 285180 409500 285236 409556
rect 289772 409164 289828 409220
rect 286300 406140 286356 406196
rect 284732 404236 284788 404292
rect 284284 399420 284340 399476
rect 283948 384412 284004 384468
rect 288316 399644 288372 399700
rect 286860 390796 286916 390852
rect 284732 382060 284788 382116
rect 285516 382844 285572 382900
rect 286076 382508 286132 382564
rect 288092 381948 288148 382004
rect 295596 408940 295652 408996
rect 295596 406588 295652 406644
rect 298172 409164 298228 409220
rect 297052 396956 297108 397012
rect 294924 392812 294980 392868
rect 293580 392588 293636 392644
rect 291564 387660 291620 387716
rect 289772 384524 289828 384580
rect 290220 387548 290276 387604
rect 289548 382732 289604 382788
rect 290556 381948 290612 382004
rect 292236 382060 292292 382116
rect 293468 381948 293524 382004
rect 292908 380156 292964 380212
rect 294252 390908 294308 390964
rect 295820 391132 295876 391188
rect 296828 387772 296884 387828
rect 298060 387884 298116 387940
rect 305788 409612 305844 409668
rect 300636 408044 300692 408100
rect 300412 401660 300468 401716
rect 299740 399868 299796 399924
rect 299068 396844 299124 396900
rect 298172 382620 298228 382676
rect 298284 394716 298340 394772
rect 303772 398188 303828 398244
rect 302540 396060 302596 396116
rect 301644 394604 301700 394660
rect 301532 382732 301588 382788
rect 305004 394940 305060 394996
rect 304332 394044 304388 394100
rect 303548 382620 303604 382676
rect 305900 394828 305956 394884
rect 310940 409724 310996 409780
rect 307132 408268 307188 408324
rect 308252 404124 308308 404180
rect 307692 394268 307748 394324
rect 306572 380604 306628 380660
rect 306908 382060 306964 382116
rect 310492 397740 310548 397796
rect 309820 396620 309876 396676
rect 308252 382844 308308 382900
rect 308364 393820 308420 393876
rect 309260 391244 309316 391300
rect 311052 391356 311108 391412
rect 313740 390460 313796 390516
rect 313068 382844 313124 382900
rect 311612 380716 311668 380772
rect 312396 381948 312452 382004
rect 313628 381948 313684 382004
rect 320908 389788 320964 389844
rect 324604 397516 324660 397572
rect 323932 397404 323988 397460
rect 321244 389788 321300 389844
rect 321804 391020 321860 391076
rect 320908 388892 320964 388948
rect 318444 388108 318500 388164
rect 315868 384748 315924 384804
rect 315868 384300 315924 384356
rect 316092 386092 316148 386148
rect 315084 381948 315140 382004
rect 315196 380940 315252 380996
rect 315868 380492 315924 380548
rect 316652 383516 316708 383572
rect 320012 382956 320068 383012
rect 320012 382060 320068 382116
rect 319340 380268 319396 380324
rect 320908 380044 320964 380100
rect 320572 379932 320628 379988
rect 322700 385532 322756 385588
rect 329308 397628 329364 397684
rect 328636 397292 328692 397348
rect 325164 392364 325220 392420
rect 322924 381948 322980 382004
rect 325836 384860 325892 384916
rect 327180 392252 327236 392308
rect 325948 384076 326004 384132
rect 325836 380492 325892 380548
rect 326284 383964 326340 384020
rect 327628 383852 327684 383908
rect 336700 383852 336756 383908
rect 341180 409276 341236 409332
rect 331548 381276 331604 381332
rect 339388 383068 339444 383124
rect 319228 379820 319284 379876
rect 200844 379708 200900 379764
rect 202188 379708 202244 379764
rect 220444 379596 220500 379652
rect 222012 379484 222068 379540
rect 224028 379484 224084 379540
rect 227612 379484 227668 379540
rect 229068 379484 229124 379540
rect 230524 379484 230580 379540
rect 235452 379484 235508 379540
rect 317884 379372 317940 379428
rect 221116 379260 221172 379316
rect 221788 379260 221844 379316
rect 225148 379260 225204 379316
rect 225820 379260 225876 379316
rect 227836 379260 227892 379316
rect 232540 379260 232596 379316
rect 340172 380156 340228 380212
rect 339388 344204 339444 344260
rect 339612 356300 339668 356356
rect 189756 270060 189812 270116
rect 339500 271180 339556 271236
rect 189532 268940 189588 268996
rect 339388 267708 339444 267764
rect 194908 240156 194964 240212
rect 189308 229852 189364 229908
rect 196700 232876 196756 232932
rect 195804 224252 195860 224308
rect 189196 219436 189252 219492
rect 189084 217868 189140 217924
rect 188076 214732 188132 214788
rect 199388 227836 199444 227892
rect 198492 227724 198548 227780
rect 200284 224476 200340 224532
rect 201180 217532 201236 217588
rect 203868 229516 203924 229572
rect 205660 234444 205716 234500
rect 208348 236908 208404 236964
rect 207452 234556 207508 234612
rect 206556 234332 206612 234388
rect 210140 231756 210196 231812
rect 209244 231532 209300 231588
rect 211932 231644 211988 231700
rect 211036 231420 211092 231476
rect 212828 230860 212884 230916
rect 216412 228396 216468 228452
rect 215516 228284 215572 228340
rect 214620 227836 214676 227892
rect 213724 227724 213780 227780
rect 217308 227500 217364 227556
rect 204764 224364 204820 224420
rect 219100 225036 219156 225092
rect 221788 224476 221844 224532
rect 220892 224364 220948 224420
rect 219996 224252 220052 224308
rect 218204 224140 218260 224196
rect 202972 222684 203028 222740
rect 223580 234444 223636 234500
rect 224476 221564 224532 221620
rect 222684 221452 222740 221508
rect 226268 236908 226324 236964
rect 228060 232764 228116 232820
rect 227164 221004 227220 221060
rect 228956 215852 229012 215908
rect 230748 214396 230804 214452
rect 229852 214284 229908 214340
rect 225372 214172 225428 214228
rect 202076 212716 202132 212772
rect 197596 212604 197652 212660
rect 233436 236908 233492 236964
rect 235228 237020 235284 237076
rect 236684 236908 236740 236964
rect 237020 236908 237076 236964
rect 234332 234220 234388 234276
rect 238812 236908 238868 236964
rect 240604 236908 240660 236964
rect 239708 232876 239764 232932
rect 237916 232764 237972 232820
rect 232540 225932 232596 225988
rect 242396 237020 242452 237076
rect 244188 238476 244244 238532
rect 245084 238476 245140 238532
rect 246876 238252 246932 238308
rect 250460 238364 250516 238420
rect 252252 238476 252308 238532
rect 251356 238140 251412 238196
rect 249564 238028 249620 238084
rect 248668 237916 248724 237972
rect 247772 237804 247828 237860
rect 245980 237692 246036 237748
rect 253148 237468 253204 237524
rect 243516 236908 243572 236964
rect 254044 214956 254100 215012
rect 255836 215852 255892 215908
rect 254940 214284 254996 214340
rect 241500 213276 241556 213332
rect 231644 212492 231700 212548
rect 259420 216524 259476 216580
rect 258524 214396 258580 214452
rect 257628 214060 257684 214116
rect 260316 212492 260372 212548
rect 256732 212380 256788 212436
rect 262108 216636 262164 216692
rect 263900 211484 263956 211540
rect 263004 210700 263060 210756
rect 267484 237020 267540 237076
rect 267036 236908 267092 236964
rect 268604 236908 268660 236964
rect 265692 211596 265748 211652
rect 264796 210028 264852 210084
rect 261212 209916 261268 209972
rect 269052 209580 269108 209636
rect 269052 209132 269108 209188
rect 269724 238476 269780 238532
rect 269612 237468 269668 237524
rect 269276 145292 269332 145348
rect 269388 227500 269444 227556
rect 41132 49644 41188 49700
rect 45612 50092 45668 50148
rect 41020 49532 41076 49588
rect 40796 47964 40852 48020
rect 40236 46956 40292 47012
rect 45388 46956 45444 47012
rect 45388 5852 45444 5908
rect 40124 4956 40180 5012
rect 40012 4844 40068 4900
rect 42028 4620 42084 4676
rect 41804 4172 41860 4228
rect 42028 4172 42084 4228
rect 49868 49756 49924 49812
rect 49644 49644 49700 49700
rect 46956 47852 47012 47908
rect 46956 47068 47012 47124
rect 47516 4284 47572 4340
rect 49644 4284 49700 4340
rect 49420 4172 49476 4228
rect 87500 49532 87556 49588
rect 49868 4172 49924 4228
rect 53228 48188 53284 48244
rect 77980 48076 78036 48132
rect 62748 46172 62804 46228
rect 60844 4956 60900 5012
rect 58940 4060 58996 4116
rect 55132 3388 55188 3444
rect 57148 3388 57204 3444
rect 68460 42812 68516 42868
rect 64652 4844 64708 4900
rect 66556 4732 66612 4788
rect 76076 4620 76132 4676
rect 72268 4508 72324 4564
rect 70364 4396 70420 4452
rect 74396 4060 74452 4116
rect 81788 47964 81844 48020
rect 79884 41132 79940 41188
rect 85708 41244 85764 41300
rect 83692 37772 83748 37828
rect 95116 49532 95172 49588
rect 91308 41356 91364 41412
rect 89628 4060 89684 4116
rect 93212 4284 93268 4340
rect 161756 50092 161812 50148
rect 156044 49980 156100 50036
rect 150332 49868 150388 49924
rect 144620 49756 144676 49812
rect 97356 48636 97412 48692
rect 97356 47852 97412 47908
rect 112252 49644 112308 49700
rect 106540 44604 106596 44660
rect 100828 44492 100884 44548
rect 97244 4844 97300 4900
rect 98924 4172 98980 4228
rect 102956 4172 103012 4228
rect 104860 4060 104916 4116
rect 108444 41468 108500 41524
rect 110796 4172 110852 4228
rect 138908 48188 138964 48244
rect 133196 48076 133252 48132
rect 127484 47964 127540 48020
rect 121772 47852 121828 47908
rect 119868 43036 119924 43092
rect 114268 42924 114324 42980
rect 117964 41580 118020 41636
rect 116284 4284 116340 4340
rect 125580 46284 125636 46340
rect 123676 41692 123732 41748
rect 131292 46396 131348 46452
rect 129388 41916 129444 41972
rect 135324 4396 135380 4452
rect 137228 3388 137284 3444
rect 142828 43148 142884 43204
rect 140812 38220 140868 38276
rect 146524 38108 146580 38164
rect 148652 3388 148708 3444
rect 152236 44716 152292 44772
rect 154476 4060 154532 4116
rect 158172 5852 158228 5908
rect 160076 4508 160132 4564
rect 201740 48524 201796 48580
rect 196028 48300 196084 48356
rect 190316 45276 190372 45332
rect 184604 45164 184660 45220
rect 178892 45052 178948 45108
rect 173180 44940 173236 44996
rect 167468 44828 167524 44884
rect 163884 7532 163940 7588
rect 165788 4732 165844 4788
rect 169372 29372 169428 29428
rect 171500 4620 171556 4676
rect 175084 43372 175140 43428
rect 176988 43260 177044 43316
rect 180796 41020 180852 41076
rect 182700 37884 182756 37940
rect 188412 37996 188468 38052
rect 186508 31052 186564 31108
rect 192332 41804 192388 41860
rect 192220 12572 192276 12628
rect 192332 4844 192388 4900
rect 194348 4844 194404 4900
rect 199948 46508 200004 46564
rect 197932 39452 197988 39508
rect 203644 48412 203700 48468
rect 269388 50092 269444 50148
rect 269500 224140 269556 224196
rect 212268 47740 212324 47796
rect 269500 44828 269556 44884
rect 207452 44380 207508 44436
rect 205772 4956 205828 5012
rect 209356 31164 209412 31220
rect 269836 210812 269892 210868
rect 269836 207900 269892 207956
rect 270172 146972 270228 147028
rect 270508 238364 270564 238420
rect 269724 48412 269780 48468
rect 269612 31164 269668 31220
rect 270844 228396 270900 228452
rect 270732 227724 270788 227780
rect 270620 225036 270676 225092
rect 270844 49980 270900 50036
rect 270956 228284 271012 228340
rect 271292 230972 271348 231028
rect 271068 133532 271124 133588
rect 271180 227836 271236 227892
rect 270956 49868 271012 49924
rect 271292 196364 271348 196420
rect 271180 49756 271236 49812
rect 271292 145404 271348 145460
rect 270732 48188 270788 48244
rect 270620 44940 270676 44996
rect 272860 238252 272916 238308
rect 273420 239820 273476 239876
rect 272300 235116 272356 235172
rect 272188 209468 272244 209524
rect 272188 180796 272244 180852
rect 272300 153580 272356 153636
rect 272412 211260 272468 211316
rect 272524 209804 272580 209860
rect 272748 209580 272804 209636
rect 272636 209468 272692 209524
rect 272860 209132 272916 209188
rect 272860 177884 272916 177940
rect 272972 203084 273028 203140
rect 272748 174972 272804 175028
rect 272636 166236 272692 166292
rect 272524 157500 272580 157556
rect 272412 148764 272468 148820
rect 272188 131292 272244 131348
rect 272300 143612 272356 143668
rect 271964 106652 272020 106708
rect 272412 140252 272468 140308
rect 273308 154364 273364 154420
rect 273084 154140 273140 154196
rect 273084 134204 273140 134260
rect 273196 144508 273252 144564
rect 273308 137116 273364 137172
rect 273196 128380 273252 128436
rect 273756 237580 273812 237636
rect 273980 238028 274036 238084
rect 273756 234444 273812 234500
rect 273756 202412 273812 202468
rect 273868 213276 273924 213332
rect 273420 105084 273476 105140
rect 272972 99260 273028 99316
rect 273084 91532 273140 91588
rect 272972 89852 273028 89908
rect 273084 78876 273140 78932
rect 272972 73052 273028 73108
rect 272412 50316 272468 50372
rect 272972 70140 273028 70196
rect 272300 50204 272356 50260
rect 273196 67228 273252 67284
rect 273084 64316 273140 64372
rect 273084 49980 273140 50036
rect 272972 48076 273028 48132
rect 273756 58492 273812 58548
rect 273756 49868 273812 49924
rect 273196 47964 273252 48020
rect 271292 36764 271348 36820
rect 270508 12572 270564 12628
rect 274092 237916 274148 237972
rect 274764 227612 274820 227668
rect 274764 200732 274820 200788
rect 274652 104972 274708 105028
rect 274764 128492 274820 128548
rect 276332 239708 276388 239764
rect 275548 125132 275604 125188
rect 275660 238140 275716 238196
rect 274764 81788 274820 81844
rect 274876 107100 274932 107156
rect 274876 75964 274932 76020
rect 274204 52668 274260 52724
rect 274204 49756 274260 49812
rect 274092 41020 274148 41076
rect 275884 224476 275940 224532
rect 275772 224252 275828 224308
rect 275884 45276 275940 45332
rect 275996 224364 276052 224420
rect 275996 45164 276052 45220
rect 276108 221564 276164 221620
rect 275772 45052 275828 45108
rect 276220 221452 276276 221508
rect 276332 199836 276388 199892
rect 277340 131852 277396 131908
rect 278012 238924 278068 238980
rect 276444 115052 276500 115108
rect 276220 48300 276276 48356
rect 276108 44380 276164 44436
rect 275660 39452 275716 39508
rect 273980 31052 274036 31108
rect 273868 4396 273924 4452
rect 211484 4060 211540 4116
rect 278236 135212 278292 135268
rect 278908 237692 278964 237748
rect 279132 152236 279188 152292
rect 279692 239596 279748 239652
rect 278908 7532 278964 7588
rect 279916 237580 279972 237636
rect 279804 214060 279860 214116
rect 280028 152684 280084 152740
rect 280588 237804 280644 237860
rect 279916 131964 279972 132020
rect 279804 103292 279860 103348
rect 280924 236908 280980 236964
rect 280700 234556 280756 234612
rect 280700 203084 280756 203140
rect 281372 214956 281428 215012
rect 282716 237468 282772 237524
rect 281820 160188 281876 160244
rect 283052 235004 283108 235060
rect 283052 233436 283108 233492
rect 281372 103740 281428 103796
rect 284508 160636 284564 160692
rect 284732 237692 284788 237748
rect 283612 160300 283668 160356
rect 283052 90524 283108 90580
rect 280588 43372 280644 43428
rect 284956 214172 285012 214228
rect 284844 212380 284900 212436
rect 284844 103628 284900 103684
rect 284732 4956 284788 5012
rect 279692 4732 279748 4788
rect 285404 152124 285460 152180
rect 287196 237580 287252 237636
rect 287980 239820 288036 239876
rect 286300 148988 286356 149044
rect 286412 219772 286468 219828
rect 286412 48188 286468 48244
rect 286524 214732 286580 214788
rect 286524 45276 286580 45332
rect 288428 236908 288484 236964
rect 288204 152572 288260 152628
rect 288316 216524 288372 216580
rect 288428 155820 288484 155876
rect 289100 239260 289156 239316
rect 289100 238476 289156 238532
rect 289772 217980 289828 218036
rect 288988 150892 289044 150948
rect 289660 216636 289716 216692
rect 288316 103516 288372 103572
rect 289660 103404 289716 103460
rect 288204 61404 288260 61460
rect 288204 49644 288260 49700
rect 288988 55580 289044 55636
rect 288988 49532 289044 49588
rect 289884 149100 289940 149156
rect 289996 239260 290052 239316
rect 289772 33628 289828 33684
rect 290780 236908 290836 236964
rect 291564 238252 291620 238308
rect 290332 216300 290388 216356
rect 290108 216188 290164 216244
rect 290108 48524 290164 48580
rect 291452 214396 291508 214452
rect 290332 48412 290388 48468
rect 290556 213164 290612 213220
rect 291788 237468 291844 237524
rect 291788 160076 291844 160132
rect 291676 155932 291732 155988
rect 293244 237580 293300 237636
rect 292572 155596 292628 155652
rect 293132 215852 293188 215908
rect 291564 138572 291620 138628
rect 293244 162092 293300 162148
rect 293468 155484 293524 155540
rect 294924 236908 294980 236964
rect 294364 151004 294420 151060
rect 294812 214284 294868 214340
rect 293132 104076 293188 104132
rect 291452 103852 291508 103908
rect 294924 155708 294980 155764
rect 295036 212492 295092 212548
rect 295260 152796 295316 152852
rect 296940 197372 296996 197428
rect 296940 157276 296996 157332
rect 297164 237356 297220 237412
rect 297164 158844 297220 158900
rect 297276 237244 297332 237300
rect 297276 158732 297332 158788
rect 297052 155372 297108 155428
rect 298732 204092 298788 204148
rect 298620 200844 298676 200900
rect 298508 199164 298564 199220
rect 298396 195692 298452 195748
rect 298508 157388 298564 157444
rect 298844 159404 298900 159460
rect 298956 237804 299012 237860
rect 300412 237916 300468 237972
rect 299740 159292 299796 159348
rect 299964 197708 300020 197764
rect 298956 158956 299012 159012
rect 298732 157500 298788 157556
rect 300188 197260 300244 197316
rect 300076 196476 300132 196532
rect 300412 160748 300468 160804
rect 300524 237468 300580 237524
rect 300076 157724 300132 157780
rect 299964 157164 300020 157220
rect 298620 157052 298676 157108
rect 298396 156940 298452 156996
rect 297948 150780 298004 150836
rect 296156 150220 296212 150276
rect 303324 237804 303380 237860
rect 302428 237356 302484 237412
rect 301532 236908 301588 236964
rect 305116 237468 305172 237524
rect 306012 237244 306068 237300
rect 304220 236908 304276 236964
rect 307804 237916 307860 237972
rect 307356 236908 307412 236964
rect 309036 236908 309092 236964
rect 309596 236908 309652 236964
rect 302764 234892 302820 234948
rect 301644 217868 301700 217924
rect 300972 211596 301028 211652
rect 300636 159180 300692 159236
rect 300860 205772 300916 205828
rect 300860 156828 300916 156884
rect 300524 149548 300580 149604
rect 301196 211484 301252 211540
rect 301084 199052 301140 199108
rect 301084 157612 301140 157668
rect 307244 234780 307300 234836
rect 305004 222908 305060 222964
rect 303884 219548 303940 219604
rect 306124 221228 306180 221284
rect 308364 233212 308420 233268
rect 309484 215964 309540 216020
rect 310492 197932 310548 197988
rect 310604 229964 310660 230020
rect 311388 197820 311444 197876
rect 311724 224812 311780 224868
rect 312284 197484 312340 197540
rect 312844 217756 312900 217812
rect 314076 237804 314132 237860
rect 313180 201068 313236 201124
rect 313964 219436 314020 219492
rect 314972 200956 315028 201012
rect 315084 228172 315140 228228
rect 315868 197596 315924 197652
rect 316204 219324 316260 219380
rect 317660 236908 317716 236964
rect 318444 222796 318500 222852
rect 316764 201180 316820 201236
rect 317324 217644 317380 217700
rect 321244 238028 321300 238084
rect 320348 237916 320404 237972
rect 321804 233100 321860 233156
rect 320684 231308 320740 231364
rect 319452 198156 319508 198212
rect 319564 224700 319620 224756
rect 318556 197148 318612 197204
rect 322140 197260 322196 197316
rect 322924 229740 322980 229796
rect 323932 199276 323988 199332
rect 324044 222572 324100 222628
rect 324828 198044 324884 198100
rect 325164 228060 325220 228116
rect 325276 197148 325332 197204
rect 326284 221116 326340 221172
rect 326620 205772 326676 205828
rect 327404 231196 327460 231252
rect 323820 196476 323876 196532
rect 328412 199164 328468 199220
rect 328524 234668 328580 234724
rect 329308 204092 329364 204148
rect 329644 224588 329700 224644
rect 330204 197708 330260 197764
rect 330764 229852 330820 229908
rect 331100 199052 331156 199108
rect 331884 232988 331940 233044
rect 334236 236908 334292 236964
rect 337372 238028 337428 238084
rect 334684 236908 334740 236964
rect 337148 237916 337204 237972
rect 335244 231084 335300 231140
rect 332892 200844 332948 200900
rect 333004 229628 333060 229684
rect 331996 197372 332052 197428
rect 335132 229404 335188 229460
rect 334124 227948 334180 228004
rect 335132 207452 335188 207508
rect 336924 214620 336980 214676
rect 336812 212604 336868 212660
rect 327516 196476 327572 196532
rect 336364 162428 336420 162484
rect 304332 160524 304388 160580
rect 302876 160412 302932 160468
rect 306572 157836 306628 157892
rect 308140 156940 308196 156996
rect 311276 157724 311332 157780
rect 314412 157500 314468 157556
rect 312844 157388 312900 157444
rect 317548 157612 317604 157668
rect 319116 157276 319172 157332
rect 315980 157164 316036 157220
rect 322252 157836 322308 157892
rect 323820 157164 323876 157220
rect 320684 157052 320740 157108
rect 309708 156828 309764 156884
rect 326956 157500 327012 157556
rect 328524 157388 328580 157444
rect 333228 157724 333284 157780
rect 334796 157612 334852 157668
rect 331660 157276 331716 157332
rect 330092 156940 330148 156996
rect 325388 156828 325444 156884
rect 335916 154476 335972 154532
rect 334684 151340 334740 151396
rect 330092 151228 330148 151284
rect 323372 146188 323428 146244
rect 323372 122556 323428 122612
rect 301196 106988 301252 107044
rect 300972 106876 301028 106932
rect 295036 103964 295092 104020
rect 294812 103180 294868 103236
rect 331772 149660 331828 149716
rect 330876 145516 330932 145572
rect 330876 140252 330932 140308
rect 334684 143612 334740 143668
rect 335132 122668 335188 122724
rect 336364 145404 336420 145460
rect 335916 122668 335972 122724
rect 335132 89852 335188 89908
rect 331772 87612 331828 87668
rect 330092 84700 330148 84756
rect 327516 52892 327572 52948
rect 293580 48636 293636 48692
rect 290556 48300 290612 48356
rect 327516 48636 327572 48692
rect 322252 48524 322308 48580
rect 315084 48412 315140 48468
rect 307916 48300 307972 48356
rect 300748 48188 300804 48244
rect 289996 4844 290052 4900
rect 288092 4620 288148 4676
rect 337036 212716 337092 212772
rect 337148 149436 337204 149492
rect 337260 197932 337316 197988
rect 337596 237804 337652 237860
rect 337596 165452 337652 165508
rect 337372 152348 337428 152404
rect 337260 142604 337316 142660
rect 337036 74844 337092 74900
rect 336924 48636 336980 48692
rect 338940 240492 338996 240548
rect 338604 240380 338660 240436
rect 338604 46284 338660 46340
rect 338716 240268 338772 240324
rect 338828 197820 338884 197876
rect 338828 137676 338884 137732
rect 339724 350140 339780 350196
rect 339724 164108 339780 164164
rect 339836 336028 339892 336084
rect 339612 162764 339668 162820
rect 339948 277004 340004 277060
rect 339948 240156 340004 240212
rect 340060 273868 340116 273924
rect 340060 238476 340116 238532
rect 341068 337260 341124 337316
rect 340284 246652 340340 246708
rect 340956 245308 341012 245364
rect 345212 407260 345268 407316
rect 342748 407036 342804 407092
rect 342748 406700 342804 406756
rect 343532 393148 343588 393204
rect 341852 383068 341908 383124
rect 343196 389004 343252 389060
rect 343084 365036 343140 365092
rect 341180 294252 341236 294308
rect 341852 356076 341908 356132
rect 341292 280476 341348 280532
rect 341180 250012 341236 250068
rect 341292 250348 341348 250404
rect 341292 246876 341348 246932
rect 340396 241554 340452 241556
rect 340396 241502 340398 241554
rect 340398 241502 340450 241554
rect 340450 241502 340452 241554
rect 340396 241500 340452 241502
rect 340956 239484 341012 239540
rect 340508 237692 340564 237748
rect 340284 236236 340340 236292
rect 340396 237580 340452 237636
rect 340172 177100 340228 177156
rect 340284 186508 340340 186564
rect 340956 237580 341012 237636
rect 341068 236348 341124 236404
rect 340508 189196 340564 189252
rect 339836 157052 339892 157108
rect 339948 154476 340004 154532
rect 341852 162652 341908 162708
rect 341964 352492 342020 352548
rect 342972 340844 343028 340900
rect 342636 298956 342692 299012
rect 342524 277228 342580 277284
rect 342412 268716 342468 268772
rect 341964 161084 342020 161140
rect 342076 256172 342132 256228
rect 341068 156828 341124 156884
rect 340396 153468 340452 153524
rect 340396 151340 340452 151396
rect 342188 248220 342244 248276
rect 342188 237692 342244 237748
rect 342188 201068 342244 201124
rect 342188 163772 342244 163828
rect 342300 198156 342356 198212
rect 342300 162204 342356 162260
rect 342300 157164 342356 157220
rect 342300 156828 342356 156884
rect 342076 151116 342132 151172
rect 342524 248444 342580 248500
rect 342412 150668 342468 150724
rect 342524 247772 342580 247828
rect 342524 95676 342580 95732
rect 342748 263788 342804 263844
rect 342748 239708 342804 239764
rect 342860 249452 342916 249508
rect 342860 236012 342916 236068
rect 343308 387212 343364 387268
rect 343420 379708 343476 379764
rect 345212 385756 345268 385812
rect 345548 384412 345604 384468
rect 343532 372204 343588 372260
rect 345436 381276 345492 381332
rect 345324 365932 345380 365988
rect 345212 357868 345268 357924
rect 343980 342636 344036 342692
rect 343868 341740 343924 341796
rect 343644 339948 343700 340004
rect 343420 293132 343476 293188
rect 343532 339052 343588 339108
rect 343308 292460 343364 292516
rect 343196 291340 343252 291396
rect 343084 268716 343140 268772
rect 343196 272748 343252 272804
rect 343308 270956 343364 271012
rect 343420 267372 343476 267428
rect 343644 264572 343700 264628
rect 343532 250348 343588 250404
rect 343420 239820 343476 239876
rect 343308 239260 343364 239316
rect 343196 237916 343252 237972
rect 343532 238700 343588 238756
rect 342972 157276 343028 157332
rect 342748 157052 342804 157108
rect 342748 150332 342804 150388
rect 342636 48412 342692 48468
rect 339500 46508 339556 46564
rect 339388 43260 339444 43316
rect 338940 43148 338996 43204
rect 338716 42812 338772 42868
rect 338492 41244 338548 41300
rect 343756 238588 343812 238644
rect 343644 209916 343700 209972
rect 343644 107324 343700 107380
rect 343868 157724 343924 157780
rect 344092 273644 344148 273700
rect 344092 238924 344148 238980
rect 344428 254828 344484 254884
rect 344540 252588 344596 252644
rect 344540 245084 344596 245140
rect 344652 245196 344708 245252
rect 344652 240268 344708 240324
rect 344428 238588 344484 238644
rect 344316 208348 344372 208404
rect 343980 157612 344036 157668
rect 344204 177212 344260 177268
rect 344204 157500 344260 157556
rect 344316 156940 344372 156996
rect 345100 195804 345156 195860
rect 345100 149212 345156 149268
rect 345436 358540 345492 358596
rect 345324 163660 345380 163716
rect 345436 348908 345492 348964
rect 345772 383852 345828 383908
rect 345772 366156 345828 366212
rect 346892 380604 346948 380660
rect 348572 409948 348628 410004
rect 351260 409388 351316 409444
rect 351148 409276 351204 409332
rect 348684 407932 348740 407988
rect 350588 407820 350644 407876
rect 350364 407708 350420 407764
rect 348684 385868 348740 385924
rect 350252 404348 350308 404404
rect 348572 382844 348628 382900
rect 350364 387436 350420 387492
rect 350476 399980 350532 400036
rect 350252 382396 350308 382452
rect 350364 384524 350420 384580
rect 347004 377468 347060 377524
rect 348572 370412 348628 370468
rect 347004 359660 347060 359716
rect 346780 328300 346836 328356
rect 345548 309036 345604 309092
rect 346108 314860 346164 314916
rect 345548 299068 345604 299124
rect 345996 283836 346052 283892
rect 345884 282156 345940 282212
rect 345772 262332 345828 262388
rect 345548 256956 345604 257012
rect 345660 258636 345716 258692
rect 345436 158620 345492 158676
rect 345548 197484 345604 197540
rect 345212 147532 345268 147588
rect 345660 154476 345716 154532
rect 345884 154252 345940 154308
rect 345772 150444 345828 150500
rect 345548 139356 345604 139412
rect 346892 308588 346948 308644
rect 346444 285292 346500 285348
rect 346220 255724 346276 255780
rect 346220 240156 346276 240212
rect 346332 248444 346388 248500
rect 346668 276332 346724 276388
rect 346444 246764 346500 246820
rect 346556 250348 346612 250404
rect 346332 160972 346388 161028
rect 346108 157836 346164 157892
rect 346668 229292 346724 229348
rect 346556 157388 346612 157444
rect 347004 147644 347060 147700
rect 347228 280476 347284 280532
rect 348012 272972 348068 273028
rect 347788 245196 347844 245252
rect 347900 262892 347956 262948
rect 348012 253932 348068 253988
rect 348012 241500 348068 241556
rect 347900 240492 347956 240548
rect 347228 159516 347284 159572
rect 347340 197596 347396 197652
rect 350252 364140 350308 364196
rect 348572 165004 348628 165060
rect 348684 362348 348740 362404
rect 348796 354284 348852 354340
rect 349020 346220 349076 346276
rect 348796 164220 348852 164276
rect 348908 345324 348964 345380
rect 349580 270060 349636 270116
rect 349468 260204 349524 260260
rect 349356 246876 349412 246932
rect 349244 244860 349300 244916
rect 349020 165116 349076 165172
rect 349132 238588 349188 238644
rect 348908 162876 348964 162932
rect 348684 161980 348740 162036
rect 347340 148652 347396 148708
rect 347116 116732 347172 116788
rect 349244 162428 349300 162484
rect 349132 102172 349188 102228
rect 349580 252588 349636 252644
rect 349468 240380 349524 240436
rect 351148 407036 351204 407092
rect 351260 406700 351316 406756
rect 351148 406588 351204 406644
rect 352044 406588 352100 406644
rect 350588 387324 350644 387380
rect 351820 389788 351876 389844
rect 350476 382732 350532 382788
rect 350588 383068 350644 383124
rect 350588 370636 350644 370692
rect 350812 381388 350868 381444
rect 350364 312508 350420 312564
rect 350476 358764 350532 358820
rect 350252 164444 350308 164500
rect 350364 247884 350420 247940
rect 349356 101388 349412 101444
rect 346892 50204 346948 50260
rect 350476 164332 350532 164388
rect 350588 355180 350644 355236
rect 350700 348012 350756 348068
rect 350924 380716 350980 380772
rect 351820 346444 351876 346500
rect 351932 370636 351988 370692
rect 350924 334348 350980 334404
rect 351260 284396 351316 284452
rect 351260 278908 351316 278964
rect 350812 248220 350868 248276
rect 350924 252028 350980 252084
rect 350700 164556 350756 164612
rect 350588 162540 350644 162596
rect 350812 151116 350868 151172
rect 350812 149660 350868 149716
rect 350812 146076 350868 146132
rect 350924 110124 350980 110180
rect 351036 249452 351092 249508
rect 351260 236460 351316 236516
rect 351372 264684 351428 264740
rect 351372 234556 351428 234612
rect 351484 264572 351540 264628
rect 351820 261212 351876 261268
rect 351820 256956 351876 257012
rect 351820 245196 351876 245252
rect 351820 239484 351876 239540
rect 351484 208348 351540 208404
rect 351148 200732 351204 200788
rect 351148 171276 351204 171332
rect 351148 170380 351204 170436
rect 351260 196364 351316 196420
rect 351260 195244 351316 195300
rect 351260 167692 351316 167748
rect 355516 408044 355572 408100
rect 353724 407596 353780 407652
rect 352716 407148 352772 407204
rect 352156 382732 352212 382788
rect 352156 381388 352212 381444
rect 352268 406700 352324 406756
rect 352156 380492 352212 380548
rect 352156 352492 352212 352548
rect 352604 404908 352660 404964
rect 352604 388780 352660 388836
rect 352380 384748 352436 384804
rect 352380 340396 352436 340452
rect 352492 377468 352548 377524
rect 352380 312508 352436 312564
rect 352380 310156 352436 310212
rect 352380 309036 352436 309092
rect 352380 304108 352436 304164
rect 352268 268716 352324 268772
rect 352044 261772 352100 261828
rect 352156 233436 352212 233492
rect 352380 256956 352436 257012
rect 352380 255724 352436 255780
rect 352044 225484 352100 225540
rect 352044 181356 352100 181412
rect 352156 219436 352212 219492
rect 352268 207340 352324 207396
rect 352044 178444 352100 178500
rect 352380 198156 352436 198212
rect 352268 173628 352324 173684
rect 352268 173068 352324 173124
rect 352044 163884 352100 163940
rect 351932 154364 351988 154420
rect 352380 171276 352436 171332
rect 353612 404460 353668 404516
rect 355180 407484 355236 407540
rect 353724 385644 353780 385700
rect 353836 399532 353892 399588
rect 354844 397404 354900 397460
rect 354732 394156 354788 394212
rect 354060 393932 354116 393988
rect 354956 397292 355012 397348
rect 355068 397068 355124 397124
rect 355068 394156 355124 394212
rect 355404 406476 355460 406532
rect 355292 403004 355348 403060
rect 355292 398076 355348 398132
rect 354956 391132 355012 391188
rect 354844 390908 354900 390964
rect 355180 393708 355236 393764
rect 355180 392588 355236 392644
rect 355068 390684 355124 390740
rect 354732 387884 354788 387940
rect 354060 382620 354116 382676
rect 353836 382508 353892 382564
rect 355404 397180 355460 397236
rect 367612 408156 367668 408212
rect 372764 408044 372820 408100
rect 379596 408604 379652 408660
rect 379596 408156 379652 408212
rect 377916 407932 377972 407988
rect 383068 407484 383124 407540
rect 383292 407484 383348 407540
rect 362460 407260 362516 407316
rect 357308 404908 357364 404964
rect 398524 407820 398580 407876
rect 399756 407820 399812 407876
rect 393372 407596 393428 407652
rect 397292 407596 397348 407652
rect 388220 404796 388276 404852
rect 383292 399756 383348 399812
rect 371980 397404 372036 397460
rect 361228 396732 361284 396788
rect 361228 395164 361284 395220
rect 358204 395052 358260 395108
rect 365148 395052 365204 395108
rect 386428 397292 386484 397348
rect 379820 395052 379876 395108
rect 393148 397180 393204 397236
rect 408828 407708 408884 407764
rect 403676 407372 403732 407428
rect 403900 407372 403956 407428
rect 399756 404684 399812 404740
rect 419132 407820 419188 407876
rect 413980 406476 414036 406532
rect 419356 407708 419412 407764
rect 403900 402892 403956 402948
rect 414092 399868 414148 399924
rect 414092 397404 414148 397460
rect 406812 397068 406868 397124
rect 397292 396284 397348 396340
rect 400204 396956 400260 397012
rect 403116 396508 403172 396564
rect 413756 396508 413812 396564
rect 430108 408380 430164 408436
rect 430108 408044 430164 408100
rect 429436 407484 429492 407540
rect 424284 407372 424340 407428
rect 424956 407372 425012 407428
rect 421596 401660 421652 401716
rect 439740 408156 439796 408212
rect 444892 407820 444948 407876
rect 455196 407708 455252 407764
rect 450044 407596 450100 407652
rect 434588 404572 434644 404628
rect 445116 407484 445172 407540
rect 424956 399644 425012 399700
rect 442092 399980 442148 400036
rect 421596 397292 421652 397348
rect 427644 397404 427700 397460
rect 419356 396172 419412 396228
rect 420700 396844 420756 396900
rect 435148 397292 435204 397348
rect 429212 396844 429268 396900
rect 403116 394716 403172 394772
rect 445116 399420 445172 399476
rect 448588 396844 448644 396900
rect 455308 396508 455364 396564
rect 460348 395948 460404 396004
rect 464492 406588 464548 406644
rect 465500 406588 465556 406644
rect 464492 395836 464548 395892
rect 466172 406028 466228 406084
rect 466172 395836 466228 395892
rect 469196 398188 469252 398244
rect 472892 406588 472948 406644
rect 472892 403004 472948 403060
rect 470652 395724 470708 395780
rect 486108 408044 486164 408100
rect 496412 407596 496468 407652
rect 501564 407484 501620 407540
rect 504700 408268 504756 408324
rect 490588 406700 490644 406756
rect 480956 404236 481012 404292
rect 475804 395612 475860 395668
rect 497644 401548 497700 401604
rect 511868 410060 511924 410116
rect 522172 407484 522228 407540
rect 527324 407484 527380 407540
rect 517020 407372 517076 407428
rect 529340 402780 529396 402836
rect 529452 489132 529508 489188
rect 529564 479836 529620 479892
rect 529564 402444 529620 402500
rect 529676 470428 529732 470484
rect 529452 401324 529508 401380
rect 506716 399532 506772 399588
rect 562604 590492 562660 590548
rect 584668 590156 584724 590212
rect 540540 575484 540596 575540
rect 537628 546252 537684 546308
rect 532588 541548 532644 541604
rect 530908 513324 530964 513380
rect 529788 409276 529844 409332
rect 529900 465612 529956 465668
rect 529676 399308 529732 399364
rect 529900 399196 529956 399252
rect 530012 460796 530068 460852
rect 530012 399084 530068 399140
rect 530124 414540 530180 414596
rect 530124 398972 530180 399028
rect 518028 396732 518084 396788
rect 483868 394940 483924 394996
rect 525532 394940 525588 394996
rect 490812 394828 490868 394884
rect 476924 394716 476980 394772
rect 511644 394716 511700 394772
rect 429212 394604 429268 394660
rect 463036 394604 463092 394660
rect 531020 452172 531076 452228
rect 531244 423948 531300 424004
rect 531020 405916 531076 405972
rect 531132 419244 531188 419300
rect 531244 405692 531300 405748
rect 534268 536844 534324 536900
rect 532700 456876 532756 456932
rect 532700 409164 532756 409220
rect 532812 447468 532868 447524
rect 532924 438060 532980 438116
rect 533036 433356 533092 433412
rect 534380 532140 534436 532196
rect 535948 522732 536004 522788
rect 534380 409052 534436 409108
rect 534492 503916 534548 503972
rect 534268 406252 534324 406308
rect 533036 405804 533092 405860
rect 532924 404460 532980 404516
rect 532812 404348 532868 404404
rect 532588 404124 532644 404180
rect 534492 401212 534548 401268
rect 534604 494508 534660 494564
rect 534604 400988 534660 401044
rect 534716 485100 534772 485156
rect 535948 402668 536004 402724
rect 536060 518028 536116 518084
rect 536060 402556 536116 402612
rect 536172 508620 536228 508676
rect 536172 401100 536228 401156
rect 536284 499212 536340 499268
rect 545132 482860 545188 482916
rect 537628 406140 537684 406196
rect 540092 456428 540148 456484
rect 587132 443212 587188 443268
rect 545132 409836 545188 409892
rect 560252 409948 560308 410004
rect 540092 402332 540148 402388
rect 536284 400876 536340 400932
rect 534716 400764 534772 400820
rect 531132 400652 531188 400708
rect 539308 397740 539364 397796
rect 531804 396620 531860 396676
rect 546252 396844 546308 396900
rect 553196 396620 553252 396676
rect 587132 406588 587188 406644
rect 583884 404012 583940 404068
rect 583772 403228 583828 403284
rect 574028 396844 574084 396900
rect 567084 396508 567140 396564
rect 580972 396732 581028 396788
rect 582988 395836 583044 395892
rect 582988 394828 583044 394884
rect 583660 394828 583716 394884
rect 530908 394492 530964 394548
rect 355516 390572 355572 390628
rect 355404 387772 355460 387828
rect 355292 382284 355348 382340
rect 353612 382172 353668 382228
rect 353612 366828 353668 366884
rect 353500 310156 353556 310212
rect 352716 245196 352772 245252
rect 352828 272076 352884 272132
rect 352828 238588 352884 238644
rect 353500 236796 353556 236852
rect 352716 213388 352772 213444
rect 352716 175756 352772 175812
rect 353500 173852 353556 173908
rect 352380 165340 352436 165396
rect 352716 171052 352772 171108
rect 352604 162316 352660 162372
rect 352604 154364 352660 154420
rect 352604 153692 352660 153748
rect 352268 153020 352324 153076
rect 352380 145516 352436 145572
rect 351036 104300 351092 104356
rect 351148 58716 351204 58772
rect 353500 165564 353556 165620
rect 355404 361452 355460 361508
rect 353612 156156 353668 156212
rect 353724 353388 353780 353444
rect 355292 351596 355348 351652
rect 353836 349804 353892 349860
rect 354508 338156 354564 338212
rect 354060 316988 354116 317044
rect 353948 298060 354004 298116
rect 353948 272076 354004 272132
rect 353836 160972 353892 161028
rect 353948 252028 354004 252084
rect 353724 147196 353780 147252
rect 354396 284732 354452 284788
rect 354284 273868 354340 273924
rect 354060 234444 354116 234500
rect 354060 234108 354116 234164
rect 354172 238588 354228 238644
rect 354060 183260 354116 183316
rect 354172 173852 354228 173908
rect 354172 173628 354228 173684
rect 354172 165228 354228 165284
rect 354284 163996 354340 164052
rect 354060 159516 354116 159572
rect 354620 287308 354676 287364
rect 355068 279356 355124 279412
rect 355068 238252 355124 238308
rect 354620 234332 354676 234388
rect 354620 234108 354676 234164
rect 354508 177212 354564 177268
rect 354732 166236 354788 166292
rect 355180 183372 355236 183428
rect 354396 107212 354452 107268
rect 353948 99036 354004 99092
rect 352716 58716 352772 58772
rect 351148 57148 351204 57204
rect 351148 52892 351204 52948
rect 350364 50092 350420 50148
rect 345996 48188 346052 48244
rect 355404 161196 355460 161252
rect 355516 238252 355572 238308
rect 486444 165564 486500 165620
rect 422716 165340 422772 165396
rect 365820 165116 365876 165172
rect 358204 162876 358260 162932
rect 379820 164556 379876 164612
rect 372092 162428 372148 162484
rect 399868 164108 399924 164164
rect 393484 160972 393540 161028
rect 386540 158620 386596 158676
rect 355516 155260 355572 155316
rect 366268 155260 366324 155316
rect 355292 147084 355348 147140
rect 414316 161084 414372 161140
rect 420812 164668 420868 164724
rect 421820 163884 421876 163940
rect 420812 154252 420868 154308
rect 421820 153916 421876 153972
rect 422492 156940 422548 156996
rect 422492 154252 422548 154308
rect 421372 147196 421428 147252
rect 407484 147084 407540 147140
rect 366268 145852 366324 145908
rect 401884 146972 401940 147028
rect 400316 145292 400372 145348
rect 386092 107324 386148 107380
rect 376572 104076 376628 104132
rect 372988 103740 373044 103796
rect 374668 103180 374724 103236
rect 383964 103964 384020 104020
rect 381388 103852 381444 103908
rect 378028 103628 378084 103684
rect 379708 103292 379764 103348
rect 383180 103516 383236 103572
rect 390796 106988 390852 107044
rect 387100 103404 387156 103460
rect 389228 103180 389284 103236
rect 393932 106876 393988 106932
rect 392364 103292 392420 103348
rect 395500 106764 395556 106820
rect 396508 104076 396564 104132
rect 398188 104076 398244 104132
rect 421820 144620 421876 144676
rect 421708 144508 421764 144564
rect 406588 138572 406644 138628
rect 403452 133532 403508 133588
rect 415996 135212 416052 135268
rect 408156 131964 408212 132020
rect 404908 106652 404964 106708
rect 406588 104972 406644 105028
rect 406588 102508 406644 102564
rect 414428 131852 414484 131908
rect 411292 125132 411348 125188
rect 408940 102508 408996 102564
rect 412860 115052 412916 115108
rect 366268 93436 366324 93492
rect 366268 91420 366324 91476
rect 420028 81564 420084 81620
rect 367836 58268 367892 58324
rect 367836 57148 367892 57204
rect 367948 50988 368004 51044
rect 419356 52108 419412 52164
rect 419356 49756 419412 49812
rect 420028 48076 420084 48132
rect 420140 77308 420196 77364
rect 421932 122556 421988 122612
rect 421932 87164 421988 87220
rect 421820 82236 421876 82292
rect 421708 77308 421764 77364
rect 420252 72380 420308 72436
rect 422268 72380 422324 72436
rect 421932 68796 421988 68852
rect 421932 67452 421988 67508
rect 420252 49980 420308 50036
rect 420364 62524 420420 62580
rect 420364 49868 420420 49924
rect 421708 57596 421764 57652
rect 466172 165340 466228 165396
rect 422716 154140 422772 154196
rect 422940 165228 422996 165284
rect 422940 154028 422996 154084
rect 423164 164892 423220 164948
rect 427644 164220 427700 164276
rect 448588 162764 448644 162820
rect 441868 162652 441924 162708
rect 435148 162540 435204 162596
rect 462364 164332 462420 164388
rect 464940 164108 464996 164164
rect 463596 163884 463652 163940
rect 458220 162428 458276 162484
rect 457772 161308 457828 161364
rect 423164 154364 423220 154420
rect 456092 147532 456148 147588
rect 458108 159852 458164 159908
rect 457884 159628 457940 159684
rect 457996 157948 458052 158004
rect 459452 154588 459508 154644
rect 458220 147644 458276 147700
rect 458556 148316 458612 148372
rect 458108 146076 458164 146132
rect 458556 142604 458612 142660
rect 457996 141036 458052 141092
rect 463596 154252 463652 154308
rect 477036 162876 477092 162932
rect 481068 163996 481124 164052
rect 469308 162428 469364 162484
rect 464940 154140 464996 154196
rect 479724 159852 479780 159908
rect 470316 157836 470372 157892
rect 466060 154028 466116 154084
rect 467628 154364 467684 154420
rect 468972 153916 469028 153972
rect 473788 156940 473844 156996
rect 473004 154700 473060 154756
rect 470316 153916 470372 153972
rect 471660 153916 471716 153972
rect 470316 152908 470372 152964
rect 471660 151340 471716 151396
rect 473788 152908 473844 152964
rect 474348 156268 474404 156324
rect 475692 152908 475748 152964
rect 478380 151228 478436 151284
rect 477036 149884 477092 149940
rect 483980 161196 484036 161252
rect 482412 158060 482468 158116
rect 483756 154476 483812 154532
rect 485100 152908 485156 152964
rect 557900 165452 557956 165508
rect 490700 161980 490756 162036
rect 495852 163212 495908 163268
rect 487788 154476 487844 154532
rect 488908 154476 488964 154532
rect 490476 154476 490532 154532
rect 491820 154476 491876 154532
rect 493164 154476 493220 154532
rect 494732 153244 494788 153300
rect 494508 152908 494564 152964
rect 470316 149660 470372 149716
rect 553308 165004 553364 165060
rect 504028 164444 504084 164500
rect 497868 162876 497924 162932
rect 502796 162316 502852 162372
rect 497196 161644 497252 161700
rect 508732 160188 508788 160244
rect 502796 154476 502852 154532
rect 506604 154476 506660 154532
rect 500108 154028 500164 154084
rect 497308 153580 497364 153636
rect 497308 152684 497364 152740
rect 498540 152908 498596 152964
rect 499884 152908 499940 152964
rect 494732 149660 494788 149716
rect 501228 153804 501284 153860
rect 500668 153356 500724 153412
rect 500668 150892 500724 150948
rect 502572 153692 502628 153748
rect 505260 153468 505316 153524
rect 503916 153020 503972 153076
rect 505596 152908 505652 152964
rect 505596 152572 505652 152628
rect 510748 155932 510804 155988
rect 508732 154476 508788 154532
rect 510636 155820 510692 155876
rect 509292 153580 509348 153636
rect 507276 153468 507332 153524
rect 507276 150780 507332 150836
rect 507948 152236 508004 152292
rect 510748 153692 510804 153748
rect 517916 163660 517972 163716
rect 520044 162092 520100 162148
rect 516012 160636 516068 160692
rect 514668 160300 514724 160356
rect 513324 160076 513380 160132
rect 511532 150668 511588 150724
rect 511980 154476 512036 154532
rect 518700 153244 518756 153300
rect 517356 152124 517412 152180
rect 522508 159404 522564 159460
rect 532364 162876 532420 162932
rect 539308 162876 539364 162932
rect 546476 162876 546532 162932
rect 557004 164668 557060 164724
rect 554652 162204 554708 162260
rect 540876 160524 540932 160580
rect 525420 156156 525476 156212
rect 532588 159292 532644 159348
rect 525420 155708 525476 155764
rect 522508 153804 522564 153860
rect 524076 154028 524132 154084
rect 522732 153356 522788 153412
rect 520828 153244 520884 153300
rect 520828 151004 520884 151060
rect 521388 152908 521444 152964
rect 524188 152908 524244 152964
rect 524188 150220 524244 150276
rect 528108 155596 528164 155652
rect 526764 153692 526820 153748
rect 529452 155484 529508 155540
rect 535948 159180 536004 159236
rect 532588 154476 532644 154532
rect 534828 155372 534884 155428
rect 530796 153244 530852 153300
rect 533484 153020 533540 153076
rect 532140 152908 532196 152964
rect 539196 159068 539252 159124
rect 535948 154364 536004 154420
rect 538860 154476 538916 154532
rect 537516 153804 537572 153860
rect 536172 153468 536228 153524
rect 539196 154252 539252 154308
rect 540204 154364 540260 154420
rect 550956 160412 551012 160468
rect 544236 158956 544292 159012
rect 542892 158844 542948 158900
rect 540876 153692 540932 153748
rect 541548 154252 541604 154308
rect 548268 158732 548324 158788
rect 545580 152012 545636 152068
rect 549612 153692 549668 153748
rect 554540 157724 554596 157780
rect 554428 150332 554484 150388
rect 500108 149660 500164 149716
rect 546924 149548 546980 149604
rect 459452 139356 459508 139412
rect 457884 139132 457940 139188
rect 457772 137676 457828 137732
rect 554540 140476 554596 140532
rect 554428 130956 554484 131012
rect 556892 161420 556948 161476
rect 555100 161308 555156 161364
rect 554988 157948 555044 158004
rect 554876 148652 554932 148708
rect 554652 125916 554708 125972
rect 554764 148316 554820 148372
rect 554876 120204 554932 120260
rect 554764 112140 554820 112196
rect 556332 159628 556388 159684
rect 555212 157612 555268 157668
rect 556220 157276 556276 157332
rect 555212 141372 555268 141428
rect 556108 157164 556164 157220
rect 556220 138236 556276 138292
rect 556108 131964 556164 132020
rect 555100 113148 555156 113204
rect 556780 157500 556836 157556
rect 556444 154588 556500 154644
rect 556556 149772 556612 149828
rect 556668 149212 556724 149268
rect 556780 133532 556836 133588
rect 556668 124124 556724 124180
rect 556556 120988 556612 121044
rect 556444 114716 556500 114772
rect 556332 110012 556388 110068
rect 554988 108780 555044 108836
rect 554316 104076 554372 104132
rect 458556 99932 458612 99988
rect 457660 98700 457716 98756
rect 449372 98364 449428 98420
rect 449372 97804 449428 97860
rect 457660 92652 457716 92708
rect 458444 97804 458500 97860
rect 458444 72156 458500 72212
rect 423164 68796 423220 68852
rect 422940 62524 422996 62580
rect 422716 57596 422772 57652
rect 554316 99932 554372 99988
rect 557788 149436 557844 149492
rect 567756 162764 567812 162820
rect 581196 164668 581252 164724
rect 574476 162652 574532 162708
rect 560700 162540 560756 162596
rect 558348 159740 558404 159796
rect 558236 152348 558292 152404
rect 557900 142940 557956 142996
rect 558012 151116 558068 151172
rect 557788 127260 557844 127316
rect 558012 88060 558068 88116
rect 558124 147868 558180 147924
rect 558236 128828 558292 128884
rect 558124 86492 558180 86548
rect 583772 377132 583828 377188
rect 583660 157836 583716 157892
rect 559468 157388 559524 157444
rect 558460 152796 558516 152852
rect 559580 157052 559636 157108
rect 590604 394828 590660 394884
rect 584668 393148 584724 393204
rect 590492 392812 590548 392868
rect 590604 364140 590660 364196
rect 590492 324492 590548 324548
rect 590492 284620 590548 284676
rect 590492 165340 590548 165396
rect 590604 244972 590660 245028
rect 590604 164108 590660 164164
rect 590828 205324 590884 205380
rect 590828 163884 590884 163940
rect 584668 162764 584724 162820
rect 583884 156940 583940 156996
rect 559580 136668 559636 136724
rect 559468 135100 559524 135156
rect 558460 83356 558516 83412
rect 558348 78652 558404 78708
rect 557004 75516 557060 75572
rect 556892 70812 556948 70868
rect 590492 73164 590548 73220
rect 557788 69244 557844 69300
rect 458556 54796 458612 54852
rect 554428 56028 554484 56084
rect 422492 52668 422548 52724
rect 421932 49644 421988 49700
rect 421708 49532 421764 49588
rect 420140 47964 420196 48020
rect 355180 45164 355236 45220
rect 558348 66108 558404 66164
rect 558124 62972 558180 63028
rect 557788 50316 557844 50372
rect 557900 59836 557956 59892
rect 557900 50204 557956 50260
rect 558012 58268 558068 58324
rect 558236 61404 558292 61460
rect 558236 50092 558292 50148
rect 558124 48412 558180 48468
rect 558012 48300 558068 48356
rect 558348 48188 558404 48244
rect 590604 59948 590660 60004
rect 590604 48636 590660 48692
rect 590492 45276 590548 45332
rect 554428 45164 554484 45220
rect 343756 41356 343812 41412
rect 343532 41132 343588 41188
rect 336812 4284 336868 4340
rect 580860 4956 580916 5012
rect 284956 4172 285012 4228
rect 278012 4060 278068 4116
rect 582540 4284 582596 4340
rect 584444 4172 584500 4228
<< metal3 >>
rect 201506 591276 201516 591332
rect 201572 591276 231644 591332
rect 231700 591276 231710 591332
rect 203186 591164 203196 591220
rect 203252 591164 297836 591220
rect 297892 591164 297902 591220
rect 208114 591052 208124 591108
rect 208180 591052 319900 591108
rect 319956 591052 319966 591108
rect 204642 590940 204652 590996
rect 204708 590940 364028 590996
rect 364084 590940 364094 590996
rect 121538 590828 121548 590884
rect 121604 590828 168812 590884
rect 168868 590828 168878 590884
rect 208002 590828 208012 590884
rect 208068 590828 386092 590884
rect 386148 590828 386158 590884
rect 99474 590716 99484 590772
rect 99540 590716 153692 590772
rect 153748 590716 153758 590772
rect 206322 590716 206332 590772
rect 206388 590716 430220 590772
rect 430276 590716 430286 590772
rect 55346 590604 55356 590660
rect 55412 590604 152012 590660
rect 152068 590604 152078 590660
rect 208226 590604 208236 590660
rect 208292 590604 496412 590660
rect 496468 590604 496478 590660
rect 518690 590604 518700 590660
rect 518756 590604 529788 590660
rect 529844 590604 529854 590660
rect 33282 590492 33292 590548
rect 33348 590492 155372 590548
rect 155428 590492 155438 590548
rect 186386 590492 186396 590548
rect 186452 590492 562604 590548
rect 562660 590492 562670 590548
rect 444322 590156 444332 590212
rect 444388 590156 452284 590212
rect 452340 590156 452350 590212
rect 584658 590156 584668 590212
rect 584724 590156 584762 590212
rect 189746 588812 189756 588868
rect 189812 588812 408268 588868
rect 408324 588812 408334 588868
rect 595560 588644 597000 588840
rect 590482 588588 590492 588644
rect 590548 588616 597000 588644
rect 590548 588588 595672 588616
rect -960 587188 480 587384
rect -960 587160 157052 587188
rect 392 587132 157052 587160
rect 157108 587132 157118 587188
rect 77298 583772 77308 583828
rect 77364 583772 173852 583828
rect 173908 583772 173918 583828
rect 143378 582092 143388 582148
rect 143444 582092 170492 582148
rect 170548 582092 170558 582148
rect 183026 578732 183036 578788
rect 183092 578732 209580 578788
rect 209636 578732 209646 578788
rect 189634 577052 189644 577108
rect 189700 577052 341964 577108
rect 342020 577052 342030 577108
rect 184706 575484 184716 575540
rect 184772 575484 540540 575540
rect 540596 575484 540606 575540
rect 595560 575428 597000 575624
rect 189298 575372 189308 575428
rect 189364 575400 597000 575428
rect 189364 575372 595672 575400
rect 181346 573692 181356 573748
rect 181412 573692 590492 573748
rect 590548 573692 590558 573748
rect -960 573076 480 573272
rect -960 573048 57932 573076
rect 392 573020 57932 573048
rect 57988 573020 57998 573076
rect 189522 572012 189532 572068
rect 189588 572012 474348 572068
rect 474404 572012 474414 572068
rect 189410 570332 189420 570388
rect 189476 570332 275772 570388
rect 275828 570332 275838 570388
rect 209458 568652 209468 568708
rect 209524 568652 253708 568708
rect 253764 568652 253774 568708
rect 183026 567868 183036 567924
rect 183092 567868 590604 567924
rect 590660 567868 590670 567924
rect 186274 566076 186284 566132
rect 186340 566076 187516 566132
rect 187572 566076 187582 566132
rect 187954 565068 187964 565124
rect 188020 565068 190120 565124
rect 529928 565068 532924 565124
rect 532980 565068 532990 565124
rect 595560 562212 597000 562408
rect 590482 562156 590492 562212
rect 590548 562184 597000 562212
rect 590548 562156 595672 562184
rect 529928 560364 535948 560420
rect 536004 560364 536014 560420
rect -960 558964 480 559160
rect -960 558936 4172 558964
rect 392 558908 4172 558936
rect 4228 558908 4238 558964
rect 187954 557900 187964 557956
rect 188020 557900 190120 557956
rect 529928 555660 532700 555716
rect 532756 555660 532766 555716
rect 529928 550956 537628 551012
rect 537684 550956 537694 551012
rect 186386 550732 186396 550788
rect 186452 550732 190120 550788
rect 590594 549164 590604 549220
rect 590660 549192 595672 549220
rect 590660 549164 597000 549192
rect 595560 548968 597000 549164
rect 529928 546252 537628 546308
rect 537684 546252 537694 546308
rect -960 544852 480 545048
rect -960 544824 7532 544852
rect 392 544796 7532 544824
rect 7588 544796 7598 544852
rect 186162 543564 186172 543620
rect 186228 543564 190120 543620
rect 529928 541548 532588 541604
rect 532644 541548 532654 541604
rect 529928 536844 534268 536900
rect 534324 536844 534334 536900
rect 187842 536396 187852 536452
rect 187908 536396 190120 536452
rect 595560 535780 597000 535976
rect 543442 535724 543452 535780
rect 543508 535752 597000 535780
rect 543508 535724 595672 535752
rect 529928 532140 534380 532196
rect 534436 532140 534446 532196
rect -960 530740 480 530936
rect -960 530712 56252 530740
rect 392 530684 56252 530712
rect 56308 530684 56318 530740
rect 186050 529228 186060 529284
rect 186116 529228 190120 529284
rect 529340 526820 529396 527464
rect 529330 526764 529340 526820
rect 529396 526764 529406 526820
rect 529928 522732 535948 522788
rect 536004 522732 536014 522788
rect 595560 522564 597000 522760
rect 590706 522508 590716 522564
rect 590772 522536 597000 522564
rect 590772 522508 595672 522536
rect 189522 522060 189532 522116
rect 189588 522060 190120 522116
rect 529928 518028 536060 518084
rect 536116 518028 536126 518084
rect -960 516628 480 516824
rect -960 516600 4284 516628
rect 392 516572 4284 516600
rect 4340 516572 4350 516628
rect 187730 514892 187740 514948
rect 187796 514892 190120 514948
rect 529928 513324 530908 513380
rect 530964 513324 530974 513380
rect 595560 509348 597000 509544
rect 590594 509292 590604 509348
rect 590660 509320 597000 509348
rect 590660 509292 595672 509320
rect 529928 508620 536172 508676
rect 536228 508620 536238 508676
rect 187282 507724 187292 507780
rect 187348 507724 190120 507780
rect 529928 503916 534492 503972
rect 534548 503916 534558 503972
rect -960 502516 480 502712
rect -960 502488 4172 502516
rect 392 502460 4172 502488
rect 4228 502460 4238 502516
rect 183922 500556 183932 500612
rect 183988 500556 190120 500612
rect 529928 499212 536284 499268
rect 536340 499212 536350 499268
rect 595560 496132 597000 496328
rect 541762 496076 541772 496132
rect 541828 496104 597000 496132
rect 541828 496076 595672 496104
rect 529928 494508 534604 494564
rect 534660 494508 534670 494564
rect 187394 493388 187404 493444
rect 187460 493388 190120 493444
rect 529452 489188 529508 489832
rect 529442 489132 529452 489188
rect 529508 489132 529518 489188
rect -960 488404 480 488600
rect -960 488376 14252 488404
rect 392 488348 14252 488376
rect 14308 488348 14318 488404
rect 187506 486220 187516 486276
rect 187572 486220 190120 486276
rect 529928 485100 534716 485156
rect 534772 485100 534782 485156
rect 595560 482916 597000 483112
rect 545122 482860 545132 482916
rect 545188 482888 597000 482916
rect 545188 482860 595672 482888
rect 529564 479892 529620 480424
rect 529554 479836 529564 479892
rect 529620 479836 529630 479892
rect 187730 479052 187740 479108
rect 187796 479052 190120 479108
rect 529928 475692 534268 475748
rect 534324 475692 534334 475748
rect -960 474292 480 474488
rect -960 474264 4172 474292
rect 392 474236 4172 474264
rect 4228 474236 4238 474292
rect 187058 471884 187068 471940
rect 187124 471884 190120 471940
rect 4162 471212 4172 471268
rect 4228 471212 178892 471268
rect 178948 471212 178958 471268
rect 529676 470484 529732 471016
rect 529666 470428 529676 470484
rect 529732 470428 529742 470484
rect 595560 469700 597000 469896
rect 590818 469644 590828 469700
rect 590884 469672 597000 469700
rect 590884 469644 595672 469672
rect 4162 469532 4172 469588
rect 4228 469532 150332 469588
rect 150388 469532 150398 469588
rect 4162 467852 4172 467908
rect 4228 467852 172172 467908
rect 172228 467852 172238 467908
rect 4274 466172 4284 466228
rect 4340 466172 175532 466228
rect 175588 466172 175598 466228
rect 529900 465668 529956 466312
rect 529890 465612 529900 465668
rect 529956 465612 529966 465668
rect 187618 464716 187628 464772
rect 187684 464716 190120 464772
rect 529900 460852 529956 461608
rect 529900 460796 530012 460852
rect 530068 460796 530078 460852
rect -960 460180 480 460376
rect -960 460152 93212 460180
rect 392 460124 93212 460152
rect 93268 460124 93278 460180
rect 187842 457548 187852 457604
rect 187908 457548 190120 457604
rect 529928 456876 532700 456932
rect 532756 456876 532766 456932
rect 595560 456484 597000 456680
rect 540082 456428 540092 456484
rect 540148 456456 597000 456484
rect 540148 456428 595672 456456
rect 529928 452172 531020 452228
rect 531076 452172 531086 452228
rect 187282 450380 187292 450436
rect 187348 450380 190120 450436
rect 529928 447468 532812 447524
rect 532868 447468 532878 447524
rect -960 446068 480 446264
rect -960 446040 160412 446068
rect 392 446012 160412 446040
rect 160468 446012 160478 446068
rect 595560 443268 597000 443464
rect 187394 443212 187404 443268
rect 187460 443212 190120 443268
rect 587122 443212 587132 443268
rect 587188 443240 597000 443268
rect 587188 443212 595672 443240
rect 529928 442764 532812 442820
rect 532868 442764 532878 442820
rect 529928 438060 532924 438116
rect 532980 438060 532990 438116
rect 187618 436044 187628 436100
rect 187684 436044 190120 436100
rect 529928 433356 533036 433412
rect 533092 433356 533102 433412
rect -960 431956 480 432152
rect -960 431928 167132 431956
rect 392 431900 167132 431928
rect 167188 431900 167198 431956
rect 595560 430164 597000 430248
rect 590930 430108 590940 430164
rect 590996 430108 597000 430164
rect 595560 430024 597000 430108
rect 168802 428876 168812 428932
rect 168868 428876 190120 428932
rect 529218 428652 529228 428708
rect 529284 428652 529294 428708
rect 529928 423948 531244 424004
rect 531300 423948 531310 424004
rect 189410 421708 189420 421764
rect 189476 421708 190120 421764
rect 529928 419244 531132 419300
rect 531188 419244 531198 419300
rect -960 417844 480 418040
rect -960 417816 4172 417844
rect 392 417788 4172 417816
rect 4228 417788 4238 417844
rect 66322 417564 66332 417620
rect 66388 417564 88172 417620
rect 88228 417564 88238 417620
rect 68562 417452 68572 417508
rect 68628 417452 91532 417508
rect 91588 417452 91598 417508
rect 73042 417340 73052 417396
rect 73108 417340 85036 417396
rect 85092 417340 85102 417396
rect 70802 417228 70812 417284
rect 70868 417228 180572 417284
rect 180628 417228 180638 417284
rect 75282 417116 75292 417172
rect 75348 417116 86492 417172
rect 86548 417116 86558 417172
rect 64082 417004 64092 417060
rect 64148 417004 85260 417060
rect 85316 417004 85326 417060
rect 79762 416892 79772 416948
rect 79828 416892 86716 416948
rect 86772 416892 86782 416948
rect 595560 416836 597000 417032
rect 82002 416780 82012 416836
rect 82068 416780 177212 416836
rect 177268 416780 177278 416836
rect 540082 416780 540092 416836
rect 540148 416808 597000 416836
rect 540148 416780 595672 416808
rect 77522 416668 77532 416724
rect 77588 416668 84812 416724
rect 84868 416668 84878 416724
rect 188066 414540 188076 414596
rect 188132 414540 190120 414596
rect 529928 414540 530124 414596
rect 530180 414540 530190 414596
rect 61814 413308 61852 413364
rect 61908 413308 61918 413364
rect 83944 411964 185612 412020
rect 185668 411964 185678 412020
rect 355394 410060 355404 410116
rect 355460 410060 511868 410116
rect 511924 410060 511934 410116
rect 348562 409948 348572 410004
rect 348628 409948 560252 410004
rect 560308 409948 560318 410004
rect 228498 409836 228508 409892
rect 228564 409836 545132 409892
rect 545188 409836 545198 409892
rect 83906 409724 83916 409780
rect 83972 409724 310940 409780
rect 310996 409724 311006 409780
rect 93202 409612 93212 409668
rect 93268 409612 305788 409668
rect 305844 409612 305854 409668
rect 152002 409500 152012 409556
rect 152068 409500 283948 409556
rect 284004 409500 285180 409556
rect 285236 409500 285246 409556
rect 168802 409388 168812 409444
rect 168868 409388 280476 409444
rect 280532 409388 280542 409444
rect 351250 409388 351260 409444
rect 351316 409388 444332 409444
rect 444388 409388 444398 409444
rect 187954 409276 187964 409332
rect 188020 409276 341180 409332
rect 341236 409276 341246 409332
rect 351138 409276 351148 409332
rect 351204 409276 529788 409332
rect 529844 409276 529854 409332
rect 289734 409164 289772 409220
rect 289828 409164 289838 409220
rect 298162 409164 298172 409220
rect 298228 409164 532700 409220
rect 532756 409164 532766 409220
rect 83944 409052 87276 409108
rect 87332 409052 87342 409108
rect 282258 409052 282268 409108
rect 282324 409052 534380 409108
rect 534436 409052 534446 409108
rect 295558 408940 295596 408996
rect 295652 408940 295662 408996
rect 268146 408604 268156 408660
rect 268212 408604 379596 408660
rect 379652 408604 379662 408660
rect 207890 408492 207900 408548
rect 207956 408492 356748 408548
rect 356804 408492 466956 408548
rect 467012 408492 467022 408548
rect 280242 408380 280252 408436
rect 280308 408380 430108 408436
rect 430164 408380 430174 408436
rect 307122 408268 307132 408324
rect 307188 408268 504700 408324
rect 504756 408268 504766 408324
rect 356514 408156 356524 408212
rect 356580 408156 367612 408212
rect 367668 408156 367678 408212
rect 379586 408156 379596 408212
rect 379652 408156 439740 408212
rect 439796 408156 439806 408212
rect 208002 408044 208012 408100
rect 208068 408044 259420 408100
rect 259476 408044 259486 408100
rect 300598 408044 300636 408100
rect 300692 408044 300702 408100
rect 337652 408044 352492 408100
rect 352548 408044 352558 408100
rect 355506 408044 355516 408100
rect 355572 408044 372764 408100
rect 372820 408044 372830 408100
rect 430098 408044 430108 408100
rect 430164 408044 486108 408100
rect 486164 408044 486174 408100
rect 186274 407932 186284 407988
rect 186340 407932 274652 407988
rect 274708 407932 274718 407988
rect 209458 407820 209468 407876
rect 209524 407820 268940 407876
rect 268996 407820 269006 407876
rect 208114 407708 208124 407764
rect 208180 407708 263788 407764
rect 263844 407708 263854 407764
rect 337652 407652 337708 408044
rect 348674 407932 348684 407988
rect 348740 407932 377916 407988
rect 377972 407932 377982 407988
rect 350578 407820 350588 407876
rect 350644 407820 398524 407876
rect 398580 407820 398590 407876
rect 399746 407820 399756 407876
rect 399812 407820 419132 407876
rect 419188 407820 419198 407876
rect 444854 407820 444892 407876
rect 444948 407820 444958 407876
rect 350354 407708 350364 407764
rect 350420 407708 408828 407764
rect 408884 407708 408894 407764
rect 419346 407708 419356 407764
rect 419412 407708 455196 407764
rect 455252 407708 455262 407764
rect 243954 407596 243964 407652
rect 244020 407596 337708 407652
rect 353714 407596 353724 407652
rect 353780 407596 393372 407652
rect 393428 407596 393438 407652
rect 397282 407596 397292 407652
rect 397348 407596 450044 407652
rect 450100 407596 450110 407652
rect 496374 407596 496412 407652
rect 496468 407596 496478 407652
rect 238802 407484 238812 407540
rect 238868 407484 352604 407540
rect 352660 407484 352670 407540
rect 355170 407484 355180 407540
rect 355236 407484 383068 407540
rect 383124 407484 383134 407540
rect 383282 407484 383292 407540
rect 383348 407484 429436 407540
rect 429492 407484 429502 407540
rect 445106 407484 445116 407540
rect 445172 407484 501564 407540
rect 501620 407484 501630 407540
rect 522134 407484 522172 407540
rect 522228 407484 522238 407540
rect 527286 407484 527324 407540
rect 527380 407484 527390 407540
rect 352604 407428 352660 407484
rect 87266 407372 87276 407428
rect 87332 407372 168028 407428
rect 168084 407372 168094 407428
rect 189298 407372 189308 407428
rect 189364 407372 210364 407428
rect 210420 407372 210430 407428
rect 233650 407372 233660 407428
rect 233716 407372 342916 407428
rect 352604 407372 356076 407428
rect 356132 407372 356142 407428
rect 356402 407372 356412 407428
rect 356468 407372 403676 407428
rect 403732 407372 403742 407428
rect 403890 407372 403900 407428
rect 403956 407372 424284 407428
rect 424340 407372 424350 407428
rect 424946 407372 424956 407428
rect 425012 407372 517020 407428
rect 517076 407372 517086 407428
rect 342860 407204 342916 407372
rect 345202 407260 345212 407316
rect 345268 407260 362460 407316
rect 362516 407260 362526 407316
rect 254258 407148 254268 407204
rect 254324 407148 342804 407204
rect 342860 407148 352716 407204
rect 352772 407148 357756 407204
rect 357812 407148 357822 407204
rect 342748 407092 342804 407148
rect 249106 407036 249116 407092
rect 249172 407036 337708 407092
rect 342738 407036 342748 407092
rect 342804 407036 342814 407092
rect 342972 407036 351148 407092
rect 351204 407036 351214 407092
rect 337652 406868 337708 407036
rect 342972 406868 343028 407036
rect 337652 406812 343028 406868
rect 206658 406700 206668 406756
rect 206724 406700 207900 406756
rect 207956 406700 207966 406756
rect 342738 406700 342748 406756
rect 342804 406700 351260 406756
rect 351316 406700 352268 406756
rect 352324 406700 352334 406756
rect 490578 406700 490588 406756
rect 490644 406700 490682 406756
rect 168018 406588 168028 406644
rect 168084 406588 218204 406644
rect 218260 406588 218270 406644
rect 228498 406588 228508 406644
rect 228564 406588 229964 406644
rect 230020 406588 230030 406644
rect 259410 406588 259420 406644
rect 259476 406588 260428 406644
rect 260484 406588 260494 406644
rect 280438 406588 280476 406644
rect 280532 406588 280542 406644
rect 295558 406588 295596 406644
rect 295652 406588 295662 406644
rect 351138 406588 351148 406644
rect 351204 406588 352044 406644
rect 352100 406588 352110 406644
rect 352482 406588 352492 406644
rect 352548 406588 354396 406644
rect 354452 406588 354462 406644
rect 464482 406588 464492 406644
rect 464548 406588 465500 406644
rect 465556 406588 465566 406644
rect 472882 406588 472892 406644
rect 472948 406588 581756 406644
rect 581812 406588 587132 406644
rect 587188 406588 587198 406644
rect 355394 406476 355404 406532
rect 355460 406476 413980 406532
rect 414036 406476 414046 406532
rect 252690 406364 252700 406420
rect 252756 406364 446012 406420
rect 446068 406364 446078 406420
rect 283602 406252 283612 406308
rect 283668 406252 534268 406308
rect 534324 406252 534334 406308
rect 83916 405412 83972 406168
rect 286290 406140 286300 406196
rect 286356 406140 537628 406196
rect 537684 406140 537694 406196
rect 196532 406028 213052 406084
rect 213108 406028 466172 406084
rect 466228 406028 466238 406084
rect 196532 405748 196588 406028
rect 259410 405916 259420 405972
rect 259476 405916 531020 405972
rect 531076 405916 531086 405972
rect 218194 405804 218204 405860
rect 218260 405804 252028 405860
rect 252084 405804 252094 405860
rect 261202 405804 261212 405860
rect 261268 405804 533036 405860
rect 533092 405804 533102 405860
rect 168018 405692 168028 405748
rect 168084 405692 196588 405748
rect 251346 405692 251356 405748
rect 251412 405692 531244 405748
rect 531300 405692 531310 405748
rect 83916 405356 90748 405412
rect 90692 404964 90748 405356
rect 90692 404908 92428 404964
rect 92484 404908 168028 404964
rect 168084 404908 168094 404964
rect 352594 404908 352604 404964
rect 352660 404908 357308 404964
rect 357364 404908 357374 404964
rect 257842 404796 257852 404852
rect 257908 404796 388220 404852
rect 388276 404796 388286 404852
rect 262770 404684 262780 404740
rect 262836 404684 399756 404740
rect 399812 404684 399822 404740
rect 266802 404572 266812 404628
rect 266868 404572 434588 404628
rect 434644 404572 434654 404628
rect 353602 404460 353612 404516
rect 353668 404460 532924 404516
rect 532980 404460 532990 404516
rect 350242 404348 350252 404404
rect 350308 404348 532812 404404
rect 532868 404348 532878 404404
rect 284722 404236 284732 404292
rect 284788 404236 480956 404292
rect 481012 404236 481022 404292
rect 308242 404124 308252 404180
rect 308308 404124 532588 404180
rect 532644 404124 532654 404180
rect 186386 404012 186396 404068
rect 186452 404012 211036 404068
rect 211092 404012 211102 404068
rect 252018 404012 252028 404068
rect 252084 404012 583884 404068
rect 583940 404012 584668 404068
rect -960 403732 480 403928
rect 584612 403844 584668 404012
rect 584612 403816 595672 403844
rect 584612 403788 597000 403816
rect -960 403704 59612 403732
rect 392 403676 59612 403704
rect 59668 403676 59678 403732
rect 595560 403592 597000 403788
rect 83944 403228 89964 403284
rect 90020 403228 90030 403284
rect 206994 403228 207004 403284
rect 207060 403228 583772 403284
rect 583828 403228 583838 403284
rect 355282 403004 355292 403060
rect 355348 403004 472892 403060
rect 472948 403004 472958 403060
rect 264114 402892 264124 402948
rect 264180 402892 403900 402948
rect 403956 402892 403966 402948
rect 280914 402780 280924 402836
rect 280980 402780 529340 402836
rect 529396 402780 529406 402836
rect 279570 402668 279580 402724
rect 279636 402668 535948 402724
rect 536004 402668 536014 402724
rect 278226 402556 278236 402612
rect 278292 402556 536060 402612
rect 536116 402556 536126 402612
rect 267474 402444 267484 402500
rect 267540 402444 529564 402500
rect 529620 402444 529630 402500
rect 208338 402332 208348 402388
rect 208404 402332 540092 402388
rect 540148 402332 540158 402388
rect 300402 401660 300412 401716
rect 300468 401660 421596 401716
rect 421652 401660 421662 401716
rect 355506 401548 355516 401604
rect 355572 401548 497644 401604
rect 497700 401548 497710 401604
rect 270162 401324 270172 401380
rect 270228 401324 529452 401380
rect 529508 401324 529518 401380
rect 274194 401212 274204 401268
rect 274260 401212 534492 401268
rect 534548 401212 534558 401268
rect 275538 401100 275548 401156
rect 275604 401100 536172 401156
rect 536228 401100 536238 401156
rect 271506 400988 271516 401044
rect 271572 400988 534604 401044
rect 534660 400988 534670 401044
rect 272850 400876 272860 400932
rect 272916 400876 536284 400932
rect 536340 400876 536350 400932
rect 268818 400764 268828 400820
rect 268884 400764 534716 400820
rect 534772 400764 534782 400820
rect 250002 400652 250012 400708
rect 250068 400652 531132 400708
rect 531188 400652 531198 400708
rect 83944 400316 89852 400372
rect 89908 400316 89918 400372
rect 350466 399980 350476 400036
rect 350532 399980 442092 400036
rect 442148 399980 442158 400036
rect 299730 399868 299740 399924
rect 299796 399868 414092 399924
rect 414148 399868 414158 399924
rect 265458 399756 265468 399812
rect 265524 399756 383292 399812
rect 383348 399756 383358 399812
rect 288306 399644 288316 399700
rect 288372 399644 424956 399700
rect 425012 399644 425022 399700
rect 353826 399532 353836 399588
rect 353892 399532 506716 399588
rect 506772 399532 506782 399588
rect 284274 399420 284284 399476
rect 284340 399420 445116 399476
rect 445172 399420 445182 399476
rect 264786 399308 264796 399364
rect 264852 399308 529676 399364
rect 529732 399308 529742 399364
rect 263442 399196 263452 399252
rect 263508 399196 529900 399252
rect 529956 399196 529966 399252
rect 208226 399084 208236 399140
rect 208292 399084 211708 399140
rect 211764 399084 211774 399140
rect 262098 399084 262108 399140
rect 262164 399084 530012 399140
rect 530068 399084 530078 399140
rect 160402 398972 160412 399028
rect 160468 398972 219100 399028
rect 219156 398972 219166 399028
rect 248658 398972 248668 399028
rect 248724 398972 530124 399028
rect 530180 398972 530190 399028
rect 303762 398188 303772 398244
rect 303828 398188 469196 398244
rect 469252 398188 469262 398244
rect 220052 398076 223356 398132
rect 223412 398076 355292 398132
rect 355348 398076 355358 398132
rect 165442 397852 165452 397908
rect 165508 397852 215068 397908
rect 215124 397852 215134 397908
rect 220052 397796 220108 398076
rect 172162 397740 172172 397796
rect 172228 397740 220108 397796
rect 310482 397740 310492 397796
rect 310548 397740 539308 397796
rect 539364 397740 539374 397796
rect 177202 397628 177212 397684
rect 177268 397628 329308 397684
rect 329364 397628 329374 397684
rect 85250 397516 85260 397572
rect 85316 397516 86772 397572
rect 88162 397516 88172 397572
rect 88228 397516 324604 397572
rect 324660 397516 324670 397572
rect 86716 397460 86772 397516
rect 83944 397404 86492 397460
rect 86548 397404 86558 397460
rect 86716 397404 323932 397460
rect 323988 397404 323998 397460
rect 354834 397404 354844 397460
rect 354900 397404 371980 397460
rect 372036 397404 372046 397460
rect 414082 397404 414092 397460
rect 414148 397404 427644 397460
rect 427700 397404 427710 397460
rect 86706 397292 86716 397348
rect 86772 397292 328636 397348
rect 328692 397292 328702 397348
rect 354946 397292 354956 397348
rect 355012 397292 386428 397348
rect 386484 397292 386494 397348
rect 421586 397292 421596 397348
rect 421652 397292 435148 397348
rect 435204 397292 435214 397348
rect 355394 397180 355404 397236
rect 355460 397180 393148 397236
rect 393204 397180 393214 397236
rect 355058 397068 355068 397124
rect 355124 397068 406812 397124
rect 406868 397068 406878 397124
rect 297042 396956 297052 397012
rect 297108 396956 400204 397012
rect 400260 396956 400270 397012
rect 299058 396844 299068 396900
rect 299124 396844 420700 396900
rect 420756 396844 420766 396900
rect 429202 396844 429212 396900
rect 429268 396844 448588 396900
rect 448644 396844 448654 396900
rect 546214 396844 546252 396900
rect 546308 396844 546318 396900
rect 573990 396844 574028 396900
rect 574084 396844 574094 396900
rect 361218 396732 361228 396788
rect 361284 396732 518028 396788
rect 518084 396732 518094 396788
rect 580934 396732 580972 396788
rect 581028 396732 581038 396788
rect 309810 396620 309820 396676
rect 309876 396620 531804 396676
rect 531860 396620 531870 396676
rect 553158 396620 553196 396676
rect 553252 396620 553262 396676
rect 403106 396508 403116 396564
rect 403172 396508 413756 396564
rect 413812 396508 413822 396564
rect 451836 396508 455308 396564
rect 455364 396508 455374 396564
rect 567046 396508 567084 396564
rect 567140 396508 567150 396564
rect 270722 396284 270732 396340
rect 270788 396284 397292 396340
rect 397348 396284 397358 396340
rect 272290 396172 272300 396228
rect 272356 396172 419356 396228
rect 419412 396172 419422 396228
rect 451836 396116 451892 396508
rect 302530 396060 302540 396116
rect 302596 396060 451892 396116
rect 273410 395948 273420 396004
rect 273476 395948 460348 396004
rect 460404 395948 460414 396004
rect 203186 395836 203196 395892
rect 203252 395836 213612 395892
rect 213668 395836 213678 395892
rect 274754 395836 274764 395892
rect 274820 395836 464492 395892
rect 464548 395836 464558 395892
rect 466162 395836 466172 395892
rect 466228 395836 582988 395892
rect 583044 395836 583054 395892
rect 175522 395724 175532 395780
rect 175588 395724 197596 395780
rect 197652 395724 197662 395780
rect 201506 395724 201516 395780
rect 201572 395724 214284 395780
rect 214340 395724 214350 395780
rect 276098 395724 276108 395780
rect 276164 395724 470652 395780
rect 470708 395724 470718 395780
rect 153682 395612 153692 395668
rect 153748 395612 215628 395668
rect 215684 395612 215694 395668
rect 277442 395612 277452 395668
rect 277508 395612 475804 395668
rect 475860 395612 475870 395668
rect 354946 395164 354956 395220
rect 355012 395164 355292 395220
rect 355348 395164 355358 395220
rect 361218 395164 361228 395220
rect 361284 395164 361322 395220
rect 356626 395052 356636 395108
rect 356692 395052 358204 395108
rect 358260 395052 358270 395108
rect 365110 395052 365148 395108
rect 365204 395052 365214 395108
rect 379782 395052 379820 395108
rect 379876 395052 379886 395108
rect 304994 394940 305004 394996
rect 305060 394940 483868 394996
rect 483924 394940 483934 394996
rect 525494 394940 525532 394996
rect 525588 394940 525598 394996
rect 305890 394828 305900 394884
rect 305956 394828 490812 394884
rect 490868 394828 490878 394884
rect 582978 394828 582988 394884
rect 583044 394828 583660 394884
rect 583716 394828 590604 394884
rect 590660 394828 590670 394884
rect 298274 394716 298284 394772
rect 298340 394716 403116 394772
rect 403172 394716 403182 394772
rect 476886 394716 476924 394772
rect 476980 394716 476990 394772
rect 511606 394716 511644 394772
rect 511700 394716 511710 394772
rect 301634 394604 301644 394660
rect 301700 394604 429212 394660
rect 429268 394604 429278 394660
rect 462998 394604 463036 394660
rect 463092 394604 463102 394660
rect 463698 394604 463708 394660
rect 463764 394604 590716 394660
rect 590772 394604 590782 394660
rect 83944 394492 211596 394548
rect 211652 394492 211662 394548
rect 276770 394492 276780 394548
rect 276836 394492 530908 394548
rect 530964 394492 530974 394548
rect 502292 394380 511644 394436
rect 511700 394380 511710 394436
rect 502292 394324 502348 394380
rect 307682 394268 307692 394324
rect 307748 394268 502348 394324
rect 354722 394156 354732 394212
rect 354788 394156 355068 394212
rect 355124 394156 355134 394212
rect 455252 394156 476924 394212
rect 476980 394156 476990 394212
rect 455252 394100 455308 394156
rect 304322 394044 304332 394100
rect 304388 394044 455308 394100
rect 463026 394044 463036 394100
rect 463092 394044 463102 394100
rect 463036 393988 463092 394044
rect 354050 393932 354060 393988
rect 354116 393932 463092 393988
rect 308354 393820 308364 393876
rect 308420 393820 361228 393876
rect 361284 393820 361294 393876
rect 365138 393820 365148 393876
rect 365204 393820 365214 393876
rect 365148 393764 365204 393820
rect 355170 393708 355180 393764
rect 355236 393708 365204 393764
rect 364466 393260 364476 393316
rect 364532 393260 393148 393316
rect 393204 393260 393214 393316
rect 343522 393148 343532 393204
rect 343588 393148 584668 393204
rect 584724 393148 584734 393204
rect 393138 393036 393148 393092
rect 393204 393036 463708 393092
rect 463764 393036 463774 393092
rect 173954 392812 173964 392868
rect 174020 392812 192444 392868
rect 192500 392812 192510 392868
rect 206322 392812 206332 392868
rect 206388 392812 212268 392868
rect 212324 392812 212334 392868
rect 294914 392812 294924 392868
rect 294980 392812 379820 392868
rect 379876 392812 379886 392868
rect 466946 392812 466956 392868
rect 467012 392812 590492 392868
rect 590548 392812 590558 392868
rect 177314 392700 177324 392756
rect 177380 392700 202748 392756
rect 202804 392700 202814 392756
rect 204642 392700 204652 392756
rect 204708 392700 212940 392756
rect 212996 392700 213006 392756
rect 155362 392588 155372 392644
rect 155428 392588 216300 392644
rect 216356 392588 216366 392644
rect 293570 392588 293580 392644
rect 293636 392588 355180 392644
rect 355236 392588 355246 392644
rect 189410 392476 189420 392532
rect 189476 392476 342860 392532
rect 342916 392476 342926 392532
rect 91522 392364 91532 392420
rect 91588 392364 325164 392420
rect 325220 392364 325230 392420
rect 86482 392252 86492 392308
rect 86548 392252 327180 392308
rect 327236 392252 327246 392308
rect 83944 391580 85708 391636
rect 85764 391580 85774 391636
rect 311042 391356 311052 391412
rect 311108 391356 355180 391412
rect 355236 391356 355246 391412
rect 309250 391244 309260 391300
rect 309316 391244 355292 391300
rect 355348 391244 355358 391300
rect 295810 391132 295820 391188
rect 295876 391132 354956 391188
rect 355012 391132 355022 391188
rect 211586 391020 211596 391076
rect 211652 391020 321804 391076
rect 321860 391020 321870 391076
rect 57922 390908 57932 390964
rect 57988 390908 216972 390964
rect 217028 390908 217038 390964
rect 294242 390908 294252 390964
rect 294308 390908 354844 390964
rect 354900 390908 354910 390964
rect 59602 390796 59612 390852
rect 59668 390796 219660 390852
rect 219716 390796 219726 390852
rect 286850 390796 286860 390852
rect 286916 390796 355404 390852
rect 355460 390796 355470 390852
rect 56242 390684 56252 390740
rect 56308 390684 217644 390740
rect 217700 390684 217710 390740
rect 253250 390684 253260 390740
rect 253316 390684 355068 390740
rect 355124 390684 355134 390740
rect 14242 390572 14252 390628
rect 14308 390572 218540 390628
rect 218596 390572 218606 390628
rect 250562 390572 250572 390628
rect 250628 390572 355516 390628
rect 355572 390572 355582 390628
rect 591154 390572 591164 390628
rect 591220 390600 595672 390628
rect 591220 390572 597000 390600
rect 313730 390460 313740 390516
rect 313796 390460 355068 390516
rect 355124 390460 355134 390516
rect 595560 390376 597000 390572
rect -960 389620 480 389816
rect 320898 389788 320908 389844
rect 320964 389788 321244 389844
rect 321300 389788 351820 389844
rect 351876 389788 351886 389844
rect -960 389592 4284 389620
rect 392 389564 4284 389592
rect 4340 389564 4350 389620
rect 337652 389452 355628 389508
rect 355684 389452 355694 389508
rect 337652 389172 337708 389452
rect 205090 389116 205100 389172
rect 205156 389116 337708 389172
rect 186050 389004 186060 389060
rect 186116 389004 343196 389060
rect 343252 389004 343262 389060
rect 4498 388892 4508 388948
rect 4564 388892 320908 388948
rect 320964 388892 320974 388948
rect 352594 388780 352604 388836
rect 352660 388780 355096 388836
rect 78418 388108 78428 388164
rect 78484 388108 318444 388164
rect 318500 388108 318510 388164
rect 298050 387884 298060 387940
rect 298116 387884 354732 387940
rect 354788 387884 354798 387940
rect 296818 387772 296828 387828
rect 296884 387772 355404 387828
rect 355460 387772 355470 387828
rect 291554 387660 291564 387716
rect 291620 387660 353612 387716
rect 353668 387660 353678 387716
rect 290210 387548 290220 387604
rect 290276 387548 353836 387604
rect 353892 387548 353902 387604
rect 260306 387436 260316 387492
rect 260372 387436 350364 387492
rect 350420 387436 350430 387492
rect 257954 387324 257964 387380
rect 258020 387324 350588 387380
rect 350644 387324 350654 387380
rect 186162 387212 186172 387268
rect 186228 387212 343308 387268
rect 343364 387212 343374 387268
rect 103282 386876 103292 386932
rect 103348 386876 240828 386932
rect 240884 386876 240894 386932
rect 96562 386764 96572 386820
rect 96628 386764 242844 386820
rect 242900 386764 242910 386820
rect 94882 386652 94892 386708
rect 94948 386652 242172 386708
rect 242228 386652 242238 386708
rect 95106 386540 95116 386596
rect 95172 386540 247100 386596
rect 247156 386540 247166 386596
rect 40898 386428 40908 386484
rect 40964 386428 232764 386484
rect 232820 386428 232830 386484
rect 69682 386092 69692 386148
rect 69748 386092 316092 386148
rect 316148 386092 316158 386148
rect 235106 385980 235116 386036
rect 235172 385980 268940 386036
rect 268996 385980 269006 386036
rect 283378 385980 283388 386036
rect 283444 385980 354956 386036
rect 355012 385980 355022 386036
rect 252466 385868 252476 385924
rect 252532 385868 348684 385924
rect 348740 385868 348750 385924
rect 248546 385756 248556 385812
rect 248612 385756 345212 385812
rect 345268 385756 345278 385812
rect 256610 385644 256620 385700
rect 256676 385644 353724 385700
rect 353780 385644 353790 385700
rect 185602 385532 185612 385588
rect 185668 385532 322700 385588
rect 322756 385532 322766 385588
rect 95330 385420 95340 385476
rect 95396 385420 246204 385476
rect 246260 385420 246270 385476
rect 104962 385308 104972 385364
rect 105028 385308 242060 385364
rect 242116 385308 242126 385364
rect 100146 385196 100156 385252
rect 100212 385196 237468 385252
rect 237524 385196 237534 385252
rect 96786 385084 96796 385140
rect 96852 385084 238812 385140
rect 238868 385084 238878 385140
rect 99922 384972 99932 385028
rect 99988 384972 245420 385028
rect 245476 384972 245486 385028
rect 274642 384972 274652 385028
rect 274708 384972 352044 385028
rect 352100 384972 352110 385028
rect 238354 384860 238364 384916
rect 238420 384860 325836 384916
rect 325892 384860 325902 384916
rect 315858 384748 315868 384804
rect 315924 384748 352380 384804
rect 352436 384748 352446 384804
rect 241826 384524 241836 384580
rect 241892 384524 289772 384580
rect 289828 384524 350364 384580
rect 350420 384524 350430 384580
rect 238466 384412 238476 384468
rect 238532 384412 283948 384468
rect 284004 384412 345548 384468
rect 345604 384412 345614 384468
rect 238578 384300 238588 384356
rect 238644 384300 315868 384356
rect 315924 384300 315934 384356
rect 269938 384188 269948 384244
rect 270004 384188 348572 384244
rect 348628 384188 348638 384244
rect 180562 384076 180572 384132
rect 180628 384076 325948 384132
rect 326004 384076 326014 384132
rect 85026 383964 85036 384020
rect 85092 383964 326284 384020
rect 326340 383964 326350 384020
rect 84802 383852 84812 383908
rect 84868 383852 327628 383908
rect 327684 383852 327694 383908
rect 336690 383852 336700 383908
rect 336756 383852 345772 383908
rect 345828 383852 345838 383908
rect 185714 383516 185724 383572
rect 185780 383516 316652 383572
rect 316708 383516 316718 383572
rect 95554 383404 95564 383460
rect 95620 383404 239372 383460
rect 239428 383404 239438 383460
rect 38434 383292 38444 383348
rect 38500 383292 228732 383348
rect 228788 383292 228798 383348
rect 38546 383180 38556 383236
rect 38612 383180 229292 383236
rect 229348 383180 229358 383236
rect 24322 383068 24332 383124
rect 24388 383068 223468 383124
rect 223524 383068 223534 383124
rect 237794 383068 237804 383124
rect 237860 383068 339388 383124
rect 339444 383068 339454 383124
rect 341842 383068 341852 383124
rect 341908 383068 350588 383124
rect 350644 383068 350654 383124
rect 255042 382956 255052 383012
rect 255108 382956 257852 383012
rect 257908 382956 257918 383012
rect 320002 382956 320012 383012
rect 320068 382956 355516 383012
rect 355572 382956 355582 383012
rect 285506 382844 285516 382900
rect 285572 382844 308252 382900
rect 308308 382844 308318 382900
rect 313058 382844 313068 382900
rect 313124 382844 348572 382900
rect 348628 382844 348638 382900
rect 256946 382732 256956 382788
rect 257012 382732 288092 382788
rect 288148 382732 288158 382788
rect 289538 382732 289548 382788
rect 289604 382732 291452 382788
rect 291508 382732 291518 382788
rect 301522 382732 301532 382788
rect 301588 382732 350476 382788
rect 350532 382732 350542 382788
rect 352146 382732 352156 382788
rect 352212 382732 355096 382788
rect 111682 382620 111692 382676
rect 111748 382620 240268 382676
rect 240324 382620 240334 382676
rect 261314 382620 261324 382676
rect 261380 382620 298172 382676
rect 298228 382620 298238 382676
rect 303538 382620 303548 382676
rect 303604 382620 354060 382676
rect 354116 382620 354126 382676
rect 202738 382508 202748 382564
rect 202804 382508 203196 382564
rect 203252 382508 203262 382564
rect 204194 382508 204204 382564
rect 204260 382508 204764 382564
rect 204820 382508 204830 382564
rect 206098 382508 206108 382564
rect 206164 382508 206556 382564
rect 206612 382508 206622 382564
rect 209458 382508 209468 382564
rect 209524 382508 209916 382564
rect 209972 382508 209982 382564
rect 286066 382508 286076 382564
rect 286132 382508 353836 382564
rect 353892 382508 353902 382564
rect 201366 382396 201404 382452
rect 201460 382396 201470 382452
rect 203046 382396 203084 382452
rect 203140 382396 203150 382452
rect 204838 382396 204876 382452
rect 204932 382396 204942 382452
rect 206406 382396 206444 382452
rect 206500 382396 206510 382452
rect 208086 382396 208124 382452
rect 208180 382396 208190 382452
rect 209766 382396 209804 382452
rect 209860 382396 209870 382452
rect 258626 382396 258636 382452
rect 258692 382396 350252 382452
rect 350308 382396 350318 382452
rect 185602 382284 185612 382340
rect 185668 382284 235228 382340
rect 235284 382284 235294 382340
rect 254706 382284 254716 382340
rect 254772 382284 261212 382340
rect 261268 382284 261278 382340
rect 261986 382284 261996 382340
rect 262052 382284 355292 382340
rect 355348 382284 355358 382340
rect 170594 382172 170604 382228
rect 170660 382172 233548 382228
rect 233604 382172 233614 382228
rect 256050 382172 256060 382228
rect 256116 382172 353612 382228
rect 353668 382172 353678 382228
rect 167122 382060 167132 382116
rect 167188 382060 226492 382116
rect 226548 382060 226558 382116
rect 226678 382060 226716 382116
rect 226772 382060 226782 382116
rect 279346 382060 279356 382116
rect 279412 382060 284732 382116
rect 284788 382060 284798 382116
rect 292226 382060 292236 382116
rect 292292 382060 301532 382116
rect 301588 382060 301598 382116
rect 306898 382060 306908 382116
rect 306964 382060 320012 382116
rect 320068 382060 320078 382116
rect 168802 381948 168812 382004
rect 168868 381948 245532 382004
rect 245588 381948 245598 382004
rect 249778 381948 249788 382004
rect 249844 381948 250236 382004
rect 250292 381948 250302 382004
rect 259186 381948 259196 382004
rect 259252 381948 260316 382004
rect 260372 381948 260382 382004
rect 266578 381948 266588 382004
rect 266644 381948 267036 382004
rect 267092 381948 267102 382004
rect 281670 381948 281708 382004
rect 281764 381948 281774 382004
rect 288082 381948 288092 382004
rect 288148 381948 288876 382004
rect 288932 381948 288942 382004
rect 290518 381948 290556 382004
rect 290612 381948 290622 382004
rect 293458 381948 293468 382004
rect 293524 381948 293916 382004
rect 293972 381948 293982 382004
rect 312358 381948 312396 382004
rect 312452 381948 312462 382004
rect 313618 381948 313628 382004
rect 313684 381948 314076 382004
rect 314132 381948 314142 382004
rect 315074 381948 315084 382004
rect 315140 381948 315756 382004
rect 315812 381948 315822 382004
rect 322578 381948 322588 382004
rect 322644 381948 322924 382004
rect 322980 381948 322990 382004
rect 118402 381836 118412 381892
rect 118468 381836 238588 381892
rect 238644 381836 238654 381892
rect 113362 381724 113372 381780
rect 113428 381724 233996 381780
rect 234052 381724 234062 381780
rect 120082 381612 120092 381668
rect 120148 381612 244076 381668
rect 244132 381612 244142 381668
rect 116722 381500 116732 381556
rect 116788 381500 243740 381556
rect 243796 381500 243806 381556
rect 226482 381388 226492 381444
rect 226548 381388 230636 381444
rect 230692 381388 230702 381444
rect 232754 381388 232764 381444
rect 232820 381388 236124 381444
rect 236180 381388 236190 381444
rect 241490 381388 241500 381444
rect 241556 381388 331604 381444
rect 350802 381388 350812 381444
rect 350868 381388 352156 381444
rect 352212 381388 352222 381444
rect 331548 381332 331604 381388
rect 331538 381276 331548 381332
rect 331604 381276 345436 381332
rect 345492 381276 345502 381332
rect 55570 380940 55580 380996
rect 55636 380940 315196 380996
rect 315252 380940 315262 380996
rect 240146 380828 240156 380884
rect 240212 380828 260428 380884
rect 260484 380828 260494 380884
rect 237682 380716 237692 380772
rect 237748 380716 263788 380772
rect 263844 380716 263854 380772
rect 311602 380716 311612 380772
rect 311668 380716 350924 380772
rect 350980 380716 350990 380772
rect 170482 380604 170492 380660
rect 170548 380604 236908 380660
rect 236964 380604 236974 380660
rect 241714 380604 241724 380660
rect 241780 380604 274652 380660
rect 274708 380604 274718 380660
rect 306562 380604 306572 380660
rect 306628 380604 346892 380660
rect 346948 380604 346958 380660
rect 185938 380492 185948 380548
rect 186004 380492 315868 380548
rect 315924 380492 315934 380548
rect 325826 380492 325836 380548
rect 325892 380492 352156 380548
rect 352212 380492 352222 380548
rect 38322 380380 38332 380436
rect 38388 380380 231868 380436
rect 231924 380380 231934 380436
rect 121762 380268 121772 380324
rect 121828 380268 319340 380324
rect 319396 380268 319406 380324
rect 14242 380156 14252 380212
rect 14308 380156 222572 380212
rect 222628 380156 222638 380212
rect 292898 380156 292908 380212
rect 292964 380156 340172 380212
rect 340228 380156 340238 380212
rect 93650 380044 93660 380100
rect 93716 380044 320908 380100
rect 320964 380044 320974 380100
rect 91522 379932 91532 379988
rect 91588 379932 320572 379988
rect 320628 379932 320638 379988
rect 82226 379820 82236 379876
rect 82292 379820 319228 379876
rect 319284 379820 319294 379876
rect 200834 379708 200844 379764
rect 200900 379708 201292 379764
rect 201348 379708 201358 379764
rect 202178 379708 202188 379764
rect 202244 379708 202860 379764
rect 202916 379708 202926 379764
rect 315746 379708 315756 379764
rect 315812 379708 343420 379764
rect 343476 379708 343486 379764
rect 34402 379596 34412 379652
rect 34468 379596 214172 379652
rect 214228 379596 214238 379652
rect 214386 379596 214396 379652
rect 214452 379596 220444 379652
rect 220500 379596 220510 379652
rect 221788 379596 230580 379652
rect 221788 379540 221844 379596
rect 230524 379540 230580 379596
rect 38210 379484 38220 379540
rect 38276 379484 221844 379540
rect 221974 379484 222012 379540
rect 222068 379484 222078 379540
rect 223990 379484 224028 379540
rect 224084 379484 224094 379540
rect 227574 379484 227612 379540
rect 227668 379484 227678 379540
rect 229058 379484 229068 379540
rect 229124 379484 230076 379540
rect 230132 379484 230142 379540
rect 230514 379484 230524 379540
rect 230580 379484 230590 379540
rect 235414 379484 235452 379540
rect 235508 379484 235518 379540
rect 74610 379372 74620 379428
rect 74676 379372 317884 379428
rect 317940 379372 317950 379428
rect 196532 379260 221116 379316
rect 221172 379260 221182 379316
rect 221778 379260 221788 379316
rect 221844 379260 221854 379316
rect 225110 379260 225148 379316
rect 225204 379260 225214 379316
rect 225782 379260 225820 379316
rect 225876 379260 225886 379316
rect 227798 379260 227836 379316
rect 227892 379260 227902 379316
rect 232502 379260 232540 379316
rect 232596 379260 232606 379316
rect 196532 379092 196588 379260
rect 221788 379204 221844 379260
rect 214162 379148 214172 379204
rect 214228 379148 221844 379204
rect 49522 379036 49532 379092
rect 49588 379036 196588 379092
rect 214386 379036 214396 379092
rect 214452 379036 214462 379092
rect 214396 378980 214452 379036
rect 120194 378924 120204 378980
rect 120260 378924 214452 378980
rect 346994 377468 347004 377524
rect 347060 377468 352492 377524
rect 352548 377468 355124 377524
rect 355068 376712 355124 377468
rect 595560 377188 597000 377384
rect 583762 377132 583772 377188
rect 583828 377160 597000 377188
rect 583828 377132 595672 377160
rect 392 375704 4172 375732
rect -960 375676 4172 375704
rect 4228 375676 4238 375732
rect -960 375480 480 375676
rect 339864 373996 343196 374052
rect 343252 373996 343262 374052
rect 339864 373100 344092 373156
rect 344148 373100 344158 373156
rect 339864 372204 343532 372260
rect 343588 372204 343598 372260
rect 339864 371308 344204 371364
rect 344260 371308 344270 371364
rect 350578 370636 350588 370692
rect 350644 370636 351932 370692
rect 351988 370636 355096 370692
rect 339864 370412 348572 370468
rect 348628 370412 348638 370468
rect 339864 369516 340620 369572
rect 340676 369516 340686 369572
rect 190652 368116 190708 368648
rect 339864 368620 346892 368676
rect 346948 368620 346958 368676
rect 190642 368060 190652 368116
rect 190708 368060 190718 368116
rect 339864 367724 355292 367780
rect 355348 367724 355358 367780
rect 190652 366996 190708 367528
rect 190642 366940 190652 366996
rect 190708 366940 190718 366996
rect 339864 366828 353612 366884
rect 353668 366828 353678 366884
rect 190642 366380 190652 366436
rect 190708 366380 190718 366436
rect 345762 366156 345772 366212
rect 345828 366156 352268 366212
rect 352324 366156 352334 366212
rect 339864 365932 345324 365988
rect 345380 365932 345390 365988
rect 190652 364644 190708 365288
rect 339864 365036 343084 365092
rect 343140 365036 343150 365092
rect 190642 364588 190652 364644
rect 190708 364588 190718 364644
rect 352258 364588 352268 364644
rect 352324 364588 355096 364644
rect 86034 363916 86044 363972
rect 86100 363916 121772 363972
rect 121828 363916 121838 363972
rect 70802 363804 70812 363860
rect 70868 363804 185724 363860
rect 185780 363804 185790 363860
rect 63186 363692 63196 363748
rect 63252 363692 185948 363748
rect 186004 363692 186014 363748
rect 190092 363300 190148 364168
rect 339864 364140 350252 364196
rect 350308 364140 350318 364196
rect 590594 364140 590604 364196
rect 590660 364168 595672 364196
rect 590660 364140 597000 364168
rect 595560 363944 597000 364140
rect 165900 363244 190148 363300
rect 339490 363244 339500 363300
rect 339556 363244 339566 363300
rect 59378 363020 59388 363076
rect 59444 363020 85708 363076
rect 85764 363020 85774 363076
rect 165900 363048 165956 363244
rect 186498 363020 186508 363076
rect 186564 363020 190120 363076
rect 66994 362908 67004 362964
rect 67060 362908 69692 362964
rect 69748 362908 69758 362964
rect 89842 362908 89852 362964
rect 89908 362908 91532 362964
rect 91588 362908 91598 362964
rect 339864 362348 348684 362404
rect 348740 362348 348750 362404
rect 186610 361900 186620 361956
rect 186676 361900 190120 361956
rect -960 361396 480 361592
rect 339864 361452 355404 361508
rect 355460 361452 355470 361508
rect -960 361368 120204 361396
rect 392 361340 120204 361368
rect 120260 361340 120270 361396
rect 85698 361228 85708 361284
rect 85764 361228 91532 361284
rect 91588 361228 91598 361284
rect 179778 360780 179788 360836
rect 179844 360780 190120 360836
rect 339864 360556 353612 360612
rect 353668 360556 353678 360612
rect 173012 359772 186508 359828
rect 186564 359772 186574 359828
rect 173012 359716 173068 359772
rect 165928 359660 173068 359716
rect 186386 359660 186396 359716
rect 186452 359660 190120 359716
rect 339864 359660 347004 359716
rect 347060 359660 347070 359716
rect 339864 358764 350476 358820
rect 350532 358764 350542 358820
rect 89954 358652 89964 358708
rect 90020 358652 93324 358708
rect 93380 358652 93390 358708
rect 168914 358540 168924 358596
rect 168980 358540 190120 358596
rect 345426 358540 345436 358596
rect 345492 358540 355096 358596
rect 339864 357868 345212 357924
rect 345268 357868 345278 357924
rect 177202 357420 177212 357476
rect 177268 357420 190120 357476
rect 167020 356412 186620 356468
rect 186676 356412 186686 356468
rect 167020 356356 167076 356412
rect 339612 356356 339668 357000
rect 165928 356300 167076 356356
rect 167234 356300 167244 356356
rect 167300 356300 190120 356356
rect 339602 356300 339612 356356
rect 339668 356300 339678 356356
rect 339864 356076 341852 356132
rect 341908 356076 341918 356132
rect 176194 355180 176204 355236
rect 176260 355180 190120 355236
rect 339864 355180 350588 355236
rect 350644 355180 350654 355236
rect 339864 354284 348796 354340
rect 348852 354284 348862 354340
rect 184594 354060 184604 354116
rect 184660 354060 190120 354116
rect 339864 353388 353724 353444
rect 353780 353388 353790 353444
rect 165928 352940 179788 352996
rect 179844 352940 179854 352996
rect 181346 352940 181356 352996
rect 181412 352940 190120 352996
rect 339864 352492 341964 352548
rect 342020 352492 342030 352548
rect 352146 352492 352156 352548
rect 352212 352492 355096 352548
rect 177874 351820 177884 351876
rect 177940 351820 190120 351876
rect 339864 351596 355292 351652
rect 355348 351596 355358 351652
rect 591042 350924 591052 350980
rect 591108 350952 595672 350980
rect 591108 350924 597000 350952
rect 189298 350700 189308 350756
rect 189364 350700 190120 350756
rect 595560 350728 597000 350924
rect 339724 350196 339780 350728
rect 339714 350140 339724 350196
rect 339780 350140 339790 350196
rect 339864 349804 353836 349860
rect 353892 349804 353902 349860
rect 165928 349580 186396 349636
rect 186452 349580 186462 349636
rect 187404 349580 190120 349636
rect 187404 349524 187460 349580
rect 176306 349468 176316 349524
rect 176372 349468 187460 349524
rect 339864 348908 345436 348964
rect 345492 348908 345502 348964
rect 179442 348460 179452 348516
rect 179508 348460 190120 348516
rect 339864 348012 350700 348068
rect 350756 348012 350766 348068
rect -960 347284 480 347480
rect 176082 347340 176092 347396
rect 176148 347340 190120 347396
rect -960 347256 4396 347284
rect 392 347228 4396 347256
rect 4452 347228 4462 347284
rect 339266 347116 339276 347172
rect 339332 347116 339342 347172
rect 351810 346444 351820 346500
rect 351876 346444 352716 346500
rect 352772 346444 355096 346500
rect 165928 346220 168140 346276
rect 168196 346220 168206 346276
rect 177986 346220 177996 346276
rect 178052 346220 190120 346276
rect 339864 346220 349020 346276
rect 349076 346220 349086 346276
rect 339864 345324 348908 345380
rect 348964 345324 348974 345380
rect 177762 345100 177772 345156
rect 177828 345100 190120 345156
rect 339864 344428 342860 344484
rect 342916 344428 342926 344484
rect 339378 344204 339388 344260
rect 339444 344204 339454 344260
rect 179666 343980 179676 344036
rect 179732 343980 190120 344036
rect 339388 343560 339444 344204
rect 165928 342860 168028 342916
rect 168084 342860 168094 342916
rect 181122 342860 181132 342916
rect 181188 342860 190120 342916
rect 339864 342636 343980 342692
rect 344036 342636 344046 342692
rect 182690 341740 182700 341796
rect 182756 341740 190120 341796
rect 339864 341740 343868 341796
rect 343924 341740 343934 341796
rect 339864 340844 342972 340900
rect 343028 340844 343038 340900
rect 179330 340620 179340 340676
rect 179396 340620 190120 340676
rect 351922 340396 351932 340452
rect 351988 340396 352380 340452
rect 352436 340396 355096 340452
rect 339864 339948 343644 340004
rect 343700 339948 343710 340004
rect 165928 339500 168028 339556
rect 168084 339500 168094 339556
rect 179554 339500 179564 339556
rect 179620 339500 190120 339556
rect 339864 339052 343532 339108
rect 343588 339052 343598 339108
rect 181234 338380 181244 338436
rect 181300 338380 190120 338436
rect 339864 338156 354508 338212
rect 354564 338156 354574 338212
rect 595560 337652 597000 337736
rect 590818 337596 590828 337652
rect 590884 337596 597000 337652
rect 595560 337512 597000 337596
rect 184482 337260 184492 337316
rect 184548 337260 190120 337316
rect 339864 337260 341068 337316
rect 341124 337260 341134 337316
rect 165900 336812 168140 336868
rect 168196 336812 177324 336868
rect 177380 336812 177390 336868
rect 165900 336168 165956 336812
rect 182914 336140 182924 336196
rect 182980 336140 190120 336196
rect 339836 336084 339892 336392
rect 339826 336028 339836 336084
rect 339892 336028 339902 336084
rect 339864 335468 346780 335524
rect 346836 335468 346846 335524
rect 181010 335020 181020 335076
rect 181076 335020 190120 335076
rect 339864 334572 346556 334628
rect 346612 334572 346622 334628
rect 350018 334348 350028 334404
rect 350084 334348 350924 334404
rect 350980 334348 355096 334404
rect 189186 333900 189196 333956
rect 189252 333900 190120 333956
rect 339864 333676 348684 333732
rect 348740 333676 348750 333732
rect 392 333368 4508 333396
rect -960 333340 4508 333368
rect 4564 333340 4574 333396
rect -960 333144 480 333340
rect 165928 332780 168252 332836
rect 168308 332780 175532 332836
rect 175588 332780 175598 332836
rect 186386 332780 186396 332836
rect 186452 332780 190120 332836
rect 339864 332780 346108 332836
rect 346164 332780 346174 332836
rect 339864 331884 346668 331940
rect 346724 331884 346734 331940
rect 172946 331660 172956 331716
rect 173012 331660 190120 331716
rect 339864 330988 345548 331044
rect 345604 330988 345614 331044
rect 168690 330876 168700 330932
rect 168756 330876 173964 330932
rect 174020 330876 174030 330932
rect 174402 330540 174412 330596
rect 174468 330540 190120 330596
rect 339836 329476 339892 330120
rect 165928 329420 168364 329476
rect 168420 329420 168700 329476
rect 168756 329420 168766 329476
rect 182802 329420 182812 329476
rect 182868 329420 190120 329476
rect 339836 329420 340116 329476
rect 340060 329364 340116 329420
rect 340050 329308 340060 329364
rect 340116 329308 340126 329364
rect 339864 329196 353724 329252
rect 353780 329196 353790 329252
rect 175970 328300 175980 328356
rect 176036 328300 190120 328356
rect 339864 328300 344988 328356
rect 345044 328300 345054 328356
rect 346770 328300 346780 328356
rect 346836 328300 355068 328356
rect 355124 328300 355134 328356
rect 339864 327404 348908 327460
rect 348964 327404 348974 327460
rect 179218 327180 179228 327236
rect 179284 327180 190120 327236
rect 339864 326508 342076 326564
rect 342132 326508 342142 326564
rect 165928 326060 168924 326116
rect 168980 326060 168990 326116
rect 174626 326060 174636 326116
rect 174692 326060 190120 326116
rect 339864 325612 341964 325668
rect 342020 325612 342030 325668
rect 174514 324940 174524 324996
rect 174580 324940 190120 324996
rect 339864 324716 345324 324772
rect 345380 324716 345390 324772
rect 590482 324492 590492 324548
rect 590548 324520 595672 324548
rect 590548 324492 597000 324520
rect 595560 324296 597000 324492
rect 182578 323820 182588 323876
rect 182644 323820 190120 323876
rect 339864 323820 350588 323876
rect 350644 323820 350654 323876
rect 339864 322924 350364 322980
rect 350420 322924 350430 322980
rect 165928 322728 172172 322756
rect 165900 322700 172172 322728
rect 172228 322700 172238 322756
rect 186274 322700 186284 322756
rect 186340 322700 190120 322756
rect 165900 322084 165956 322700
rect 354386 322252 354396 322308
rect 354452 322252 355096 322308
rect 165890 322028 165900 322084
rect 165956 322028 165966 322084
rect 339864 322028 349020 322084
rect 349076 322028 349086 322084
rect 152786 321804 152796 321860
rect 152852 321804 167244 321860
rect 167300 321804 167310 321860
rect 108322 321692 108332 321748
rect 108388 321692 165900 321748
rect 165956 321692 165966 321748
rect 189074 321580 189084 321636
rect 189140 321580 190120 321636
rect 339864 321132 341068 321188
rect 341124 321132 341134 321188
rect 342402 320908 342412 320964
rect 342468 320908 354396 320964
rect 354452 320908 354462 320964
rect 184482 320460 184492 320516
rect 184548 320460 190120 320516
rect 339864 320236 344092 320292
rect 344148 320236 344158 320292
rect 106642 320012 106652 320068
rect 106708 320012 168140 320068
rect 168196 320012 168206 320068
rect 190642 319340 190652 319396
rect 190708 319340 190718 319396
rect 339864 319340 341180 319396
rect 341236 319340 341246 319396
rect -960 319060 480 319256
rect -960 319032 49532 319060
rect 392 319004 49532 319032
rect 49588 319004 49598 319060
rect 339864 318444 349132 318500
rect 349188 318444 349198 318500
rect 167234 318220 167244 318276
rect 167300 318220 190120 318276
rect 339864 317548 344876 317604
rect 344932 317548 344942 317604
rect 182802 317100 182812 317156
rect 182868 317100 190120 317156
rect 339378 316988 339388 317044
rect 339444 316988 354060 317044
rect 354116 316988 355124 317044
rect 339864 316652 344652 316708
rect 344708 316652 344718 316708
rect 355068 316232 355124 316988
rect 181234 315980 181244 316036
rect 181300 315980 190120 316036
rect 339864 315756 344540 315812
rect 344596 315756 344606 315812
rect 186386 314860 186396 314916
rect 186452 314860 190120 314916
rect 339864 314860 346108 314916
rect 346164 314860 346174 314916
rect 339864 313964 341292 314020
rect 341348 313964 341358 314020
rect 177986 313740 177996 313796
rect 178052 313740 190120 313796
rect 4274 313292 4284 313348
rect 4340 313292 168924 313348
rect 168980 313292 168990 313348
rect 339864 313068 350812 313124
rect 350868 313068 350878 313124
rect 179666 312620 179676 312676
rect 179732 312620 190120 312676
rect 350354 312508 350364 312564
rect 350420 312508 352380 312564
rect 352436 312508 352446 312564
rect 339864 312172 344764 312228
rect 344820 312172 344830 312228
rect 184370 311500 184380 311556
rect 184436 311500 190120 311556
rect 339864 311276 340396 311332
rect 340452 311276 340462 311332
rect 590706 311276 590716 311332
rect 590772 311304 595672 311332
rect 590772 311276 597000 311304
rect 595560 311080 597000 311276
rect 190418 310380 190428 310436
rect 190484 310380 190494 310436
rect 339864 310380 341404 310436
rect 341460 310380 341470 310436
rect 352370 310156 352380 310212
rect 352436 310156 353500 310212
rect 353556 310156 355096 310212
rect 339266 309484 339276 309540
rect 339332 309484 339342 309540
rect 181010 309260 181020 309316
rect 181076 309260 190120 309316
rect 345538 309036 345548 309092
rect 345604 309036 352380 309092
rect 352436 309036 352446 309092
rect 339864 308588 346892 308644
rect 346948 308588 346958 308644
rect 189522 308140 189532 308196
rect 189588 308140 190120 308196
rect 339864 307692 344428 307748
rect 344484 307692 344494 307748
rect 181122 307020 181132 307076
rect 181188 307020 190120 307076
rect 339864 306796 354508 306852
rect 354564 306796 354574 306852
rect 182690 305900 182700 305956
rect 182756 305900 190120 305956
rect 339864 305900 354060 305956
rect 354116 305900 354126 305956
rect -960 304948 480 305144
rect 339864 305004 342300 305060
rect 342356 305004 342366 305060
rect -960 304920 165452 304948
rect 392 304892 165452 304920
rect 165508 304892 165518 304948
rect 186162 304780 186172 304836
rect 186228 304780 190120 304836
rect 339836 304332 349468 304388
rect 339836 304136 339892 304332
rect 349412 304276 349468 304332
rect 349412 304220 354732 304276
rect 354788 304220 354798 304276
rect 352370 304108 352380 304164
rect 352436 304108 354844 304164
rect 354900 304108 355096 304164
rect 187730 303660 187740 303716
rect 187796 303660 190120 303716
rect 339864 303212 350476 303268
rect 350532 303212 350542 303268
rect 187954 302540 187964 302596
rect 188020 302540 190120 302596
rect 339864 302316 342188 302372
rect 342244 302316 342254 302372
rect 10994 301532 11004 301588
rect 11060 301532 175532 301588
rect 175588 301532 175598 301588
rect 177874 301420 177884 301476
rect 177940 301420 190120 301476
rect 339864 301420 345436 301476
rect 345492 301420 345502 301476
rect 339864 300524 353948 300580
rect 354004 300524 354014 300580
rect 187170 300300 187180 300356
rect 187236 300300 190120 300356
rect 339864 299628 345212 299684
rect 345268 299628 345278 299684
rect 187506 299180 187516 299236
rect 187572 299180 190120 299236
rect 344418 299068 344428 299124
rect 344484 299068 345548 299124
rect 345604 299068 345614 299124
rect 341394 298956 341404 299012
rect 341460 298956 342636 299012
rect 342692 298956 342702 299012
rect 339864 298732 341852 298788
rect 341908 298732 341918 298788
rect 179554 298060 179564 298116
rect 179620 298060 190120 298116
rect 339378 298060 339388 298116
rect 339444 298060 353948 298116
rect 354004 298060 355096 298116
rect 590594 298060 590604 298116
rect 590660 298088 595672 298116
rect 590660 298060 597000 298088
rect 339864 297836 351148 297892
rect 351204 297836 351214 297892
rect 595560 297864 597000 298060
rect 186946 296940 186956 296996
rect 187012 296940 190120 296996
rect 339826 296940 339836 296996
rect 339892 296940 339902 296996
rect 4386 296492 4396 296548
rect 4452 296492 177212 296548
rect 177268 296492 177278 296548
rect 186498 296492 186508 296548
rect 186564 296492 187068 296548
rect 187124 296492 187134 296548
rect 339864 296044 340732 296100
rect 340788 296044 340798 296100
rect 187842 295820 187852 295876
rect 187908 295820 190120 295876
rect 339836 295596 339948 295652
rect 340004 295596 340014 295652
rect 339836 295204 339892 295596
rect 339836 295176 348012 295204
rect 339864 295148 348012 295176
rect 348068 295148 348078 295204
rect 161298 294812 161308 294868
rect 161364 294812 177212 294868
rect 177268 294812 177278 294868
rect 186050 294700 186060 294756
rect 186116 294700 190120 294756
rect 339864 294252 341180 294308
rect 341236 294252 349580 294308
rect 349636 294252 349646 294308
rect 59042 293916 59052 293972
rect 59108 293916 60396 293972
rect 60452 293916 60462 293972
rect 46274 293132 46284 293188
rect 46340 293132 51660 293188
rect 51716 293132 87276 293188
rect 87332 293132 87342 293188
rect 190652 293076 190708 293608
rect 339836 293188 339892 293384
rect 339836 293132 343420 293188
rect 343476 293132 353388 293188
rect 353444 293132 353454 293188
rect 190642 293020 190652 293076
rect 190708 293020 190718 293076
rect 7522 292460 7532 292516
rect 7588 292460 190120 292516
rect 339864 292460 343308 292516
rect 343364 292460 349468 292516
rect 40226 292348 40236 292404
rect 40292 292348 46284 292404
rect 46340 292348 46350 292404
rect 71782 292348 71820 292404
rect 71876 292348 71886 292404
rect 84550 292348 84588 292404
rect 84644 292348 84654 292404
rect 349412 292348 349468 292460
rect 349524 292348 349534 292404
rect 352034 292012 352044 292068
rect 352100 292012 355180 292068
rect 355236 292012 355246 292068
rect 339602 291564 339612 291620
rect 339668 291564 347788 291620
rect 347844 291564 347854 291620
rect 349412 291452 352828 291508
rect 352884 291452 352894 291508
rect 349412 291396 349468 291452
rect 10882 291340 10892 291396
rect 10948 291340 190120 291396
rect 339836 291340 343196 291396
rect 343252 291340 349468 291396
rect 392 291032 4284 291060
rect -960 291004 4284 291032
rect 4340 291004 4350 291060
rect -960 290808 480 291004
rect 339836 290696 339892 291340
rect 26002 290556 26012 290612
rect 26068 290556 190148 290612
rect 4274 290444 4284 290500
rect 4340 290444 92316 290500
rect 92372 290444 92382 290500
rect 87266 290332 87276 290388
rect 87332 290332 144284 290388
rect 144340 290332 144350 290388
rect 190092 290248 190148 290556
rect 169138 289884 169148 289940
rect 169204 289884 187292 289940
rect 187348 289884 188076 289940
rect 188132 289884 188142 289940
rect 144274 289772 144284 289828
rect 144340 289772 188076 289828
rect 188132 289772 188142 289828
rect 339864 289772 342748 289828
rect 342804 289772 349692 289828
rect 349748 289772 349758 289828
rect 27682 289100 27692 289156
rect 27748 289100 190120 289156
rect 188066 288988 188076 289044
rect 188132 288988 188972 289044
rect 189028 288988 189038 289044
rect 90888 288876 93996 288932
rect 94052 288876 94062 288932
rect 339714 288876 339724 288932
rect 339780 288876 348572 288932
rect 348628 288876 348638 288932
rect 169250 288092 169260 288148
rect 169316 288092 187404 288148
rect 187460 288092 188076 288148
rect 188132 288092 188142 288148
rect 115042 287980 115052 288036
rect 115108 287980 190120 288036
rect 339836 287364 339892 288008
rect 187030 287308 187068 287364
rect 187124 287308 187134 287364
rect 339836 287308 354620 287364
rect 354676 287308 354686 287364
rect 339864 287084 344316 287140
rect 344372 287084 344382 287140
rect 173842 286860 173852 286916
rect 173908 286860 190120 286916
rect 169362 286524 169372 286580
rect 169428 286524 187516 286580
rect 187572 286524 188076 286580
rect 188132 286524 188142 286580
rect 93986 286412 93996 286468
rect 94052 286412 166348 286468
rect 166404 286412 166414 286468
rect 169026 286412 169036 286468
rect 169092 286412 187068 286468
rect 187124 286412 187740 286468
rect 187796 286412 187806 286468
rect 339266 286188 339276 286244
rect 339332 286216 339864 286244
rect 339332 286188 339892 286216
rect 92306 285740 92316 285796
rect 92372 285740 190120 285796
rect 339836 285684 339892 286188
rect 353490 285964 353500 286020
rect 353556 285964 355096 286020
rect 182242 285628 182252 285684
rect 182308 285628 183932 285684
rect 183988 285628 183998 285684
rect 339836 285628 355628 285684
rect 355684 285628 355694 285684
rect 93986 285404 93996 285460
rect 94052 285404 168028 285460
rect 168084 285404 168094 285460
rect 90860 285292 167468 285348
rect 167524 285292 167534 285348
rect 339864 285292 346444 285348
rect 346500 285292 346510 285348
rect 90860 284648 90916 285292
rect 168914 284732 168924 284788
rect 168980 284732 186508 284788
rect 186564 284732 188076 284788
rect 188132 284732 188142 284788
rect 353378 284732 353388 284788
rect 353444 284732 354396 284788
rect 354452 284732 354462 284788
rect 595560 284676 597000 284872
rect 165442 284620 165452 284676
rect 165508 284620 190120 284676
rect 590482 284620 590492 284676
rect 590548 284648 597000 284676
rect 590548 284620 595672 284648
rect 339864 284396 351260 284452
rect 351316 284396 351326 284452
rect 165928 283948 169148 284004
rect 169204 283948 169214 284004
rect 344754 283836 344764 283892
rect 344820 283836 345996 283892
rect 346052 283836 346062 283892
rect 177202 283500 177212 283556
rect 177268 283500 190120 283556
rect 339864 283500 347900 283556
rect 347956 283500 347966 283556
rect 175634 283052 175644 283108
rect 175700 283052 187628 283108
rect 187684 283052 187694 283108
rect 339864 282604 344764 282660
rect 344820 282604 344830 282660
rect 168914 282380 168924 282436
rect 168980 282380 190120 282436
rect 185714 282156 185724 282212
rect 185780 282156 187292 282212
rect 187348 282156 187358 282212
rect 344866 282156 344876 282212
rect 344932 282156 345884 282212
rect 345940 282156 345950 282212
rect 187030 282044 187068 282100
rect 187124 282044 187134 282100
rect 165928 281932 182252 281988
rect 182308 281932 182318 281988
rect 339714 281708 339724 281764
rect 339780 281708 355516 281764
rect 355572 281708 355582 281764
rect 167122 281260 167132 281316
rect 167188 281260 190120 281316
rect 339864 280812 344204 280868
rect 344260 280812 344270 280868
rect 188038 280588 188076 280644
rect 188132 280588 188142 280644
rect 167458 280476 167468 280532
rect 167524 280476 168140 280532
rect 168196 280476 168206 280532
rect 185602 280476 185612 280532
rect 185668 280476 187628 280532
rect 187684 280476 187694 280532
rect 341254 280476 341292 280532
rect 341348 280476 341358 280532
rect 346098 280476 346108 280532
rect 346164 280476 347228 280532
rect 347284 280476 347294 280532
rect 90888 280364 93996 280420
rect 94052 280364 94062 280420
rect 185938 280364 185948 280420
rect 186004 280364 187404 280420
rect 187460 280364 187470 280420
rect 178882 280140 178892 280196
rect 178948 280140 190120 280196
rect 165928 279916 169260 279972
rect 169316 279916 169326 279972
rect 339864 279916 341404 279972
rect 341460 279916 341470 279972
rect 355068 279412 355124 279944
rect 355058 279356 355068 279412
rect 355124 279356 355134 279412
rect 173012 279132 185948 279188
rect 186004 279132 186014 279188
rect 173012 278964 173068 279132
rect 175522 279020 175532 279076
rect 175588 279020 190120 279076
rect 339864 279020 346220 279076
rect 346276 279020 346286 279076
rect 168130 278908 168140 278964
rect 168196 278908 173068 278964
rect 351250 278908 351260 278964
rect 351316 278908 353836 278964
rect 353892 278908 353902 278964
rect 165928 277900 169372 277956
rect 169428 277900 169438 277956
rect 172162 277900 172172 277956
rect 172228 277900 190120 277956
rect 339836 277508 339892 278152
rect 339836 277452 339948 277508
rect 340004 277452 340014 277508
rect 339836 277060 339892 277256
rect 341170 277228 341180 277284
rect 341236 277228 342524 277284
rect 342580 277228 342590 277284
rect 339836 277004 339948 277060
rect 340004 277004 340014 277060
rect -960 276724 480 276920
rect 175522 276780 175532 276836
rect 175588 276780 190120 276836
rect -960 276696 34412 276724
rect 392 276668 34412 276696
rect 34468 276668 34478 276724
rect 339864 276332 346668 276388
rect 346724 276332 346734 276388
rect 90888 276108 93996 276164
rect 94052 276108 94062 276164
rect 165928 275884 169036 275940
rect 169092 275884 169102 275940
rect 173842 275660 173852 275716
rect 173908 275660 190120 275716
rect 339864 275436 351260 275492
rect 351316 275436 351326 275492
rect 170482 274540 170492 274596
rect 170548 274540 190120 274596
rect 339836 273924 339892 274568
rect 165928 273868 168924 273924
rect 168980 273868 168990 273924
rect 339836 273868 340060 273924
rect 340116 273868 340126 273924
rect 354274 273868 354284 273924
rect 354340 273868 355096 273924
rect 339864 273644 344092 273700
rect 344148 273644 344158 273700
rect 183026 273420 183036 273476
rect 183092 273420 190120 273476
rect 347974 272972 348012 273028
rect 348068 272972 348078 273028
rect 339864 272748 343196 272804
rect 343252 272748 343262 272804
rect 189410 272300 189420 272356
rect 189476 272300 190120 272356
rect 165900 272076 174636 272132
rect 174692 272076 175644 272132
rect 175700 272076 175710 272132
rect 352818 272076 352828 272132
rect 352884 272076 353948 272132
rect 354004 272076 354014 272132
rect 90888 271852 93996 271908
rect 94052 271852 94062 271908
rect 165900 271880 165956 272076
rect 339500 271236 339556 271880
rect 595560 271460 597000 271656
rect 590706 271404 590716 271460
rect 590772 271432 597000 271460
rect 590772 271404 595672 271432
rect 189634 271180 189644 271236
rect 189700 271180 190120 271236
rect 339490 271180 339500 271236
rect 339556 271180 339566 271236
rect 339864 270956 343308 271012
rect 343364 270956 343374 271012
rect 189746 270060 189756 270116
rect 189812 270060 190120 270116
rect 339864 270060 349580 270116
rect 349636 270060 349646 270116
rect 165928 269836 177996 269892
rect 178052 269836 178062 269892
rect 339266 269164 339276 269220
rect 339332 269164 339342 269220
rect 189522 268940 189532 268996
rect 189588 268940 190120 268996
rect 173012 268716 185724 268772
rect 185780 268716 185790 268772
rect 342402 268716 342412 268772
rect 342468 268716 343084 268772
rect 343140 268716 343150 268772
rect 352034 268716 352044 268772
rect 352100 268716 352268 268772
rect 352324 268716 352334 268772
rect 173012 268660 173068 268716
rect 166338 268604 166348 268660
rect 166404 268604 173068 268660
rect 165928 267820 166348 267876
rect 166404 267820 166414 267876
rect 184706 267820 184716 267876
rect 184772 267820 190120 267876
rect 339388 267764 339444 268296
rect 352034 267820 352044 267876
rect 352100 267820 355096 267876
rect 339378 267708 339388 267764
rect 339444 267708 339454 267764
rect 90888 267596 108332 267652
rect 108388 267596 108398 267652
rect 339864 267372 343420 267428
rect 343476 267372 343486 267428
rect 181346 266700 181356 266756
rect 181412 266700 190120 266756
rect 339864 266476 343084 266532
rect 343140 266476 343150 266532
rect 165928 265804 168140 265860
rect 168196 265804 168206 265860
rect 183026 265580 183036 265636
rect 183092 265580 190120 265636
rect 339864 265580 342860 265636
rect 342916 265580 342926 265636
rect 168018 265356 168028 265412
rect 168084 265356 185612 265412
rect 185668 265356 185678 265412
rect 339864 264684 351372 264740
rect 351428 264684 351438 264740
rect 343634 264572 343644 264628
rect 343700 264572 351484 264628
rect 351540 264572 351550 264628
rect 182914 264460 182924 264516
rect 182980 264460 190120 264516
rect 165928 263788 168028 263844
rect 168084 263788 168094 263844
rect 339864 263788 342748 263844
rect 342804 263788 342814 263844
rect 90888 263340 106652 263396
rect 106708 263340 106718 263396
rect 184594 263340 184604 263396
rect 184660 263340 190120 263396
rect 339864 262892 347900 262948
rect 347956 262892 347966 262948
rect 392 262808 4284 262836
rect -960 262780 4284 262808
rect 4340 262780 4350 262836
rect -960 262584 480 262780
rect 344642 262332 344652 262388
rect 344708 262332 345772 262388
rect 345828 262332 345838 262388
rect 186274 262220 186284 262276
rect 186340 262220 190120 262276
rect 344082 262108 344092 262164
rect 344148 262108 345100 262164
rect 345156 262108 345166 262164
rect 339864 261996 342972 262052
rect 343028 261996 343038 262052
rect 165928 261772 168812 261828
rect 168868 261772 168878 261828
rect 352034 261772 352044 261828
rect 352100 261772 352268 261828
rect 352324 261772 355096 261828
rect 351250 261212 351260 261268
rect 351316 261212 351820 261268
rect 351876 261212 351886 261268
rect 184706 261100 184716 261156
rect 184772 261100 190120 261156
rect 339602 261100 339612 261156
rect 339668 261100 339678 261156
rect 339864 260204 349468 260260
rect 349524 260204 349534 260260
rect 187058 259980 187068 260036
rect 187124 259980 190120 260036
rect 190642 259756 190652 259812
rect 190708 259756 190718 259812
rect 90888 259084 92428 259140
rect 92484 259084 92494 259140
rect 190652 258888 190708 259756
rect 339266 259308 339276 259364
rect 339332 259308 339342 259364
rect 344530 258636 344540 258692
rect 344596 258636 345660 258692
rect 345716 258636 345726 258692
rect 339266 258412 339276 258468
rect 339332 258412 339342 258468
rect 590482 258412 590492 258468
rect 590548 258440 595672 258468
rect 590548 258412 597000 258440
rect 595560 258216 597000 258412
rect 187618 257740 187628 257796
rect 187684 257740 190120 257796
rect 339266 257516 339276 257572
rect 339332 257516 339342 257572
rect 342626 256956 342636 257012
rect 342692 256956 344988 257012
rect 345044 256956 345054 257012
rect 345538 256956 345548 257012
rect 345604 256956 345996 257012
rect 346052 256956 346062 257012
rect 351782 256956 351820 257012
rect 351876 256956 351886 257012
rect 352370 256956 352380 257012
rect 352436 256956 352492 257012
rect 352548 256956 352558 257012
rect 339378 256844 339388 256900
rect 339444 256844 340060 256900
rect 340116 256844 340126 256900
rect 190652 255780 190708 256648
rect 339378 256620 339388 256676
rect 339444 256620 339454 256676
rect 341058 256172 341068 256228
rect 341124 256172 342076 256228
rect 342132 256172 342142 256228
rect 190642 255724 190652 255780
rect 190708 255724 190718 255780
rect 339864 255724 346220 255780
rect 346276 255724 346286 255780
rect 352370 255724 352380 255780
rect 352436 255724 355096 255780
rect 187394 255500 187404 255556
rect 187460 255500 190120 255556
rect 90888 254828 93324 254884
rect 93380 254828 93390 254884
rect 339864 254828 344428 254884
rect 344484 254828 344494 254884
rect 187282 254380 187292 254436
rect 187348 254380 190120 254436
rect 339864 253932 348012 253988
rect 348068 253932 348078 253988
rect 339378 253708 339388 253764
rect 339444 253708 340060 253764
rect 340116 253708 340126 253764
rect 190652 252420 190708 253288
rect 339864 253036 344428 253092
rect 344484 253036 344494 253092
rect 345090 252924 345100 252980
rect 345156 252924 354172 252980
rect 354228 252924 354238 252980
rect 345538 252700 345548 252756
rect 345604 252700 350140 252756
rect 350196 252700 350206 252756
rect 344530 252588 344540 252644
rect 344596 252588 349580 252644
rect 349636 252588 349646 252644
rect 190642 252364 190652 252420
rect 190708 252364 190718 252420
rect 188066 252140 188076 252196
rect 188132 252140 190120 252196
rect 339864 252140 340228 252196
rect 340172 252084 340228 252140
rect 340162 252028 340172 252084
rect 340228 252028 340238 252084
rect 349570 252028 349580 252084
rect 349636 252028 350924 252084
rect 350980 252028 350990 252084
rect 352818 252028 352828 252084
rect 352884 252028 353948 252084
rect 354004 252028 354014 252084
rect 339864 251244 344652 251300
rect 344708 251244 344718 251300
rect 187954 251020 187964 251076
rect 188020 251020 190120 251076
rect 90888 250572 93212 250628
rect 93268 250572 93660 250628
rect 93716 250572 93726 250628
rect 339864 250348 341292 250404
rect 341348 250348 341358 250404
rect 343522 250348 343532 250404
rect 343588 250348 346556 250404
rect 346612 250348 346622 250404
rect 340050 250012 340060 250068
rect 340116 250012 341180 250068
rect 341236 250012 341246 250068
rect 352594 249676 352604 249732
rect 352660 249676 355096 249732
rect 339864 249452 342860 249508
rect 342916 249452 342926 249508
rect 349458 249452 349468 249508
rect 349524 249452 351036 249508
rect 351092 249452 351102 249508
rect -960 248500 480 248696
rect 339864 248556 343196 248612
rect 343252 248556 343262 248612
rect -960 248472 40908 248500
rect 392 248444 40908 248472
rect 40964 248444 40974 248500
rect 342514 248444 342524 248500
rect 342580 248444 346332 248500
rect 346388 248444 346398 248500
rect 342178 248220 342188 248276
rect 342244 248220 350812 248276
rect 350868 248220 350878 248276
rect 339378 247884 339388 247940
rect 339444 247884 350364 247940
rect 350420 247884 350430 247940
rect 342514 247772 342524 247828
rect 342580 247772 349692 247828
rect 349748 247772 349758 247828
rect 339266 247660 339276 247716
rect 339332 247660 339342 247716
rect 340386 246988 340396 247044
rect 340452 246988 342524 247044
rect 342580 246988 342590 247044
rect 341254 246876 341292 246932
rect 341348 246876 341358 246932
rect 347778 246876 347788 246932
rect 347844 246876 349356 246932
rect 349412 246876 349422 246932
rect 339266 246764 339276 246820
rect 339332 246764 339342 246820
rect 344316 246764 346444 246820
rect 346500 246764 350252 246820
rect 350308 246764 350318 246820
rect 344316 246708 344372 246764
rect 340274 246652 340284 246708
rect 340340 246652 344372 246708
rect 344530 246652 344540 246708
rect 344596 246652 350700 246708
rect 350756 246652 350766 246708
rect 340274 246540 340284 246596
rect 340340 246540 348460 246596
rect 348516 246540 348526 246596
rect 90888 246316 93324 246372
rect 93380 246316 93436 246372
rect 93492 246316 93502 246372
rect 339864 245868 346108 245924
rect 346164 245868 346174 245924
rect 339378 245308 339388 245364
rect 339444 245308 340956 245364
rect 341012 245308 341022 245364
rect 344614 245196 344652 245252
rect 344708 245196 344718 245252
rect 345874 245196 345884 245252
rect 345940 245196 347788 245252
rect 347844 245196 347854 245252
rect 351782 245196 351820 245252
rect 351876 245196 351886 245252
rect 352482 245196 352492 245252
rect 352548 245196 352716 245252
rect 352772 245196 352782 245252
rect 339378 245084 339388 245140
rect 339444 245084 344540 245140
rect 344596 245084 344606 245140
rect 595560 245028 597000 245224
rect 590594 244972 590604 245028
rect 590660 245000 597000 245028
rect 590660 244972 595672 245000
rect 339378 244860 339388 244916
rect 339444 244860 349244 244916
rect 349300 244860 349310 244916
rect 341394 243628 341404 243684
rect 341460 243628 348796 243684
rect 348852 243628 348862 243684
rect 352482 243628 352492 243684
rect 352548 243628 355096 243684
rect 90888 242060 93492 242116
rect 93436 242004 93492 242060
rect 93398 241948 93436 242004
rect 93492 241948 93502 242004
rect 339378 241948 339388 242004
rect 339444 241948 339948 242004
rect 340004 241948 340014 242004
rect 340946 241948 340956 242004
rect 341012 241948 342524 242004
rect 342580 241948 342590 242004
rect 340386 241500 340396 241556
rect 340452 241500 348012 241556
rect 348068 241500 348078 241556
rect 90178 241164 90188 241220
rect 90244 241164 116732 241220
rect 116788 241164 116798 241220
rect 85652 241052 111692 241108
rect 111748 241052 111758 241108
rect 70532 240940 80444 240996
rect 80500 240940 80510 240996
rect 70532 240884 70588 240940
rect 85652 240884 85708 241052
rect 66220 240828 70588 240884
rect 71596 240828 85708 240884
rect 66220 240772 66276 240828
rect 71596 240772 71652 240828
rect 38434 240716 38444 240772
rect 38500 240716 41132 240772
rect 41188 240716 41198 240772
rect 66210 240716 66220 240772
rect 66276 240716 66286 240772
rect 71586 240716 71596 240772
rect 71652 240716 71662 240772
rect 80434 240716 80444 240772
rect 80500 240716 118412 240772
rect 118468 240716 118478 240772
rect 80546 240604 80556 240660
rect 80612 240604 90188 240660
rect 90244 240604 90254 240660
rect 339714 240604 339724 240660
rect 339780 240604 347900 240660
rect 347956 240604 347966 240660
rect 60834 240492 60844 240548
rect 60900 240492 232764 240548
rect 232820 240492 232830 240548
rect 236114 240492 236124 240548
rect 236180 240492 337708 240548
rect 338930 240492 338940 240548
rect 338996 240492 347900 240548
rect 347956 240492 347966 240548
rect 57250 240380 57260 240436
rect 57316 240380 185612 240436
rect 185668 240380 185678 240436
rect 337652 240324 337708 240492
rect 338594 240380 338604 240436
rect 338660 240380 349468 240436
rect 349524 240380 349534 240436
rect 53666 240268 53676 240324
rect 53732 240268 170604 240324
rect 170660 240268 170670 240324
rect 337652 240268 338548 240324
rect 338706 240268 338716 240324
rect 338772 240268 344652 240324
rect 344708 240268 344718 240324
rect 347890 240268 347900 240324
rect 347956 240268 349244 240324
rect 349300 240268 349310 240324
rect 338492 240212 338548 240268
rect 46498 240156 46508 240212
rect 46564 240156 67228 240212
rect 85922 240156 85932 240212
rect 85988 240156 168812 240212
rect 168868 240156 168878 240212
rect 188962 240156 188972 240212
rect 189028 240156 194908 240212
rect 194964 240156 194974 240212
rect 338492 240156 339724 240212
rect 339780 240156 339790 240212
rect 339910 240156 339948 240212
rect 340004 240156 340014 240212
rect 340834 240156 340844 240212
rect 340900 240156 346220 240212
rect 346276 240156 346286 240212
rect 67172 240100 67228 240156
rect 55458 240044 55468 240100
rect 55524 240044 55534 240100
rect 67172 240044 167132 240100
rect 167188 240044 167198 240100
rect 55468 239988 55524 240044
rect 55468 239932 113372 239988
rect 113428 239932 113438 239988
rect 185938 239932 185948 239988
rect 186004 239932 341404 239988
rect 341460 239932 341470 239988
rect 82338 239820 82348 239876
rect 82404 239820 120092 239876
rect 120148 239820 120158 239876
rect 238466 239820 238476 239876
rect 238532 239820 273420 239876
rect 273476 239820 273486 239876
rect 287970 239820 287980 239876
rect 288036 239820 343420 239876
rect 343476 239820 343486 239876
rect 241826 239708 241836 239764
rect 241892 239708 276332 239764
rect 276388 239708 276398 239764
rect 281362 239708 281372 239764
rect 281428 239708 342748 239764
rect 342804 239708 342814 239764
rect 187170 239596 187180 239652
rect 187236 239596 273980 239652
rect 274036 239596 274046 239652
rect 279682 239596 279692 239652
rect 279748 239596 343084 239652
rect 343140 239596 343150 239652
rect 179554 239484 179564 239540
rect 179620 239484 272972 239540
rect 273028 239484 273038 239540
rect 314132 239484 340956 239540
rect 341012 239484 341022 239540
rect 342626 239484 342636 239540
rect 342692 239484 351820 239540
rect 351876 239484 351886 239540
rect 314132 239428 314188 239484
rect 230962 239372 230972 239428
rect 231028 239372 314188 239428
rect 236786 239260 236796 239316
rect 236852 239260 289100 239316
rect 289156 239260 289166 239316
rect 289986 239260 289996 239316
rect 290052 239260 343308 239316
rect 343364 239260 343374 239316
rect 185714 239148 185724 239204
rect 185780 239148 344540 239204
rect 344596 239148 344606 239204
rect 288306 239036 288316 239092
rect 288372 239036 342972 239092
rect 343028 239036 343038 239092
rect 278002 238924 278012 238980
rect 278068 238924 344092 238980
rect 344148 238924 344158 238980
rect 343522 238700 343532 238756
rect 343588 238700 344428 238756
rect 344484 238700 344494 238756
rect 343746 238588 343756 238644
rect 343812 238588 344428 238644
rect 344484 238588 344494 238644
rect 349122 238588 349132 238644
rect 349188 238588 352828 238644
rect 352884 238588 354172 238644
rect 354228 238588 354238 238644
rect 38546 238476 38556 238532
rect 38612 238476 42924 238532
rect 42980 238476 42990 238532
rect 62598 238476 62636 238532
rect 62692 238476 62702 238532
rect 64390 238476 64428 238532
rect 64484 238476 64494 238532
rect 87714 238476 87724 238532
rect 87780 238476 95340 238532
rect 95396 238476 95406 238532
rect 244150 238476 244188 238532
rect 244244 238476 244254 238532
rect 245046 238476 245084 238532
rect 245140 238476 245150 238532
rect 252242 238476 252252 238532
rect 252308 238476 269724 238532
rect 269780 238476 269790 238532
rect 289090 238476 289100 238532
rect 289156 238476 337708 238532
rect 340022 238476 340060 238532
rect 340116 238476 340126 238532
rect 40674 238364 40684 238420
rect 40740 238364 51884 238420
rect 51940 238364 51950 238420
rect 84130 238364 84140 238420
rect 84196 238364 99932 238420
rect 99988 238364 99998 238420
rect 250450 238364 250460 238420
rect 250516 238364 270508 238420
rect 270564 238364 270574 238420
rect 337652 238308 337708 238476
rect 38210 238252 38220 238308
rect 38276 238252 44716 238308
rect 44772 238252 44782 238308
rect 89506 238252 89516 238308
rect 89572 238252 95116 238308
rect 95172 238252 95182 238308
rect 246866 238252 246876 238308
rect 246932 238252 270508 238308
rect 270564 238252 270574 238308
rect 272850 238252 272860 238308
rect 272916 238252 291564 238308
rect 291620 238252 291630 238308
rect 337652 238252 355068 238308
rect 355124 238252 355516 238308
rect 355572 238252 355582 238308
rect 38322 238140 38332 238196
rect 38388 238140 48300 238196
rect 48356 238140 48366 238196
rect 69794 238140 69804 238196
rect 69860 238140 95564 238196
rect 95620 238140 95630 238196
rect 251346 238140 251356 238196
rect 251412 238140 275660 238196
rect 275716 238140 275726 238196
rect 76962 238028 76972 238084
rect 77028 238028 94892 238084
rect 94948 238028 94958 238084
rect 249554 238028 249564 238084
rect 249620 238028 273980 238084
rect 274036 238028 274046 238084
rect 321234 238028 321244 238084
rect 321300 238028 337372 238084
rect 337428 238028 337438 238084
rect 39666 237916 39676 237972
rect 39732 237916 50092 237972
rect 50148 237916 50158 237972
rect 73378 237916 73388 237972
rect 73444 237916 103292 237972
rect 103348 237916 103358 237972
rect 248658 237916 248668 237972
rect 248724 237916 274092 237972
rect 274148 237916 274158 237972
rect 300402 237916 300412 237972
rect 300468 237916 307804 237972
rect 307860 237916 307870 237972
rect 320338 237916 320348 237972
rect 320404 237916 337148 237972
rect 337204 237916 337214 237972
rect 337820 237916 343196 237972
rect 343252 237916 343262 237972
rect 75170 237804 75180 237860
rect 75236 237804 104972 237860
rect 105028 237804 105038 237860
rect 247762 237804 247772 237860
rect 247828 237804 280588 237860
rect 280644 237804 280654 237860
rect 298946 237804 298956 237860
rect 299012 237804 303324 237860
rect 303380 237804 303390 237860
rect 314066 237804 314076 237860
rect 314132 237804 337596 237860
rect 337652 237804 337662 237860
rect 337820 237748 337876 237916
rect 78754 237692 78764 237748
rect 78820 237692 96572 237748
rect 96628 237692 96638 237748
rect 245970 237692 245980 237748
rect 246036 237692 278908 237748
rect 278964 237692 278974 237748
rect 284722 237692 284732 237748
rect 284788 237692 337876 237748
rect 340498 237692 340508 237748
rect 340564 237692 342188 237748
rect 342244 237692 342254 237748
rect 68002 237580 68012 237636
rect 68068 237580 96796 237636
rect 96852 237580 96862 237636
rect 273746 237580 273756 237636
rect 273812 237580 279916 237636
rect 279972 237580 279982 237636
rect 287186 237580 287196 237636
rect 287252 237580 293244 237636
rect 293300 237580 293310 237636
rect 340386 237580 340396 237636
rect 340452 237580 340956 237636
rect 341012 237580 355096 237636
rect 253138 237468 253148 237524
rect 253204 237468 269612 237524
rect 269668 237468 269678 237524
rect 282706 237468 282716 237524
rect 282772 237468 291788 237524
rect 291844 237468 291854 237524
rect 300514 237468 300524 237524
rect 300580 237468 305116 237524
rect 305172 237468 305182 237524
rect 297154 237356 297164 237412
rect 297220 237356 302428 237412
rect 302484 237356 302494 237412
rect 297266 237244 297276 237300
rect 297332 237244 306012 237300
rect 306068 237244 306078 237300
rect 235218 237020 235228 237076
rect 235284 237020 236796 237076
rect 236852 237020 236862 237076
rect 242386 237020 242396 237076
rect 242452 237020 243404 237076
rect 243460 237020 243470 237076
rect 267474 237020 267484 237076
rect 267540 237020 268716 237076
rect 268772 237020 268782 237076
rect 208338 236908 208348 236964
rect 208404 236908 209916 236964
rect 209972 236908 209982 236964
rect 225138 236908 225148 236964
rect 225204 236908 226268 236964
rect 226324 236908 226334 236964
rect 233398 236908 233436 236964
rect 233492 236908 233502 236964
rect 236646 236908 236684 236964
rect 236740 236908 236750 236964
rect 237010 236908 237020 236964
rect 237076 236908 238476 236964
rect 238532 236908 238542 236964
rect 238802 236908 238812 236964
rect 238868 236908 240044 236964
rect 240100 236908 240110 236964
rect 240594 236908 240604 236964
rect 240660 236908 241836 236964
rect 241892 236908 241902 236964
rect 243478 236908 243516 236964
rect 243572 236908 243582 236964
rect 266998 236908 267036 236964
rect 267092 236908 267102 236964
rect 268566 236908 268604 236964
rect 268660 236908 268670 236964
rect 280914 236908 280924 236964
rect 280980 236908 288428 236964
rect 288484 236908 288494 236964
rect 290770 236908 290780 236964
rect 290836 236908 294924 236964
rect 294980 236908 294990 236964
rect 301522 236908 301532 236964
rect 301588 236908 302316 236964
rect 302372 236908 302382 236964
rect 303426 236908 303436 236964
rect 303492 236908 304220 236964
rect 304276 236908 304286 236964
rect 307318 236908 307356 236964
rect 307412 236908 307422 236964
rect 308998 236908 309036 236964
rect 309092 236908 309102 236964
rect 309586 236908 309596 236964
rect 309652 236908 310716 236964
rect 310772 236908 310782 236964
rect 317650 236908 317660 236964
rect 317716 236908 319116 236964
rect 319172 236908 319182 236964
rect 334198 236908 334236 236964
rect 334292 236908 334302 236964
rect 334674 236908 334684 236964
rect 334740 236908 335916 236964
rect 335972 236908 335982 236964
rect 168802 236796 168812 236852
rect 168868 236796 339388 236852
rect 339444 236796 339948 236852
rect 340004 236796 340014 236852
rect 353490 236796 353500 236852
rect 353556 236796 354284 236852
rect 354340 236796 354350 236852
rect 182242 236684 182252 236740
rect 182308 236684 349468 236740
rect 349412 236628 349468 236684
rect 185602 236572 185612 236628
rect 185668 236572 345660 236628
rect 345716 236572 345726 236628
rect 349412 236572 352940 236628
rect 352996 236572 355404 236628
rect 355460 236572 355470 236628
rect 239474 236460 239484 236516
rect 239540 236460 351260 236516
rect 351316 236460 351326 236516
rect 236002 236348 236012 236404
rect 236068 236348 341068 236404
rect 341124 236348 341134 236404
rect 236226 236236 236236 236292
rect 236292 236236 340284 236292
rect 340340 236236 340350 236292
rect 35186 236124 35196 236180
rect 35252 236124 343196 236180
rect 343252 236124 343262 236180
rect 33506 236012 33516 236068
rect 33572 236012 342860 236068
rect 342916 236012 342926 236068
rect 41010 235116 41020 235172
rect 41076 235116 241500 235172
rect 241556 235116 272300 235172
rect 272356 235116 272366 235172
rect 240146 235004 240156 235060
rect 240212 235004 283052 235060
rect 283108 235004 283118 235060
rect 186274 234892 186284 234948
rect 186340 234892 302764 234948
rect 302820 234892 302830 234948
rect 179218 234780 179228 234836
rect 179284 234780 307244 234836
rect 307300 234780 307310 234836
rect 179442 234668 179452 234724
rect 179508 234668 328524 234724
rect 328580 234668 328590 234724
rect -960 234388 480 234584
rect 43474 234556 43484 234612
rect 43540 234556 207452 234612
rect 207508 234556 207518 234612
rect 241714 234556 241724 234612
rect 241780 234556 280700 234612
rect 280756 234556 280766 234612
rect 283042 234556 283052 234612
rect 283108 234556 351372 234612
rect 351428 234556 351438 234612
rect 41010 234444 41020 234500
rect 41076 234444 205660 234500
rect 205716 234444 205726 234500
rect 223570 234444 223580 234500
rect 223636 234444 266924 234500
rect 266980 234444 266990 234500
rect 273746 234444 273756 234500
rect 273812 234444 354060 234500
rect 354116 234444 354126 234500
rect -960 234360 12572 234388
rect 392 234332 12572 234360
rect 12628 234332 12638 234388
rect 41122 234332 41132 234388
rect 41188 234332 206556 234388
rect 206612 234332 206622 234388
rect 239922 234332 239932 234388
rect 239988 234332 344316 234388
rect 344372 234332 354620 234388
rect 354676 234332 354686 234388
rect 234322 234220 234332 234276
rect 234388 234220 270060 234276
rect 270116 234220 270126 234276
rect 354050 234108 354060 234164
rect 354116 234108 354620 234164
rect 354676 234108 354686 234164
rect 59042 233436 59052 233492
rect 59108 233436 235228 233492
rect 235284 233436 235294 233492
rect 283042 233436 283052 233492
rect 283108 233436 352156 233492
rect 352212 233436 352222 233492
rect 175970 233212 175980 233268
rect 176036 233212 308364 233268
rect 308420 233212 308430 233268
rect 182690 233100 182700 233156
rect 182756 233100 321804 233156
rect 321860 233100 321870 233156
rect 177874 232988 177884 233044
rect 177940 232988 331884 233044
rect 331940 232988 331950 233044
rect 22754 232876 22764 232932
rect 22820 232876 196700 232932
rect 196756 232876 196766 232932
rect 239698 232876 239708 232932
rect 239764 232876 270620 232932
rect 270676 232876 270686 232932
rect 38546 232764 38556 232820
rect 38612 232764 228060 232820
rect 228116 232764 228126 232820
rect 237906 232764 237916 232820
rect 237972 232764 271068 232820
rect 271124 232764 271134 232820
rect 34178 232652 34188 232708
rect 34244 232652 339276 232708
rect 339332 232652 339342 232708
rect 595560 231924 597000 232008
rect 590930 231868 590940 231924
rect 590996 231868 597000 231924
rect 210130 231756 210140 231812
rect 210196 231756 267260 231812
rect 267316 231756 267326 231812
rect 595560 231784 597000 231868
rect 211922 231644 211932 231700
rect 211988 231644 269500 231700
rect 269556 231644 269566 231700
rect 209234 231532 209244 231588
rect 209300 231532 267484 231588
rect 267540 231532 267550 231588
rect 351810 231532 351820 231588
rect 351876 231532 355096 231588
rect 211026 231420 211036 231476
rect 211092 231420 269612 231476
rect 269668 231420 269678 231476
rect 179330 231308 179340 231364
rect 179396 231308 320684 231364
rect 320740 231308 320750 231364
rect 176082 231196 176092 231252
rect 176148 231196 327404 231252
rect 327460 231196 327470 231252
rect 176194 231084 176204 231140
rect 176260 231084 335244 231140
rect 335300 231084 335310 231140
rect 93426 230972 93436 231028
rect 93492 230972 271292 231028
rect 271348 230972 271358 231028
rect 212818 230860 212828 230916
rect 212884 230860 269388 230916
rect 269444 230860 269454 230916
rect 174402 229964 174412 230020
rect 174468 229964 310604 230020
rect 310660 229964 310670 230020
rect 189298 229852 189308 229908
rect 189364 229852 330764 229908
rect 330820 229852 330830 229908
rect 181122 229740 181132 229796
rect 181188 229740 322924 229796
rect 322980 229740 322990 229796
rect 181346 229628 181356 229684
rect 181412 229628 333004 229684
rect 333060 229628 333070 229684
rect 43586 229516 43596 229572
rect 43652 229516 203868 229572
rect 203924 229516 203934 229572
rect 93202 229404 93212 229460
rect 93268 229404 335132 229460
rect 335188 229404 335198 229460
rect 18946 229292 18956 229348
rect 19012 229292 346668 229348
rect 346724 229292 346734 229348
rect 216402 228396 216412 228452
rect 216468 228396 270844 228452
rect 270900 228396 270910 228452
rect 215506 228284 215516 228340
rect 215572 228284 270956 228340
rect 271012 228284 271022 228340
rect 181010 228172 181020 228228
rect 181076 228172 315084 228228
rect 315140 228172 315150 228228
rect 177762 228060 177772 228116
rect 177828 228060 325164 228116
rect 325220 228060 325230 228116
rect 184594 227948 184604 228004
rect 184660 227948 334124 228004
rect 334180 227948 334190 228004
rect 40898 227836 40908 227892
rect 40964 227836 199388 227892
rect 199444 227836 199454 227892
rect 214610 227836 214620 227892
rect 214676 227836 271180 227892
rect 271236 227836 271246 227892
rect 37986 227724 37996 227780
rect 38052 227724 198492 227780
rect 198548 227724 198558 227780
rect 213714 227724 213724 227780
rect 213780 227724 270732 227780
rect 270788 227724 270798 227780
rect 93314 227612 93324 227668
rect 93380 227612 274764 227668
rect 274820 227612 274830 227668
rect 217298 227500 217308 227556
rect 217364 227500 269388 227556
rect 269444 227500 269454 227556
rect 43362 225932 43372 225988
rect 43428 225932 232540 225988
rect 232596 225932 232606 225988
rect 352034 225484 352044 225540
rect 352100 225484 355096 225540
rect 219090 225036 219100 225092
rect 219156 225036 270620 225092
rect 270676 225036 270686 225092
rect 190418 224924 190428 224980
rect 190484 224924 272860 224980
rect 272916 224924 272926 224980
rect 172946 224812 172956 224868
rect 173012 224812 311724 224868
rect 311780 224812 311790 224868
rect 179554 224700 179564 224756
rect 179620 224700 319564 224756
rect 319620 224700 319630 224756
rect 176306 224588 176316 224644
rect 176372 224588 329644 224644
rect 329700 224588 329710 224644
rect 40674 224476 40684 224532
rect 40740 224476 200284 224532
rect 200340 224476 200350 224532
rect 221778 224476 221788 224532
rect 221844 224476 275884 224532
rect 275940 224476 275950 224532
rect 40786 224364 40796 224420
rect 40852 224364 204764 224420
rect 204820 224364 204830 224420
rect 220882 224364 220892 224420
rect 220948 224364 275996 224420
rect 276052 224364 276062 224420
rect 13234 224252 13244 224308
rect 13300 224252 195804 224308
rect 195860 224252 195870 224308
rect 219986 224252 219996 224308
rect 220052 224252 275772 224308
rect 275828 224252 275838 224308
rect 218194 224140 218204 224196
rect 218260 224140 269500 224196
rect 269556 224140 269566 224196
rect 187282 223020 187292 223076
rect 187348 223020 296604 223076
rect 296660 223020 296670 223076
rect 174514 222908 174524 222964
rect 174580 222908 305004 222964
rect 305060 222908 305070 222964
rect 181234 222796 181244 222852
rect 181300 222796 318444 222852
rect 318500 222796 318510 222852
rect 36866 222684 36876 222740
rect 36932 222684 202972 222740
rect 203028 222684 203038 222740
rect 217634 222684 217644 222740
rect 217700 222684 301532 222740
rect 301588 222684 301598 222740
rect 4274 222572 4284 222628
rect 4340 222572 173852 222628
rect 173908 222572 173918 222628
rect 179666 222572 179676 222628
rect 179732 222572 324044 222628
rect 324100 222572 324110 222628
rect 224466 221564 224476 221620
rect 224532 221564 276108 221620
rect 276164 221564 276174 221620
rect 222674 221452 222684 221508
rect 222740 221452 276220 221508
rect 276276 221452 276286 221508
rect 187730 221340 187740 221396
rect 187796 221340 274428 221396
rect 274484 221340 274494 221396
rect 174626 221228 174636 221284
rect 174692 221228 306124 221284
rect 306180 221228 306190 221284
rect 177986 221116 177996 221172
rect 178052 221116 326284 221172
rect 326340 221116 326350 221172
rect 39890 221004 39900 221060
rect 39956 221004 227164 221060
rect 227220 221004 227230 221060
rect 41010 220892 41020 220948
rect 41076 220892 338380 220948
rect 338436 220892 338446 220948
rect 392 220472 4284 220500
rect -960 220444 4284 220472
rect 4340 220444 4350 220500
rect -960 220248 480 220444
rect 239362 219884 239372 219940
rect 239428 219884 301644 219940
rect 301700 219884 301710 219940
rect 214274 219772 214284 219828
rect 214340 219772 286412 219828
rect 286468 219772 286478 219828
rect 187506 219660 187516 219716
rect 187572 219660 271180 219716
rect 271236 219660 271246 219716
rect 182578 219548 182588 219604
rect 182644 219548 303884 219604
rect 303940 219548 303950 219604
rect 189186 219436 189196 219492
rect 189252 219436 313964 219492
rect 314020 219436 314030 219492
rect 352146 219436 352156 219492
rect 352212 219436 355096 219492
rect 182914 219324 182924 219380
rect 182980 219324 316204 219380
rect 316260 219324 316270 219380
rect 187394 219212 187404 219268
rect 187460 219212 337036 219268
rect 337092 219212 337102 219268
rect 592274 218764 592284 218820
rect 592340 218792 595672 218820
rect 592340 218764 597000 218792
rect 595560 218568 597000 218764
rect 184370 218092 184380 218148
rect 184436 218092 272524 218148
rect 272580 218092 272590 218148
rect 187954 217980 187964 218036
rect 188020 217980 289772 218036
rect 289828 217980 289838 218036
rect 189074 217868 189084 217924
rect 189140 217868 301644 217924
rect 301700 217868 301710 217924
rect 186386 217756 186396 217812
rect 186452 217756 312844 217812
rect 312900 217756 312910 217812
rect 154914 217644 154924 217700
rect 154980 217644 167244 217700
rect 167300 217644 167310 217700
rect 184482 217644 184492 217700
rect 184548 217644 317324 217700
rect 317380 217644 317390 217700
rect 38434 217532 38444 217588
rect 38500 217532 201180 217588
rect 201236 217532 201246 217588
rect 262098 216636 262108 216692
rect 262164 216636 289660 216692
rect 289716 216636 289726 216692
rect 259410 216524 259420 216580
rect 259476 216524 288316 216580
rect 288372 216524 288382 216580
rect 239698 216412 239708 216468
rect 239764 216412 274652 216468
rect 274708 216412 274718 216468
rect 214162 216300 214172 216356
rect 214228 216300 290332 216356
rect 290388 216300 290398 216356
rect 210802 216188 210812 216244
rect 210868 216188 290108 216244
rect 290164 216188 290174 216244
rect 177874 216076 177884 216132
rect 177940 216076 272636 216132
rect 272692 216076 272702 216132
rect 182802 215964 182812 216020
rect 182868 215964 309484 216020
rect 309540 215964 309550 216020
rect 35186 215852 35196 215908
rect 35252 215852 228956 215908
rect 229012 215852 229022 215908
rect 255826 215852 255836 215908
rect 255892 215852 293132 215908
rect 293188 215852 293198 215908
rect 254034 214956 254044 215012
rect 254100 214956 281372 215012
rect 281428 214956 281438 215012
rect 181010 214844 181020 214900
rect 181076 214844 272300 214900
rect 272356 214844 272366 214900
rect 188066 214732 188076 214788
rect 188132 214732 286524 214788
rect 286580 214732 286590 214788
rect 203186 214620 203196 214676
rect 203252 214620 336924 214676
rect 336980 214620 336990 214676
rect 187618 214508 187628 214564
rect 187684 214508 337372 214564
rect 337428 214508 337438 214564
rect 40898 214396 40908 214452
rect 40964 214396 230748 214452
rect 230804 214396 230814 214452
rect 258514 214396 258524 214452
rect 258580 214396 291452 214452
rect 291508 214396 291518 214452
rect 40114 214284 40124 214340
rect 40180 214284 229852 214340
rect 229908 214284 229918 214340
rect 254930 214284 254940 214340
rect 254996 214284 294812 214340
rect 294868 214284 294878 214340
rect 24658 214172 24668 214228
rect 24724 214172 225372 214228
rect 225428 214172 225438 214228
rect 228162 214172 228172 214228
rect 228228 214172 284956 214228
rect 285012 214172 285022 214228
rect 257618 214060 257628 214116
rect 257684 214060 279804 214116
rect 279860 214060 279870 214116
rect 352706 213388 352716 213444
rect 352772 213388 355404 213444
rect 355460 213388 355470 213444
rect 241490 213276 241500 213332
rect 241556 213276 273868 213332
rect 273924 213276 273934 213332
rect 217522 213164 217532 213220
rect 217588 213164 290556 213220
rect 290612 213164 290622 213220
rect 201394 213052 201404 213108
rect 201460 213052 276332 213108
rect 276388 213052 276398 213108
rect 186050 212940 186060 212996
rect 186116 212940 272412 212996
rect 272468 212940 272478 212996
rect 187842 212828 187852 212884
rect 187908 212828 277340 212884
rect 277396 212828 277406 212884
rect 40002 212716 40012 212772
rect 40068 212716 202076 212772
rect 202132 212716 202142 212772
rect 230066 212716 230076 212772
rect 230132 212716 337036 212772
rect 337092 212716 337102 212772
rect 30370 212604 30380 212660
rect 30436 212604 197596 212660
rect 197652 212604 197662 212660
rect 227602 212604 227612 212660
rect 227668 212604 336812 212660
rect 336868 212604 336878 212660
rect 39778 212492 39788 212548
rect 39844 212492 231644 212548
rect 231700 212492 231710 212548
rect 260306 212492 260316 212548
rect 260372 212492 295036 212548
rect 295092 212492 295102 212548
rect 256722 212380 256732 212436
rect 256788 212380 284844 212436
rect 284900 212380 284910 212436
rect 265682 211596 265692 211652
rect 265748 211596 300972 211652
rect 301028 211596 301038 211652
rect 263890 211484 263900 211540
rect 263956 211484 301196 211540
rect 301252 211484 301262 211540
rect 187954 211372 187964 211428
rect 188020 211372 271292 211428
rect 271348 211372 271358 211428
rect 186162 211260 186172 211316
rect 186228 211260 272188 211316
rect 272244 211260 272254 211316
rect 272402 211260 272412 211316
rect 272468 211260 272506 211316
rect 186946 211148 186956 211204
rect 187012 211148 274316 211204
rect 274372 211148 274382 211204
rect 181234 211036 181244 211092
rect 181300 211036 272748 211092
rect 272804 211036 272814 211092
rect 182802 210924 182812 210980
rect 182868 210924 269892 210980
rect 269836 210868 269892 210924
rect 4274 210812 4284 210868
rect 4340 210812 115052 210868
rect 115108 210812 115118 210868
rect 179666 210812 179676 210868
rect 179732 210812 267316 210868
rect 269826 210812 269836 210868
rect 269892 210812 269902 210868
rect 262994 210700 263004 210756
rect 263060 210700 267204 210756
rect 267148 210420 267204 210700
rect 267260 210532 267316 210812
rect 278852 210700 296492 210756
rect 296548 210700 296558 210756
rect 267260 210476 273196 210532
rect 273252 210476 273262 210532
rect 278852 210420 278908 210700
rect 267148 210364 278908 210420
rect 264758 210028 264796 210084
rect 264852 210028 264862 210084
rect 261202 209916 261212 209972
rect 261268 209916 343644 209972
rect 343700 209916 343710 209972
rect 189522 209804 189532 209860
rect 189588 209804 270004 209860
rect 272514 209804 272524 209860
rect 272580 209804 272972 209860
rect 273028 209804 273038 209860
rect 269948 209748 270004 209804
rect 186386 209692 186396 209748
rect 186452 209692 269332 209748
rect 269948 209692 273476 209748
rect 269276 209636 269332 209692
rect 273420 209636 273476 209692
rect 182690 209580 182700 209636
rect 182756 209580 269052 209636
rect 269108 209580 269118 209636
rect 269266 209580 269276 209636
rect 269332 209580 269342 209636
rect 272178 209580 272188 209636
rect 272244 209580 272748 209636
rect 272804 209580 272814 209636
rect 273410 209580 273420 209636
rect 273476 209580 273486 209636
rect 181122 209468 181132 209524
rect 181188 209468 272188 209524
rect 272244 209468 272254 209524
rect 272598 209468 272636 209524
rect 272692 209468 272702 209524
rect 177986 209356 177996 209412
rect 178052 209356 273084 209412
rect 273140 209356 273150 209412
rect 269042 209132 269052 209188
rect 269108 209132 272860 209188
rect 272916 209132 272926 209188
rect 264786 209020 264796 209076
rect 264852 209020 293132 209076
rect 293188 209020 293198 209076
rect 344306 208348 344316 208404
rect 344372 208348 351484 208404
rect 351540 208348 351550 208404
rect 269826 207900 269836 207956
rect 269892 207900 269902 207956
rect 269836 207032 269892 207900
rect 335122 207452 335132 207508
rect 335188 207452 337708 207508
rect 337652 207396 337708 207452
rect 337652 207340 352268 207396
rect 352324 207340 355096 207396
rect -960 206164 480 206360
rect -960 206136 41132 206164
rect 392 206108 41132 206136
rect 41188 206108 41198 206164
rect 300850 205772 300860 205828
rect 300916 205772 326620 205828
rect 326676 205772 326686 205828
rect 595560 205380 597000 205576
rect 590818 205324 590828 205380
rect 590884 205352 597000 205380
rect 590884 205324 595672 205352
rect 269864 204092 272748 204148
rect 272804 204092 272814 204148
rect 298722 204092 298732 204148
rect 298788 204092 329308 204148
rect 329364 204092 329374 204148
rect 272962 203084 272972 203140
rect 273028 203084 280700 203140
rect 280756 203084 280766 203140
rect 272850 202524 272860 202580
rect 272916 202524 273196 202580
rect 273252 202524 273262 202580
rect 272178 202412 272188 202468
rect 272244 202412 273756 202468
rect 273812 202412 273822 202468
rect 269266 201180 269276 201236
rect 269332 201180 269342 201236
rect 316754 201180 316764 201236
rect 316820 201180 339164 201236
rect 339220 201180 339230 201236
rect 313170 201068 313180 201124
rect 313236 201068 342188 201124
rect 342244 201068 342254 201124
rect 314962 200956 314972 201012
rect 315028 200956 344204 201012
rect 344260 200956 344270 201012
rect 298610 200844 298620 200900
rect 298676 200844 332892 200900
rect 332948 200844 332958 200900
rect 355068 200788 355124 201320
rect 274754 200732 274764 200788
rect 274820 200732 351148 200788
rect 351204 200732 355124 200788
rect 272962 199836 272972 199892
rect 273028 199836 276332 199892
rect 276388 199836 276398 199892
rect 300626 199276 300636 199332
rect 300692 199276 323932 199332
rect 323988 199276 323998 199332
rect 298498 199164 298508 199220
rect 298564 199164 328412 199220
rect 328468 199164 328478 199220
rect 301074 199052 301084 199108
rect 301140 199052 331100 199108
rect 331156 199052 331166 199108
rect 269864 198268 273084 198324
rect 273140 198268 273150 198324
rect 319442 198156 319452 198212
rect 319508 198156 342300 198212
rect 342356 198156 342366 198212
rect 352342 198156 352380 198212
rect 352436 198156 352446 198212
rect 298946 198044 298956 198100
rect 299012 198044 324828 198100
rect 324884 198044 324894 198100
rect 310482 197932 310492 197988
rect 310548 197932 337260 197988
rect 337316 197932 337326 197988
rect 311378 197820 311388 197876
rect 311444 197820 338828 197876
rect 338884 197820 338894 197876
rect 299954 197708 299964 197764
rect 300020 197708 330204 197764
rect 330260 197708 330270 197764
rect 315858 197596 315868 197652
rect 315924 197596 347340 197652
rect 347396 197596 347406 197652
rect 312274 197484 312284 197540
rect 312340 197484 345548 197540
rect 345604 197484 345614 197540
rect 296930 197372 296940 197428
rect 296996 197372 331996 197428
rect 332052 197372 332062 197428
rect 300178 197260 300188 197316
rect 300244 197260 322140 197316
rect 322196 197260 322206 197316
rect 318518 197148 318556 197204
rect 318612 197148 318622 197204
rect 325238 197148 325276 197204
rect 325332 197148 325342 197204
rect 323596 196588 324100 196644
rect 323596 196532 323652 196588
rect 324044 196532 324100 196588
rect 300066 196476 300076 196532
rect 300132 196476 323652 196532
rect 323782 196476 323820 196532
rect 323876 196476 323886 196532
rect 324044 196476 327516 196532
rect 327572 196476 327582 196532
rect 271282 196364 271292 196420
rect 271348 196364 351260 196420
rect 351316 196364 351326 196420
rect 314132 196252 323820 196308
rect 323876 196252 323886 196308
rect 314132 195972 314188 196252
rect 300514 195916 300524 195972
rect 300580 195916 314188 195972
rect 318546 195804 318556 195860
rect 318612 195804 345100 195860
rect 345156 195804 345166 195860
rect 298386 195692 298396 195748
rect 298452 195692 325276 195748
rect 325332 195692 325342 195748
rect 269864 195356 272748 195412
rect 272804 195356 272814 195412
rect 351250 195244 351260 195300
rect 351316 195244 355096 195300
rect 336952 194572 339948 194628
rect 340004 194572 340014 194628
rect 339938 193228 339948 193284
rect 340004 193228 340396 193284
rect 340452 193228 340462 193284
rect 269864 192444 272636 192500
rect 272692 192444 272702 192500
rect 336354 192444 336364 192500
rect 336420 192444 336430 192500
rect -960 192052 480 192248
rect -960 192024 14252 192052
rect 392 191996 14252 192024
rect 14308 191996 14318 192052
rect 336364 191912 336420 192444
rect 595560 192164 597000 192360
rect 590482 192108 590492 192164
rect 590548 192136 597000 192164
rect 590548 192108 595672 192136
rect 269864 189532 272860 189588
rect 272916 189532 272926 189588
rect 336952 189196 340508 189252
rect 340564 189196 340574 189252
rect 345650 189196 345660 189252
rect 345716 189196 354844 189252
rect 354900 189196 355096 189252
rect 269864 186620 272412 186676
rect 272468 186620 272478 186676
rect 336952 186508 340284 186564
rect 340340 186508 340350 186564
rect 336952 183820 351820 183876
rect 351876 183820 351886 183876
rect 269864 183708 273420 183764
rect 273476 183708 273486 183764
rect 354498 183372 354508 183428
rect 354564 183372 355180 183428
rect 355236 183372 355246 183428
rect 351810 183260 351820 183316
rect 351876 183260 354060 183316
rect 354116 183260 354126 183316
rect 340386 183148 340396 183204
rect 340452 183148 355404 183204
rect 355460 183148 355470 183204
rect 349412 181356 352044 181412
rect 352100 181356 352110 181412
rect 336952 181132 349356 181188
rect 349412 181132 349468 181356
rect 269864 180796 272188 180852
rect 272244 180796 272254 180852
rect 585442 179116 585452 179172
rect 585508 179144 595672 179172
rect 585508 179116 597000 179144
rect 595560 178920 597000 179116
rect 336952 178444 352044 178500
rect 352100 178444 352110 178500
rect -960 178052 480 178136
rect -960 177996 4284 178052
rect 4340 177996 4350 178052
rect -960 177912 480 177996
rect 269864 177884 272860 177940
rect 272916 177884 272926 177940
rect 344194 177212 344204 177268
rect 344260 177212 354508 177268
rect 354564 177212 354574 177268
rect 340162 177100 340172 177156
rect 340228 177100 355096 177156
rect 336952 175756 352716 175812
rect 352772 175756 352782 175812
rect 269864 174972 272748 175028
rect 272804 174972 272814 175028
rect 353490 173852 353500 173908
rect 353556 173852 354172 173908
rect 354228 173852 354238 173908
rect 352258 173628 352268 173684
rect 352324 173628 354172 173684
rect 354228 173628 354238 173684
rect 336952 173068 352268 173124
rect 352324 173068 352334 173124
rect 269864 172060 274428 172116
rect 274484 172060 274494 172116
rect 351138 171276 351148 171332
rect 351204 171276 352380 171332
rect 352436 171276 352446 171332
rect 352706 171052 352716 171108
rect 352772 171052 355096 171108
rect 336952 170380 351148 170436
rect 351204 170380 351214 170436
rect 269864 169148 271292 169204
rect 271348 169148 271358 169204
rect 336952 167692 351260 167748
rect 351316 167692 351820 167748
rect 351876 167692 351886 167748
rect 269864 166236 272636 166292
rect 272692 166236 272702 166292
rect 354722 166236 354732 166292
rect 354788 166236 356076 166292
rect 356132 166236 356142 166292
rect 345762 166124 345772 166180
rect 345828 166124 590940 166180
rect 590996 166124 591006 166180
rect 337362 165676 337372 165732
rect 337428 165676 590716 165732
rect 590772 165676 590782 165732
rect 595560 165704 597000 165928
rect 353490 165564 353500 165620
rect 353556 165564 486444 165620
rect 486500 165564 486510 165620
rect 337586 165452 337596 165508
rect 337652 165452 557900 165508
rect 557956 165452 557966 165508
rect 352370 165340 352380 165396
rect 352436 165340 422716 165396
rect 422772 165340 422782 165396
rect 466162 165340 466172 165396
rect 466228 165340 590492 165396
rect 590548 165340 590558 165396
rect 354162 165228 354172 165284
rect 354228 165228 422940 165284
rect 422996 165228 423006 165284
rect 349010 165116 349020 165172
rect 349076 165116 365820 165172
rect 365876 165116 365886 165172
rect 336952 165004 339724 165060
rect 339780 165004 339790 165060
rect 348562 165004 348572 165060
rect 348628 165004 553308 165060
rect 553364 165004 553374 165060
rect 356738 164892 356748 164948
rect 356804 164892 423164 164948
rect 423220 164892 423230 164948
rect 457874 164780 457884 164836
rect 457940 164780 557900 164836
rect 557956 164780 557966 164836
rect 420802 164668 420812 164724
rect 420868 164668 557004 164724
rect 557060 164668 557070 164724
rect 581186 164668 581196 164724
rect 581252 164668 586460 164724
rect 586516 164668 586526 164724
rect 350690 164556 350700 164612
rect 350756 164556 379820 164612
rect 379876 164556 379886 164612
rect 350242 164444 350252 164500
rect 350308 164444 504028 164500
rect 504084 164444 504094 164500
rect 350466 164332 350476 164388
rect 350532 164332 462364 164388
rect 462420 164332 462430 164388
rect 348786 164220 348796 164276
rect 348852 164220 427644 164276
rect 427700 164220 427710 164276
rect 339714 164108 339724 164164
rect 339780 164108 399868 164164
rect 399924 164108 399934 164164
rect 464930 164108 464940 164164
rect 464996 164108 590604 164164
rect 590660 164108 590670 164164
rect -960 163828 480 164024
rect 354274 163996 354284 164052
rect 354340 163996 481068 164052
rect 481124 163996 481134 164052
rect 352034 163884 352044 163940
rect 352100 163884 421820 163940
rect 421876 163884 421886 163940
rect 463586 163884 463596 163940
rect 463652 163884 590828 163940
rect 590884 163884 590894 163940
rect -960 163800 41132 163828
rect 392 163772 41132 163800
rect 41188 163772 41198 163828
rect 342178 163772 342188 163828
rect 342244 163772 553644 163828
rect 553700 163772 553710 163828
rect 345314 163660 345324 163716
rect 345380 163660 517916 163716
rect 517972 163660 517982 163716
rect 269864 163324 273980 163380
rect 274036 163324 274046 163380
rect 462802 163212 462812 163268
rect 462868 163212 495852 163268
rect 495908 163212 495918 163268
rect 460002 163100 460012 163156
rect 460068 163100 553980 163156
rect 554036 163100 554046 163156
rect 457762 162988 457772 163044
rect 457828 162988 556220 163044
rect 556276 162988 556286 163044
rect 348898 162876 348908 162932
rect 348964 162876 358204 162932
rect 358260 162876 358270 162932
rect 476998 162876 477036 162932
rect 477092 162876 477102 162932
rect 497830 162876 497868 162932
rect 497924 162876 497934 162932
rect 532326 162876 532364 162932
rect 532420 162876 532430 162932
rect 539270 162876 539308 162932
rect 539364 162876 539374 162932
rect 546438 162876 546476 162932
rect 546532 162876 546542 162932
rect 339602 162764 339612 162820
rect 339668 162764 448588 162820
rect 448644 162764 448654 162820
rect 567746 162764 567756 162820
rect 567812 162764 584668 162820
rect 584724 162764 584734 162820
rect 341842 162652 341852 162708
rect 341908 162652 441868 162708
rect 441924 162652 441934 162708
rect 574466 162652 574476 162708
rect 574532 162652 586348 162708
rect 586404 162652 586414 162708
rect 350578 162540 350588 162596
rect 350644 162540 435148 162596
rect 435204 162540 435214 162596
rect 560690 162540 560700 162596
rect 560756 162540 584780 162596
rect 584836 162540 584846 162596
rect 336354 162428 336364 162484
rect 336420 162428 336430 162484
rect 349234 162428 349244 162484
rect 349300 162428 372092 162484
rect 372148 162428 372158 162484
rect 458210 162428 458220 162484
rect 458276 162428 469308 162484
rect 469364 162428 469374 162484
rect 336364 162372 336420 162428
rect 336364 162344 352604 162372
rect 336392 162316 352604 162344
rect 352660 162316 502796 162372
rect 502852 162316 502862 162372
rect 342290 162204 342300 162260
rect 342356 162204 554652 162260
rect 554708 162204 554718 162260
rect 293234 162092 293244 162148
rect 293300 162092 520044 162148
rect 520100 162092 520110 162148
rect 348674 161980 348684 162036
rect 348740 161980 490700 162036
rect 490756 161980 490766 162036
rect 462914 161644 462924 161700
rect 462980 161644 497196 161700
rect 497252 161644 497262 161700
rect 460114 161532 460124 161588
rect 460180 161532 554652 161588
rect 554708 161532 554718 161588
rect 460226 161420 460236 161476
rect 460292 161420 556892 161476
rect 556948 161420 556958 161476
rect 457762 161308 457772 161364
rect 457828 161308 555100 161364
rect 555156 161308 555166 161364
rect 355394 161196 355404 161252
rect 355460 161196 483980 161252
rect 484036 161196 484046 161252
rect 341954 161084 341964 161140
rect 342020 161084 414316 161140
rect 414372 161084 414382 161140
rect 346294 160972 346332 161028
rect 346388 160972 346398 161028
rect 353826 160972 353836 161028
rect 353892 160972 393484 161028
rect 393540 160972 393550 161028
rect 304220 160860 314188 160916
rect 300402 160748 300412 160804
rect 300468 160748 303996 160804
rect 304052 160748 304062 160804
rect 304220 160692 304276 160860
rect 284498 160636 284508 160692
rect 284564 160636 304276 160692
rect 314132 160692 314188 160860
rect 314132 160636 516012 160692
rect 516068 160636 516078 160692
rect 300626 160524 300636 160580
rect 300692 160524 304332 160580
rect 304388 160524 304398 160580
rect 307346 160524 307356 160580
rect 307412 160524 540876 160580
rect 540932 160524 540942 160580
rect 269864 160412 271180 160468
rect 271236 160412 271246 160468
rect 300514 160412 300524 160468
rect 300580 160412 302876 160468
rect 302932 160412 302942 160468
rect 303986 160412 303996 160468
rect 304052 160412 550956 160468
rect 551012 160412 551022 160468
rect 283602 160300 283612 160356
rect 283668 160300 514668 160356
rect 514724 160300 514734 160356
rect 281810 160188 281820 160244
rect 281876 160188 508732 160244
rect 508788 160188 508798 160244
rect 291778 160076 291788 160132
rect 291844 160076 513324 160132
rect 513380 160076 513390 160132
rect 458098 159852 458108 159908
rect 458164 159852 479724 159908
rect 479780 159852 479790 159908
rect 480386 159740 480396 159796
rect 480452 159740 558348 159796
rect 558404 159740 558414 159796
rect 457874 159628 457884 159684
rect 457940 159628 556332 159684
rect 556388 159628 556398 159684
rect 346882 159516 346892 159572
rect 346948 159516 347228 159572
rect 347284 159516 347294 159572
rect 354050 159516 354060 159572
rect 354116 159516 422492 159572
rect 422548 159516 422558 159572
rect 298834 159404 298844 159460
rect 298900 159404 522508 159460
rect 522564 159404 522574 159460
rect 299730 159292 299740 159348
rect 299796 159292 532588 159348
rect 532644 159292 532654 159348
rect 300626 159180 300636 159236
rect 300692 159180 535948 159236
rect 536004 159180 536014 159236
rect 302306 159068 302316 159124
rect 302372 159068 539196 159124
rect 539252 159068 539262 159124
rect 298946 158956 298956 159012
rect 299012 158956 544236 159012
rect 544292 158956 544302 159012
rect 297154 158844 297164 158900
rect 297220 158844 542892 158900
rect 542948 158844 542958 158900
rect 297266 158732 297276 158788
rect 297332 158732 548268 158788
rect 548324 158732 548334 158788
rect 345426 158620 345436 158676
rect 345492 158620 386540 158676
rect 386596 158620 386606 158676
rect 460450 158060 460460 158116
rect 460516 158060 482412 158116
rect 482468 158060 482478 158116
rect 457986 157948 457996 158004
rect 458052 157948 554988 158004
rect 555044 157948 555054 158004
rect 306534 157836 306572 157892
rect 306628 157836 306638 157892
rect 322242 157836 322252 157892
rect 322308 157836 341068 157892
rect 341124 157836 341134 157892
rect 346070 157836 346108 157892
rect 346164 157836 346174 157892
rect 349122 157836 349132 157892
rect 349188 157836 468636 157892
rect 468692 157836 468702 157892
rect 470306 157836 470316 157892
rect 470372 157836 583660 157892
rect 583716 157836 583726 157892
rect 300066 157724 300076 157780
rect 300132 157724 311276 157780
rect 311332 157724 311342 157780
rect 333218 157724 333228 157780
rect 333284 157724 343868 157780
rect 343924 157724 554540 157780
rect 554596 157724 554606 157780
rect 301074 157612 301084 157668
rect 301140 157612 317548 157668
rect 317604 157612 317614 157668
rect 334786 157612 334796 157668
rect 334852 157612 343980 157668
rect 344036 157612 555212 157668
rect 555268 157612 555278 157668
rect 269864 157500 272524 157556
rect 272580 157500 272590 157556
rect 298722 157500 298732 157556
rect 298788 157500 314412 157556
rect 314468 157500 314478 157556
rect 326946 157500 326956 157556
rect 327012 157500 344204 157556
rect 344260 157500 556780 157556
rect 556836 157500 556846 157556
rect 298498 157388 298508 157444
rect 298564 157388 312844 157444
rect 312900 157388 312910 157444
rect 328514 157388 328524 157444
rect 328580 157388 346556 157444
rect 346612 157388 559468 157444
rect 559524 157388 559534 157444
rect 296930 157276 296940 157332
rect 296996 157276 319116 157332
rect 319172 157276 319182 157332
rect 331650 157276 331660 157332
rect 331716 157276 342972 157332
rect 343028 157276 556220 157332
rect 556276 157276 556286 157332
rect 299954 157164 299964 157220
rect 300020 157164 315980 157220
rect 316036 157164 316046 157220
rect 323810 157164 323820 157220
rect 323876 157164 337708 157220
rect 342290 157164 342300 157220
rect 342356 157164 556108 157220
rect 556164 157164 556174 157220
rect 337652 157108 337708 157164
rect 298610 157052 298620 157108
rect 298676 157052 320684 157108
rect 320740 157052 320750 157108
rect 337652 157052 339836 157108
rect 339892 157052 342748 157108
rect 342804 157052 342814 157108
rect 349412 157052 559580 157108
rect 559636 157052 559646 157108
rect 349412 156996 349468 157052
rect 298386 156940 298396 156996
rect 298452 156940 308140 156996
rect 308196 156940 308206 156996
rect 330082 156940 330092 156996
rect 330148 156940 344316 156996
rect 344372 156940 349468 156996
rect 356514 156940 356524 156996
rect 356580 156940 422492 156996
rect 422548 156940 422558 156996
rect 473778 156940 473788 156996
rect 473844 156940 583884 156996
rect 583940 156940 583950 156996
rect 300850 156828 300860 156884
rect 300916 156828 309708 156884
rect 309764 156828 309774 156884
rect 325378 156828 325388 156884
rect 325444 156828 341068 156884
rect 341124 156828 342300 156884
rect 342356 156828 342366 156884
rect 460562 156268 460572 156324
rect 460628 156268 474348 156324
rect 474404 156268 474414 156324
rect 353602 156156 353612 156212
rect 353668 156156 525420 156212
rect 525476 156156 525486 156212
rect 346658 156044 346668 156100
rect 346724 156044 460012 156100
rect 460068 156044 460078 156100
rect 291666 155932 291676 155988
rect 291732 155932 510748 155988
rect 510804 155932 510814 155988
rect 288418 155820 288428 155876
rect 288484 155820 510636 155876
rect 510692 155820 510702 155876
rect 294914 155708 294924 155764
rect 294980 155708 525420 155764
rect 525476 155708 525486 155764
rect 292562 155596 292572 155652
rect 292628 155596 528108 155652
rect 528164 155596 528174 155652
rect 293458 155484 293468 155540
rect 293524 155484 529452 155540
rect 529508 155484 529518 155540
rect 297042 155372 297052 155428
rect 297108 155372 534828 155428
rect 534884 155372 534894 155428
rect 355506 155260 355516 155316
rect 355572 155260 366268 155316
rect 366324 155260 366334 155316
rect 460674 154700 460684 154756
rect 460740 154700 473004 154756
rect 473060 154700 473070 154756
rect 269864 154588 274316 154644
rect 274372 154588 274382 154644
rect 459442 154588 459452 154644
rect 459508 154588 556444 154644
rect 556500 154588 556510 154644
rect 335906 154476 335916 154532
rect 335972 154476 339948 154532
rect 340004 154476 340014 154532
rect 345650 154476 345660 154532
rect 345716 154476 421596 154532
rect 421652 154476 421662 154532
rect 468626 154476 468636 154532
rect 468692 154476 478828 154532
rect 483718 154476 483756 154532
rect 483812 154476 483822 154532
rect 487750 154476 487788 154532
rect 487844 154476 487854 154532
rect 488870 154476 488908 154532
rect 488964 154476 488974 154532
rect 489234 154476 489244 154532
rect 489300 154476 490476 154532
rect 490532 154476 490542 154532
rect 491782 154476 491820 154532
rect 491876 154476 491886 154532
rect 493126 154476 493164 154532
rect 493220 154476 493230 154532
rect 502786 154476 502796 154532
rect 502852 154476 506604 154532
rect 506660 154476 506670 154532
rect 508722 154476 508732 154532
rect 508788 154476 511980 154532
rect 512036 154476 512046 154532
rect 532578 154476 532588 154532
rect 532644 154476 538860 154532
rect 538916 154476 538926 154532
rect 478772 154420 478828 154476
rect 273298 154364 273308 154420
rect 273364 154364 274204 154420
rect 274260 154364 351932 154420
rect 351988 154364 352604 154420
rect 352660 154364 352670 154420
rect 423154 154364 423164 154420
rect 423220 154364 467628 154420
rect 467684 154364 467694 154420
rect 478772 154364 497364 154420
rect 535938 154364 535948 154420
rect 536004 154364 540204 154420
rect 540260 154364 540270 154420
rect 497308 154308 497364 154364
rect 345874 154252 345884 154308
rect 345940 154252 420812 154308
rect 420868 154252 420878 154308
rect 422482 154252 422492 154308
rect 422548 154252 463596 154308
rect 463652 154252 463662 154308
rect 497298 154252 497308 154308
rect 497364 154252 497374 154308
rect 539186 154252 539196 154308
rect 539252 154252 541548 154308
rect 541604 154252 541614 154308
rect 273074 154140 273084 154196
rect 273140 154140 274092 154196
rect 274148 154140 337708 154196
rect 422706 154140 422716 154196
rect 422772 154140 464940 154196
rect 464996 154140 465006 154196
rect 337652 153860 337708 154140
rect 422930 154028 422940 154084
rect 422996 154028 466060 154084
rect 466116 154028 466126 154084
rect 500098 154028 500108 154084
rect 500164 154028 524076 154084
rect 524132 154028 524142 154084
rect 421810 153916 421820 153972
rect 421876 153916 468972 153972
rect 469028 153916 470316 153972
rect 470372 153916 470382 153972
rect 471650 153916 471660 153972
rect 471716 153916 581756 153972
rect 581812 153916 581822 153972
rect 337652 153804 352156 153860
rect 352212 153804 501228 153860
rect 501284 153804 501294 153860
rect 522498 153804 522508 153860
rect 522564 153804 537516 153860
rect 537572 153804 537582 153860
rect 352594 153692 352604 153748
rect 352660 153692 502572 153748
rect 502628 153692 502638 153748
rect 510738 153692 510748 153748
rect 510804 153692 526764 153748
rect 526820 153692 526830 153748
rect 540866 153692 540876 153748
rect 540932 153692 549612 153748
rect 549668 153692 549678 153748
rect 272262 153580 272300 153636
rect 272356 153580 272366 153636
rect 497298 153580 497308 153636
rect 497364 153580 509292 153636
rect 509348 153580 509358 153636
rect 340386 153468 340396 153524
rect 340452 153468 505260 153524
rect 505316 153468 505326 153524
rect 507266 153468 507276 153524
rect 507332 153468 536172 153524
rect 536228 153468 536238 153524
rect 500658 153356 500668 153412
rect 500724 153356 522732 153412
rect 522788 153356 522798 153412
rect 494722 153244 494732 153300
rect 494788 153244 518700 153300
rect 518756 153244 518766 153300
rect 520818 153244 520828 153300
rect 520884 153244 530796 153300
rect 530852 153244 530862 153300
rect 463698 153132 463708 153188
rect 463764 153132 558012 153188
rect 558068 153132 558078 153188
rect 352258 153020 352268 153076
rect 352324 153020 503916 153076
rect 503972 153020 503982 153076
rect 525812 153020 533484 153076
rect 533540 153020 533550 153076
rect 525812 152964 525868 153020
rect 470306 152908 470316 152964
rect 470372 152908 473788 152964
rect 473844 152908 473854 152964
rect 475654 152908 475692 152964
rect 475748 152908 475758 152964
rect 485062 152908 485100 152964
rect 485156 152908 485166 152964
rect 494470 152908 494508 152964
rect 494564 152908 494574 152964
rect 498502 152908 498540 152964
rect 498596 152908 498606 152964
rect 499846 152908 499884 152964
rect 499940 152908 499950 152964
rect 505586 152908 505596 152964
rect 505652 152908 521388 152964
rect 521444 152908 521454 152964
rect 524178 152908 524188 152964
rect 524244 152908 525868 152964
rect 527436 152908 532140 152964
rect 532196 152908 532206 152964
rect 527436 152852 527492 152908
rect 295250 152796 295260 152852
rect 295316 152796 527492 152852
rect 557890 152796 557900 152852
rect 557956 152796 558460 152852
rect 558516 152796 558526 152852
rect 280018 152684 280028 152740
rect 280084 152684 497308 152740
rect 497364 152684 497374 152740
rect 590146 152684 590156 152740
rect 590212 152712 595672 152740
rect 590212 152684 597000 152712
rect 288194 152572 288204 152628
rect 288260 152572 505596 152628
rect 505652 152572 505662 152628
rect 350802 152460 350812 152516
rect 350868 152460 352268 152516
rect 352324 152460 352334 152516
rect 595560 152488 597000 152684
rect 337362 152348 337372 152404
rect 337428 152348 558236 152404
rect 558292 152348 558302 152404
rect 279122 152236 279132 152292
rect 279188 152236 507948 152292
rect 508004 152236 508014 152292
rect 285394 152124 285404 152180
rect 285460 152124 517356 152180
rect 517412 152124 517422 152180
rect 303426 152012 303436 152068
rect 303492 152012 545580 152068
rect 545636 152012 545646 152068
rect 269864 151676 277340 151732
rect 277396 151676 277406 151732
rect 334674 151340 334684 151396
rect 334740 151340 340396 151396
rect 340452 151340 340462 151396
rect 461570 151340 461580 151396
rect 461636 151340 471660 151396
rect 471716 151340 471726 151396
rect 330082 151228 330092 151284
rect 330148 151228 350812 151284
rect 350868 151228 350878 151284
rect 463586 151228 463596 151284
rect 463652 151228 478380 151284
rect 478436 151228 478446 151284
rect 342038 151116 342076 151172
rect 342132 151116 342142 151172
rect 350802 151116 350812 151172
rect 350868 151116 352044 151172
rect 352100 151116 352110 151172
rect 557778 151116 557788 151172
rect 557844 151116 558012 151172
rect 558068 151116 558078 151172
rect 294354 151004 294364 151060
rect 294420 151004 520828 151060
rect 520884 151004 520894 151060
rect 288978 150892 288988 150948
rect 289044 150892 500668 150948
rect 500724 150892 500734 150948
rect 297938 150780 297948 150836
rect 298004 150780 507276 150836
rect 507332 150780 507342 150836
rect 342402 150668 342412 150724
rect 342468 150668 511532 150724
rect 511588 150668 511598 150724
rect 345762 150444 345772 150500
rect 345828 150444 461916 150500
rect 461972 150444 461982 150500
rect 342738 150332 342748 150388
rect 342804 150332 554428 150388
rect 554484 150332 554494 150388
rect 296146 150220 296156 150276
rect 296212 150220 524188 150276
rect 524244 150220 524254 150276
rect -960 149716 480 149912
rect 476998 149884 477036 149940
rect 477092 149884 477102 149940
rect 463026 149772 463036 149828
rect 463092 149772 556556 149828
rect 556612 149772 556622 149828
rect -960 149688 24332 149716
rect 392 149660 24332 149688
rect 24388 149660 24398 149716
rect 331762 149660 331772 149716
rect 331828 149660 350812 149716
rect 350868 149660 350878 149716
rect 461682 149660 461692 149716
rect 461748 149660 470316 149716
rect 470372 149660 470382 149716
rect 494694 149660 494732 149716
rect 494788 149660 494798 149716
rect 500070 149660 500108 149716
rect 500164 149660 500174 149716
rect 300514 149548 300524 149604
rect 300580 149548 546924 149604
rect 546980 149548 546990 149604
rect 337138 149436 337148 149492
rect 337204 149436 557788 149492
rect 557844 149436 557854 149492
rect 349010 149324 349020 149380
rect 349076 149324 457884 149380
rect 457940 149324 457950 149380
rect 494498 149324 494508 149380
rect 494564 149324 500108 149380
rect 500164 149324 500174 149380
rect 345090 149212 345100 149268
rect 345156 149212 556668 149268
rect 556724 149212 556734 149268
rect 289874 149100 289884 149156
rect 289940 149100 494508 149156
rect 494564 149100 494574 149156
rect 494722 149100 494732 149156
rect 494788 149100 494798 149156
rect 494732 149044 494788 149100
rect 286290 148988 286300 149044
rect 286356 148988 494788 149044
rect 269864 148764 272412 148820
rect 272468 148764 272478 148820
rect 461906 148764 461916 148820
rect 461972 148764 554092 148820
rect 554148 148764 554158 148820
rect 347330 148652 347340 148708
rect 347396 148652 554876 148708
rect 554932 148652 554942 148708
rect 458546 148316 458556 148372
rect 458612 148316 554764 148372
rect 554820 148316 554830 148372
rect 459340 147924 460040 147980
rect 457650 147868 457660 147924
rect 457716 147868 459396 147924
rect 558114 147868 558124 147924
rect 558180 147868 558236 147924
rect 558292 147868 558302 147924
rect 342514 147756 342524 147812
rect 342580 147756 456988 147812
rect 457044 147756 457054 147812
rect 346994 147644 347004 147700
rect 347060 147644 458220 147700
rect 458276 147644 458286 147700
rect 345202 147532 345212 147588
rect 345268 147532 456092 147588
rect 456148 147532 456158 147588
rect 348898 147420 348908 147476
rect 348964 147420 458444 147476
rect 458500 147420 458510 147476
rect 354050 147308 354060 147364
rect 354116 147308 457660 147364
rect 457716 147308 457726 147364
rect 353714 147196 353724 147252
rect 353780 147196 421372 147252
rect 421428 147196 421438 147252
rect 355282 147084 355292 147140
rect 355348 147084 407484 147140
rect 407540 147084 407550 147140
rect 270162 146972 270172 147028
rect 270228 146972 401884 147028
rect 401940 146972 401950 147028
rect 323362 146188 323372 146244
rect 323428 146188 351036 146244
rect 351092 146188 351932 146244
rect 351988 146188 351998 146244
rect 350802 146076 350812 146132
rect 350868 146076 458108 146132
rect 458164 146076 458174 146132
rect 269836 145460 269892 145880
rect 366230 145852 366268 145908
rect 366324 145852 366334 145908
rect 330866 145516 330876 145572
rect 330932 145516 352380 145572
rect 352436 145516 352446 145572
rect 269836 145404 271292 145460
rect 271348 145404 336364 145460
rect 336420 145404 336430 145460
rect 269266 145292 269276 145348
rect 269332 145292 400316 145348
rect 400372 145292 400382 145348
rect 342290 145068 342300 145124
rect 342356 145068 459396 145124
rect 459340 145012 460040 145068
rect 421810 144620 421820 144676
rect 421876 144620 422492 144676
rect 422548 144620 422558 144676
rect 273186 144508 273196 144564
rect 273252 144508 274652 144564
rect 274708 144508 274718 144564
rect 421670 144508 421708 144564
rect 421764 144508 421774 144564
rect 557778 143836 557788 143892
rect 557844 143836 558236 143892
rect 558292 143836 558302 143892
rect 269836 143612 272300 143668
rect 272356 143612 334684 143668
rect 334740 143612 334750 143668
rect 558114 143612 558124 143668
rect 558180 143612 558190 143668
rect 269836 142968 269892 143612
rect 558124 143556 558180 143612
rect 557890 143500 557900 143556
rect 557956 143500 558180 143556
rect 557778 143388 557788 143444
rect 557844 143388 558124 143444
rect 558180 143388 558190 143444
rect 554904 142940 557900 142996
rect 557956 142940 557966 142996
rect 301634 142716 301644 142772
rect 301700 142716 457212 142772
rect 457268 142716 457278 142772
rect 337250 142604 337260 142660
rect 337316 142604 458556 142660
rect 458612 142604 458622 142660
rect 354722 142156 354732 142212
rect 354788 142156 459396 142212
rect 459340 142100 460040 142156
rect 554904 141372 555212 141428
rect 555268 141372 555278 141428
rect 338370 141036 338380 141092
rect 338436 141036 457996 141092
rect 458052 141036 458062 141092
rect 353714 140924 353724 140980
rect 353780 140924 457772 140980
rect 457828 140924 457838 140980
rect 554530 140476 554540 140532
rect 554596 140476 554606 140532
rect 269836 140252 272412 140308
rect 272468 140252 330876 140308
rect 330932 140252 330942 140308
rect 269836 140056 269892 140252
rect 554540 139832 554596 140476
rect 595560 139412 597000 139496
rect 345538 139356 345548 139412
rect 345604 139356 459452 139412
rect 459508 139356 459518 139412
rect 587346 139356 587356 139412
rect 587412 139356 597000 139412
rect 350466 139244 350476 139300
rect 350532 139244 459396 139300
rect 595560 139272 597000 139356
rect 459340 139188 460040 139244
rect 344082 139132 344092 139188
rect 344148 139132 457884 139188
rect 457940 139132 457950 139188
rect 291554 138572 291564 138628
rect 291620 138572 406588 138628
rect 406644 138572 406654 138628
rect 554904 138236 556220 138292
rect 556276 138236 556286 138292
rect 338818 137676 338828 137732
rect 338884 137676 457772 137732
rect 457828 137676 457838 137732
rect 269864 137116 273308 137172
rect 273364 137116 273374 137172
rect 554904 136668 559580 136724
rect 559636 136668 559646 136724
rect 342178 136332 342188 136388
rect 342244 136332 459396 136388
rect 459340 136276 460040 136332
rect -960 135604 480 135800
rect -960 135576 27692 135604
rect 392 135548 27692 135576
rect 27748 135548 27758 135604
rect 278226 135212 278236 135268
rect 278292 135212 415996 135268
rect 416052 135212 416062 135268
rect 554904 135100 559468 135156
rect 559524 135100 559534 135156
rect 269864 134204 273084 134260
rect 273140 134204 273150 134260
rect 271058 133532 271068 133588
rect 271124 133532 403452 133588
rect 403508 133532 403518 133588
rect 554904 133532 556780 133588
rect 556836 133532 556846 133588
rect 345426 133420 345436 133476
rect 345492 133420 459396 133476
rect 459340 133364 460040 133420
rect 279906 131964 279916 132020
rect 279972 131964 408156 132020
rect 408212 131964 408222 132020
rect 554904 131964 556108 132020
rect 556164 131964 556174 132020
rect 277330 131852 277340 131908
rect 277396 131852 414428 131908
rect 414484 131852 414494 131908
rect 269864 131292 272188 131348
rect 272244 131292 272254 131348
rect 554418 130956 554428 131012
rect 554484 130956 554494 131012
rect 353938 130508 353948 130564
rect 354004 130508 459396 130564
rect 459340 130452 460040 130508
rect 554428 130424 554484 130956
rect 554904 128828 558236 128884
rect 558292 128828 558302 128884
rect 274754 128492 274764 128548
rect 274820 128492 352044 128548
rect 352100 128492 352110 128548
rect 269864 128380 273196 128436
rect 273252 128380 273262 128436
rect 345202 127596 345212 127652
rect 345268 127596 459396 127652
rect 459340 127540 460040 127596
rect 554904 127260 557788 127316
rect 557844 127260 557854 127316
rect 595560 126056 597000 126280
rect 554642 125916 554652 125972
rect 554708 125916 554718 125972
rect 554652 125720 554708 125916
rect 269864 125468 293244 125524
rect 293300 125468 293310 125524
rect 275538 125132 275548 125188
rect 275604 125132 411292 125188
rect 411348 125132 411358 125188
rect 341842 124684 341852 124740
rect 341908 124684 459396 124740
rect 459340 124628 460040 124684
rect 554904 124124 556668 124180
rect 556724 124124 556734 124180
rect 335122 122668 335132 122724
rect 335188 122668 335916 122724
rect 335972 122668 423276 122724
rect 423332 122668 423342 122724
rect 421932 122612 421988 122668
rect 269864 122556 323372 122612
rect 323428 122556 323438 122612
rect 421922 122556 421932 122612
rect 421988 122556 421998 122612
rect 554904 122556 555212 122612
rect 555268 122556 555278 122612
rect 350914 121772 350924 121828
rect 350980 121772 459396 121828
rect 459340 121716 460040 121772
rect -960 121492 480 121688
rect -960 121464 4172 121492
rect 392 121436 4172 121464
rect 4228 121436 4238 121492
rect 554904 120988 556556 121044
rect 556612 120988 556622 121044
rect 554866 120204 554876 120260
rect 554932 120204 554942 120260
rect 269864 119644 311612 119700
rect 311668 119644 311678 119700
rect 554876 119448 554932 120204
rect 339826 118860 339836 118916
rect 339892 118860 459396 118916
rect 459340 118804 460040 118860
rect 554904 117852 556332 117908
rect 556388 117852 556398 117908
rect 554876 116844 555212 116900
rect 555268 116844 555278 116900
rect 269864 116732 347116 116788
rect 347172 116732 347182 116788
rect 554876 116312 554932 116844
rect 459340 115892 460040 115948
rect 340722 115836 340732 115892
rect 340788 115836 459396 115892
rect 276434 115052 276444 115108
rect 276500 115052 412860 115108
rect 412916 115052 412926 115108
rect 554904 114716 556444 114772
rect 556500 114716 556510 114772
rect 269864 113820 337260 113876
rect 337316 113820 337326 113876
rect 554904 113148 555100 113204
rect 555156 113148 555166 113204
rect 345874 113036 345884 113092
rect 345940 113036 459396 113092
rect 590482 113036 590492 113092
rect 590548 113064 595672 113092
rect 590548 113036 597000 113064
rect 459340 112980 460040 113036
rect 595560 112840 597000 113036
rect 554754 112140 554764 112196
rect 554820 112140 554830 112196
rect 554764 111608 554820 112140
rect 269864 110908 272188 110964
rect 272244 110908 272254 110964
rect 350914 110124 350924 110180
rect 350980 110124 459396 110180
rect 459340 110068 460040 110124
rect 355618 110012 355628 110068
rect 355684 110012 458108 110068
rect 458164 110012 458174 110068
rect 554904 110012 556332 110068
rect 556388 110012 556398 110068
rect 554876 108780 554988 108836
rect 555044 108780 555054 108836
rect 554876 108472 554932 108780
rect 269864 107996 272972 108052
rect 273028 107996 273038 108052
rect -960 107380 480 107576
rect -960 107352 31052 107380
rect 392 107324 31052 107352
rect 31108 107324 31118 107380
rect 343634 107324 343644 107380
rect 343700 107324 386092 107380
rect 386148 107324 386158 107380
rect 354386 107212 354396 107268
rect 354452 107212 459396 107268
rect 459340 107156 460040 107212
rect 274866 107100 274876 107156
rect 274932 107100 352156 107156
rect 352212 107100 352222 107156
rect 301186 106988 301196 107044
rect 301252 106988 390796 107044
rect 390852 106988 390862 107044
rect 300962 106876 300972 106932
rect 301028 106876 393932 106932
rect 393988 106876 393998 106932
rect 554904 106876 558236 106932
rect 558292 106876 558302 106932
rect 298162 106764 298172 106820
rect 298228 106764 395500 106820
rect 395556 106764 395566 106820
rect 271954 106652 271964 106708
rect 272020 106652 404908 106708
rect 404964 106652 404974 106708
rect 554904 105308 558124 105364
rect 558180 105308 558190 105364
rect 269864 105084 273420 105140
rect 273476 105084 273486 105140
rect 353826 105084 353836 105140
rect 353892 105084 458220 105140
rect 458276 105084 458286 105140
rect 274642 104972 274652 105028
rect 274708 104972 406588 105028
rect 406644 104972 406654 105028
rect 351026 104300 351036 104356
rect 351092 104300 459396 104356
rect 459340 104244 460040 104300
rect 293122 104076 293132 104132
rect 293188 104076 376572 104132
rect 376628 104076 376638 104132
rect 396498 104076 396508 104132
rect 396564 104076 396602 104132
rect 398150 104076 398188 104132
rect 398244 104076 398254 104132
rect 554306 104076 554316 104132
rect 554372 104076 554410 104132
rect 295026 103964 295036 104020
rect 295092 103964 383964 104020
rect 384020 103964 384030 104020
rect 291442 103852 291452 103908
rect 291508 103852 381388 103908
rect 381444 103852 381454 103908
rect 281362 103740 281372 103796
rect 281428 103740 372988 103796
rect 373044 103740 373054 103796
rect 554904 103740 558012 103796
rect 558068 103740 558078 103796
rect 284834 103628 284844 103684
rect 284900 103628 378028 103684
rect 378084 103628 378094 103684
rect 288306 103516 288316 103572
rect 288372 103516 383180 103572
rect 383236 103516 383246 103572
rect 289650 103404 289660 103460
rect 289716 103404 387100 103460
rect 387156 103404 387166 103460
rect 279794 103292 279804 103348
rect 279860 103292 379708 103348
rect 379764 103292 379774 103348
rect 392326 103292 392364 103348
rect 392420 103292 392430 103348
rect 294802 103180 294812 103236
rect 294868 103180 374668 103236
rect 374724 103180 374734 103236
rect 389190 103180 389228 103236
rect 389284 103180 389294 103236
rect 406578 102508 406588 102564
rect 406644 102508 408940 102564
rect 408996 102508 409006 102564
rect 269864 102172 349132 102228
rect 349188 102172 349198 102228
rect 554306 102172 554316 102228
rect 554372 102172 554382 102228
rect 355506 101612 355516 101668
rect 355572 101612 457884 101668
rect 457940 101612 457950 101668
rect 349346 101388 349356 101444
rect 349412 101388 459396 101444
rect 459340 101332 460040 101388
rect 554306 100604 554316 100660
rect 554372 100604 554382 100660
rect 301522 99932 301532 99988
rect 301588 99932 458556 99988
rect 458612 99932 458622 99988
rect 554306 99932 554316 99988
rect 554372 99932 554410 99988
rect 587122 99820 587132 99876
rect 587188 99848 595672 99876
rect 587188 99820 597000 99848
rect 595560 99624 597000 99820
rect 269864 99260 272972 99316
rect 273028 99260 273038 99316
rect 353910 99036 353948 99092
rect 354004 99036 354014 99092
rect 354834 99036 354844 99092
rect 354900 99036 419356 99092
rect 419412 99036 419422 99092
rect 554904 99036 557900 99092
rect 557956 99036 557966 99092
rect 350690 98924 350700 98980
rect 350756 98924 457996 98980
rect 458052 98924 458062 98980
rect 350242 98812 350252 98868
rect 350308 98812 457436 98868
rect 457492 98812 457502 98868
rect 348562 98700 348572 98756
rect 348628 98700 457660 98756
rect 457716 98700 457726 98756
rect 349234 98588 349244 98644
rect 349300 98588 458332 98644
rect 458388 98588 458398 98644
rect 348786 98476 348796 98532
rect 348852 98476 457772 98532
rect 457828 98476 457838 98532
rect 459340 98420 460040 98476
rect 345538 98364 345548 98420
rect 345604 98364 449372 98420
rect 449428 98364 449438 98420
rect 457650 98364 457660 98420
rect 457716 98364 459396 98420
rect 344306 98252 344316 98308
rect 344372 98252 457324 98308
rect 457380 98252 457390 98308
rect 355394 98140 355404 98196
rect 355460 98140 421708 98196
rect 421764 98140 421774 98196
rect 449362 97804 449372 97860
rect 449428 97804 458444 97860
rect 458500 97804 458510 97860
rect 554904 97468 559132 97524
rect 559188 97468 559198 97524
rect 356626 97244 356636 97300
rect 356692 97244 457548 97300
rect 457604 97244 457614 97300
rect 419346 97020 419356 97076
rect 419412 97020 419422 97076
rect 419356 96628 419412 97020
rect 419356 96572 425852 96628
rect 425908 96572 425918 96628
rect 269266 96348 269276 96404
rect 269332 96348 269342 96404
rect 554904 95900 556220 95956
rect 556276 95900 556286 95956
rect 342486 95676 342524 95732
rect 342580 95676 342590 95732
rect 459340 95508 460040 95564
rect 457650 95452 457660 95508
rect 457716 95452 459396 95508
rect 554306 94332 554316 94388
rect 554372 94332 554382 94388
rect -960 93268 480 93464
rect 269864 93436 366268 93492
rect 366324 93436 366334 93492
rect -960 93240 26012 93268
rect 392 93212 26012 93240
rect 26068 93212 26078 93268
rect 554904 92764 555100 92820
rect 555156 92764 555166 92820
rect 457650 92652 457660 92708
rect 457716 92652 459396 92708
rect 459340 92596 460040 92652
rect 419916 91588 419972 92120
rect 273074 91532 273084 91588
rect 273140 91532 351932 91588
rect 351988 91532 351998 91588
rect 419916 91532 421708 91588
rect 421764 91532 424172 91588
rect 424228 91532 424238 91588
rect 366258 91420 366268 91476
rect 366324 91420 370104 91476
rect 554754 91196 554764 91252
rect 554820 91196 554830 91252
rect 269864 90524 283052 90580
rect 283108 90524 283118 90580
rect 272962 89852 272972 89908
rect 273028 89852 335132 89908
rect 335188 89852 335198 89908
rect 457314 89740 457324 89796
rect 457380 89740 459396 89796
rect 459340 89684 460040 89740
rect 554642 89628 554652 89684
rect 554708 89628 554718 89684
rect 554904 88060 558012 88116
rect 558068 88060 558078 88116
rect 269864 87612 331772 87668
rect 331828 87612 331838 87668
rect 419944 87164 421932 87220
rect 421988 87164 421998 87220
rect 457650 86828 457660 86884
rect 457716 86828 459396 86884
rect 459340 86772 460040 86828
rect 554904 86492 558124 86548
rect 558180 86492 558190 86548
rect 595560 86408 597000 86632
rect 554876 85260 554988 85316
rect 555044 85260 555054 85316
rect 554876 84952 554932 85260
rect 269864 84700 330092 84756
rect 330148 84700 330158 84756
rect 458098 83916 458108 83972
rect 458164 83916 459396 83972
rect 459340 83860 460040 83916
rect 554904 83356 558460 83412
rect 558516 83356 558526 83412
rect 554306 82292 554316 82348
rect 554372 82292 554382 82348
rect 419944 82264 421820 82292
rect 419916 82236 421820 82264
rect 421876 82236 421886 82292
rect 554316 82236 554652 82292
rect 554708 82236 554718 82292
rect 269864 81788 274764 81844
rect 274820 81788 274830 81844
rect 419916 81620 419972 82236
rect 554866 81788 554876 81844
rect 554932 81788 554942 81844
rect 419916 81564 420028 81620
rect 420084 81564 420094 81620
rect 457426 81004 457436 81060
rect 457492 81004 459396 81060
rect 459340 80948 460040 81004
rect 554530 80220 554540 80276
rect 554596 80220 554606 80276
rect -960 79156 480 79352
rect -960 79128 27692 79156
rect 392 79100 27692 79128
rect 27748 79100 27758 79156
rect 269864 78876 273084 78932
rect 273140 78876 273150 78932
rect 554904 78652 558348 78708
rect 558404 78652 558414 78708
rect 458210 78092 458220 78148
rect 458276 78092 459396 78148
rect 459340 78036 460040 78092
rect 419944 77308 420140 77364
rect 420196 77308 421708 77364
rect 421764 77308 421774 77364
rect 554904 77084 556108 77140
rect 556164 77084 556174 77140
rect 269864 75964 274876 76020
rect 274932 75964 274942 76020
rect 554904 75516 557004 75572
rect 557060 75516 557070 75572
rect 458322 75180 458332 75236
rect 458388 75180 459396 75236
rect 459340 75124 460040 75180
rect 337026 74844 337036 74900
rect 337092 74844 370104 74900
rect 554306 73948 554316 74004
rect 554372 73948 554382 74004
rect 595560 73220 597000 73416
rect 590482 73164 590492 73220
rect 590548 73192 597000 73220
rect 590548 73164 595672 73192
rect 269864 73052 272972 73108
rect 273028 73052 273038 73108
rect 419944 72380 420252 72436
rect 420308 72380 422268 72436
rect 422324 72380 422334 72436
rect 554418 72380 554428 72436
rect 554484 72380 554494 72436
rect 459340 72212 460040 72268
rect 458434 72156 458444 72212
rect 458500 72156 459396 72212
rect 554904 70812 556892 70868
rect 556948 70812 556958 70868
rect 269864 70140 272972 70196
rect 273028 70140 273038 70196
rect 457874 69356 457884 69412
rect 457940 69356 459396 69412
rect 459340 69300 460040 69356
rect 554904 69244 557788 69300
rect 557844 69244 557854 69300
rect 421922 68796 421932 68852
rect 421988 68796 423164 68852
rect 423220 68796 423230 68852
rect 554306 67676 554316 67732
rect 554372 67676 554382 67732
rect 419944 67452 421932 67508
rect 421988 67452 421998 67508
rect 269864 67228 273196 67284
rect 273252 67228 273262 67284
rect 457986 66444 457996 66500
rect 458052 66444 459396 66500
rect 459340 66388 460040 66444
rect 425842 66332 425852 66388
rect 425908 66332 457548 66388
rect 457604 66332 457614 66388
rect 554904 66108 558348 66164
rect 558404 66108 558414 66164
rect -960 65044 480 65240
rect -960 65016 29372 65044
rect 392 64988 29372 65016
rect 29428 64988 29438 65044
rect 554904 64540 557788 64596
rect 557844 64540 557854 64596
rect 269864 64316 273084 64372
rect 273140 64316 273150 64372
rect 457762 63532 457772 63588
rect 457828 63532 459396 63588
rect 459340 63476 460040 63532
rect 554904 62972 558124 63028
rect 558180 62972 558190 63028
rect 419944 62524 420364 62580
rect 420420 62524 422940 62580
rect 422996 62524 423006 62580
rect 269864 61404 288204 61460
rect 288260 61404 288270 61460
rect 554904 61404 558236 61460
rect 558292 61404 558302 61460
rect 424162 61292 424172 61348
rect 424228 61292 457660 61348
rect 457716 61292 457726 61348
rect 457538 60620 457548 60676
rect 457604 60620 459396 60676
rect 459340 60564 460040 60620
rect 595560 60004 597000 60200
rect 590594 59948 590604 60004
rect 590660 59976 597000 60004
rect 590660 59948 595672 59976
rect 554904 59836 557900 59892
rect 557956 59836 557966 59892
rect 351138 58716 351148 58772
rect 351204 58716 352716 58772
rect 352772 58716 352782 58772
rect 269864 58492 273756 58548
rect 273812 58492 273822 58548
rect 367826 58268 367836 58324
rect 367892 58268 370104 58324
rect 554904 58268 558012 58324
rect 558068 58268 558078 58324
rect 457650 57708 457660 57764
rect 457716 57708 459396 57764
rect 459340 57652 460040 57708
rect 419944 57596 421708 57652
rect 421764 57596 422716 57652
rect 422772 57596 422782 57652
rect 351138 57148 351148 57204
rect 351204 57148 367836 57204
rect 367892 57148 367902 57204
rect 554428 56084 554484 56728
rect 554418 56028 554428 56084
rect 554484 56028 554494 56084
rect 269864 55580 288988 55636
rect 289044 55580 289054 55636
rect 458546 54796 458556 54852
rect 458612 54796 459396 54852
rect 459340 54740 460040 54796
rect 327506 52892 327516 52948
rect 327572 52892 351148 52948
rect 351204 52892 351214 52948
rect 269864 52668 274204 52724
rect 274260 52668 274270 52724
rect 419384 52696 422492 52724
rect 419356 52668 422492 52696
rect 422548 52668 422558 52724
rect 419356 52164 419412 52668
rect 419346 52108 419356 52164
rect 419412 52108 419422 52164
rect 459340 51828 460040 51884
rect 392 51128 10892 51156
rect -960 51100 10892 51128
rect 10948 51100 10958 51156
rect -960 50904 480 51100
rect 459340 51044 459396 51828
rect 367938 50988 367948 51044
rect 368004 50988 459396 51044
rect 4162 50316 4172 50372
rect 4228 50316 272412 50372
rect 272468 50316 272478 50372
rect 338034 50316 338044 50372
rect 338100 50316 557788 50372
rect 557844 50316 557854 50372
rect 27682 50204 27692 50260
rect 27748 50204 272300 50260
rect 272356 50204 272366 50260
rect 346882 50204 346892 50260
rect 346948 50204 557900 50260
rect 557956 50204 557966 50260
rect 40898 50092 40908 50148
rect 40964 50092 45612 50148
rect 45668 50092 45678 50148
rect 161746 50092 161756 50148
rect 161812 50092 269388 50148
rect 269444 50092 269454 50148
rect 350354 50092 350364 50148
rect 350420 50092 558236 50148
rect 558292 50092 558302 50148
rect 156034 49980 156044 50036
rect 156100 49980 270844 50036
rect 270900 49980 270910 50036
rect 273074 49980 273084 50036
rect 273140 49980 420252 50036
rect 420308 49980 420318 50036
rect 150322 49868 150332 49924
rect 150388 49868 270956 49924
rect 271012 49868 271022 49924
rect 273746 49868 273756 49924
rect 273812 49868 420364 49924
rect 420420 49868 420430 49924
rect 43474 49756 43484 49812
rect 43540 49756 49868 49812
rect 49924 49756 49934 49812
rect 144610 49756 144620 49812
rect 144676 49756 271180 49812
rect 271236 49756 271246 49812
rect 274194 49756 274204 49812
rect 274260 49756 419356 49812
rect 419412 49756 419422 49812
rect 41122 49644 41132 49700
rect 41188 49644 49644 49700
rect 49700 49644 49710 49700
rect 112242 49644 112252 49700
rect 112308 49644 271068 49700
rect 271124 49644 271134 49700
rect 288194 49644 288204 49700
rect 288260 49644 421932 49700
rect 421988 49644 421998 49700
rect 41010 49532 41020 49588
rect 41076 49532 87500 49588
rect 87556 49532 87566 49588
rect 95106 49532 95116 49588
rect 95172 49532 269724 49588
rect 269780 49532 269790 49588
rect 288978 49532 288988 49588
rect 289044 49532 421708 49588
rect 421764 49532 421774 49588
rect 97346 48636 97356 48692
rect 97412 48636 293580 48692
rect 293636 48636 327516 48692
rect 327572 48636 327582 48692
rect 336914 48636 336924 48692
rect 336980 48636 590604 48692
rect 590660 48636 590670 48692
rect 201730 48524 201740 48580
rect 201796 48524 266924 48580
rect 266980 48524 266990 48580
rect 290098 48524 290108 48580
rect 290164 48524 322252 48580
rect 322308 48524 322318 48580
rect 340946 48524 340956 48580
rect 341012 48524 557788 48580
rect 557844 48524 557854 48580
rect 203634 48412 203644 48468
rect 203700 48412 269724 48468
rect 269780 48412 269790 48468
rect 290322 48412 290332 48468
rect 290388 48412 315084 48468
rect 315140 48412 315150 48468
rect 342626 48412 342636 48468
rect 342692 48412 558124 48468
rect 558180 48412 558190 48468
rect 196018 48300 196028 48356
rect 196084 48300 276220 48356
rect 276276 48300 276286 48356
rect 290546 48300 290556 48356
rect 290612 48300 307916 48356
rect 307972 48300 307982 48356
rect 345986 48300 345996 48356
rect 346052 48300 558012 48356
rect 558068 48300 558078 48356
rect 40674 48188 40684 48244
rect 40740 48188 53228 48244
rect 53284 48188 53294 48244
rect 138898 48188 138908 48244
rect 138964 48188 270732 48244
rect 270788 48188 270798 48244
rect 286402 48188 286412 48244
rect 286468 48188 300748 48244
rect 300804 48188 300814 48244
rect 345986 48188 345996 48244
rect 346052 48188 558348 48244
rect 558404 48188 558414 48244
rect 43362 48076 43372 48132
rect 43428 48076 77980 48132
rect 78036 48076 78046 48132
rect 133186 48076 133196 48132
rect 133252 48076 269388 48132
rect 269444 48076 269454 48132
rect 272962 48076 272972 48132
rect 273028 48076 420028 48132
rect 420084 48076 420094 48132
rect 40786 47964 40796 48020
rect 40852 47964 81788 48020
rect 81844 47964 81854 48020
rect 127474 47964 127484 48020
rect 127540 47964 269500 48020
rect 269556 47964 269566 48020
rect 273186 47964 273196 48020
rect 273252 47964 420140 48020
rect 420196 47964 420206 48020
rect 46946 47852 46956 47908
rect 47012 47852 97356 47908
rect 97412 47852 97422 47908
rect 121762 47852 121772 47908
rect 121828 47852 269612 47908
rect 269668 47852 269678 47908
rect 212258 47740 212268 47796
rect 212324 47740 267596 47796
rect 267652 47740 267662 47796
rect 46946 47068 46956 47124
rect 47012 47068 47022 47124
rect 46956 47012 47012 47068
rect 40226 46956 40236 47012
rect 40292 46956 45388 47012
rect 45444 46956 47012 47012
rect 595560 46760 597000 46984
rect 199938 46508 199948 46564
rect 200004 46508 339500 46564
rect 339556 46508 339566 46564
rect 131282 46396 131292 46452
rect 131348 46396 337148 46452
rect 337204 46396 337214 46452
rect 125570 46284 125580 46340
rect 125636 46284 338604 46340
rect 338660 46284 338670 46340
rect 62738 46172 62748 46228
rect 62804 46172 336924 46228
rect 336980 46172 336990 46228
rect 190306 45276 190316 45332
rect 190372 45276 275884 45332
rect 275940 45276 275950 45332
rect 286514 45276 286524 45332
rect 286580 45276 590492 45332
rect 590548 45276 590558 45332
rect 184594 45164 184604 45220
rect 184660 45164 275996 45220
rect 276052 45164 276062 45220
rect 355170 45164 355180 45220
rect 355236 45164 554428 45220
rect 554484 45164 554494 45220
rect 178882 45052 178892 45108
rect 178948 45052 275772 45108
rect 275828 45052 275838 45108
rect 173170 44940 173180 44996
rect 173236 44940 270620 44996
rect 270676 44940 270686 44996
rect 167458 44828 167468 44884
rect 167524 44828 269500 44884
rect 269556 44828 269566 44884
rect 152226 44716 152236 44772
rect 152292 44716 277228 44772
rect 277284 44716 277294 44772
rect 106530 44604 106540 44660
rect 106596 44604 270956 44660
rect 271012 44604 271022 44660
rect 100818 44492 100828 44548
rect 100884 44492 269948 44548
rect 270004 44492 270014 44548
rect 207442 44380 207452 44436
rect 207508 44380 276108 44436
rect 276164 44380 276174 44436
rect 175074 43372 175084 43428
rect 175140 43372 280588 43428
rect 280644 43372 280654 43428
rect 176978 43260 176988 43316
rect 177044 43260 339388 43316
rect 339444 43260 339454 43316
rect 142818 43148 142828 43204
rect 142884 43148 338940 43204
rect 338996 43148 339006 43204
rect 119858 43036 119868 43092
rect 119924 43036 338828 43092
rect 338884 43036 338894 43092
rect 114258 42924 114268 42980
rect 114324 42924 338604 42980
rect 338660 42924 338670 42980
rect 68450 42812 68460 42868
rect 68516 42812 338716 42868
rect 338772 42812 338782 42868
rect 129378 41916 129388 41972
rect 129444 41916 270732 41972
rect 270788 41916 270798 41972
rect 192322 41804 192332 41860
rect 192388 41804 336812 41860
rect 336868 41804 336878 41860
rect 123666 41692 123676 41748
rect 123732 41692 270620 41748
rect 270676 41692 270686 41748
rect 117954 41580 117964 41636
rect 118020 41580 270844 41636
rect 270900 41580 270910 41636
rect 108434 41468 108444 41524
rect 108500 41468 338940 41524
rect 338996 41468 339006 41524
rect 91298 41356 91308 41412
rect 91364 41356 343756 41412
rect 343812 41356 343822 41412
rect 85698 41244 85708 41300
rect 85764 41244 338492 41300
rect 338548 41244 338558 41300
rect 79874 41132 79884 41188
rect 79940 41132 343532 41188
rect 343588 41132 343598 41188
rect 180786 41020 180796 41076
rect 180852 41020 274092 41076
rect 274148 41020 274158 41076
rect 197922 39452 197932 39508
rect 197988 39452 275660 39508
rect 275716 39452 275726 39508
rect 140802 38220 140812 38276
rect 140868 38220 267372 38276
rect 267428 38220 267438 38276
rect 146514 38108 146524 38164
rect 146580 38108 275548 38164
rect 275604 38108 275614 38164
rect 188402 37996 188412 38052
rect 188468 37996 338492 38052
rect 338548 37996 338558 38052
rect 182690 37884 182700 37940
rect 182756 37884 339052 37940
rect 339108 37884 339118 37940
rect 83682 37772 83692 37828
rect 83748 37772 273868 37828
rect 273924 37772 273934 37828
rect -960 36820 480 37016
rect -960 36792 271292 36820
rect 392 36764 271292 36792
rect 271348 36764 271358 36820
rect 595560 33684 597000 33768
rect 289762 33628 289772 33684
rect 289828 33628 597000 33684
rect 595560 33544 597000 33628
rect 209346 31164 209356 31220
rect 209412 31164 269612 31220
rect 269668 31164 269678 31220
rect 186498 31052 186508 31108
rect 186564 31052 273980 31108
rect 274036 31052 274046 31108
rect 169362 29372 169372 29428
rect 169428 29372 270508 29428
rect 270564 29372 270574 29428
rect 392 22904 4172 22932
rect -960 22876 4172 22904
rect 4228 22876 4238 22932
rect -960 22680 480 22876
rect 592162 20524 592172 20580
rect 592228 20552 595672 20580
rect 592228 20524 597000 20552
rect 595560 20328 597000 20524
rect 3714 14140 3724 14196
rect 3780 14140 7532 14196
rect 7588 14140 7598 14196
rect 192210 12572 192220 12628
rect 192276 12572 270508 12628
rect 270564 12572 270574 12628
rect 392 8792 3724 8820
rect -960 8764 3724 8792
rect 3780 8764 3790 8820
rect -960 8568 480 8764
rect 163874 7532 163884 7588
rect 163940 7532 278908 7588
rect 278964 7532 278974 7588
rect 595560 7140 597000 7336
rect 276322 7084 276332 7140
rect 276388 7112 597000 7140
rect 276388 7084 595672 7112
rect 11554 5852 11564 5908
rect 11620 5852 45388 5908
rect 45444 5852 45454 5908
rect 158162 5852 158172 5908
rect 158228 5852 269836 5908
rect 269892 5852 269902 5908
rect 40114 4956 40124 5012
rect 40180 4956 60844 5012
rect 60900 4956 60910 5012
rect 205762 4956 205772 5012
rect 205828 4956 284732 5012
rect 284788 4956 284798 5012
rect 580850 4956 580860 5012
rect 580916 4956 584668 5012
rect 584724 4956 584734 5012
rect 40002 4844 40012 4900
rect 40068 4844 64652 4900
rect 64708 4844 64718 4900
rect 97234 4844 97244 4900
rect 97300 4844 192332 4900
rect 192388 4844 192398 4900
rect 194338 4844 194348 4900
rect 194404 4844 289996 4900
rect 290052 4844 290062 4900
rect 40898 4732 40908 4788
rect 40964 4732 66556 4788
rect 66612 4732 66622 4788
rect 165778 4732 165788 4788
rect 165844 4732 279692 4788
rect 279748 4732 279758 4788
rect 35186 4620 35196 4676
rect 35252 4620 42028 4676
rect 42084 4620 42094 4676
rect 43586 4620 43596 4676
rect 43652 4620 76076 4676
rect 76132 4620 76142 4676
rect 171490 4620 171500 4676
rect 171556 4620 288092 4676
rect 288148 4620 288158 4676
rect 39778 4508 39788 4564
rect 39844 4508 72268 4564
rect 72324 4508 72334 4564
rect 160066 4508 160076 4564
rect 160132 4508 289772 4564
rect 289828 4508 289838 4564
rect 36866 4396 36876 4452
rect 36932 4396 70364 4452
rect 70420 4396 70430 4452
rect 135314 4396 135324 4452
rect 135380 4396 273868 4452
rect 273924 4396 273934 4452
rect 38546 4284 38556 4340
rect 38612 4284 47516 4340
rect 47572 4284 47582 4340
rect 49634 4284 49644 4340
rect 49700 4284 93212 4340
rect 93268 4284 93278 4340
rect 116274 4284 116284 4340
rect 116340 4284 267260 4340
rect 267316 4284 267326 4340
rect 336802 4284 336812 4340
rect 336868 4284 582540 4340
rect 582596 4284 582606 4340
rect 15362 4172 15372 4228
rect 15428 4172 16716 4228
rect 16772 4172 16782 4228
rect 17266 4172 17276 4228
rect 17332 4172 18396 4228
rect 18452 4172 18462 4228
rect 21074 4172 21084 4228
rect 21140 4172 21756 4228
rect 21812 4172 21822 4228
rect 26758 4172 26796 4228
rect 26852 4172 26862 4228
rect 32498 4172 32508 4228
rect 32564 4172 33404 4228
rect 33460 4172 33470 4228
rect 41010 4172 41020 4228
rect 41076 4172 41804 4228
rect 41860 4172 41870 4228
rect 42018 4172 42028 4228
rect 42084 4172 49420 4228
rect 49476 4172 49486 4228
rect 49858 4172 49868 4228
rect 49924 4172 98924 4228
rect 98980 4172 98990 4228
rect 102946 4172 102956 4228
rect 103012 4172 104076 4228
rect 104132 4172 104142 4228
rect 110758 4172 110796 4228
rect 110852 4172 110862 4228
rect 114212 4172 267148 4228
rect 267204 4172 267214 4228
rect 284946 4172 284956 4228
rect 285012 4172 584444 4228
rect 584500 4172 584510 4228
rect 114212 4116 114268 4172
rect 38434 4060 38444 4116
rect 38500 4060 58940 4116
rect 58996 4060 59006 4116
rect 74386 4060 74396 4116
rect 74452 4060 75516 4116
rect 75572 4060 75582 4116
rect 89618 4060 89628 4116
rect 89684 4060 90636 4116
rect 90692 4060 90702 4116
rect 104850 4060 104860 4116
rect 104916 4060 114268 4116
rect 154438 4060 154476 4116
rect 154532 4060 154542 4116
rect 211474 4060 211484 4116
rect 211540 4060 278012 4116
rect 278068 4060 278078 4116
rect 55094 3388 55132 3444
rect 55188 3388 55198 3444
rect 57110 3388 57148 3444
rect 57204 3388 57214 3444
rect 137190 3388 137228 3444
rect 137284 3388 137294 3444
rect 148614 3388 148652 3444
rect 148708 3388 148718 3444
<< via3 >>
rect 201516 591276 201572 591332
rect 203196 591164 203252 591220
rect 208124 591052 208180 591108
rect 204652 590940 204708 590996
rect 208012 590828 208068 590884
rect 206332 590716 206388 590772
rect 208236 590604 208292 590660
rect 444332 590156 444388 590212
rect 584668 590156 584724 590212
rect 590492 588588 590548 588644
rect 157052 587132 157108 587188
rect 181356 573692 181412 573748
rect 590492 573692 590548 573748
rect 209468 568652 209524 568708
rect 183036 567868 183092 567924
rect 590604 567868 590660 567924
rect 187964 565068 188020 565124
rect 532924 565068 532980 565124
rect 590492 562156 590548 562212
rect 535948 560364 536004 560420
rect 4172 558908 4228 558964
rect 532700 555660 532756 555716
rect 537628 550956 537684 551012
rect 186396 550732 186452 550788
rect 590604 549164 590660 549220
rect 7532 544796 7588 544852
rect 187852 536396 187908 536452
rect 543452 535724 543508 535780
rect 590716 522508 590772 522564
rect 189532 522060 189588 522116
rect 4284 516572 4340 516628
rect 187740 514892 187796 514948
rect 590604 509292 590660 509348
rect 183932 500556 183988 500612
rect 541772 496076 541828 496132
rect 534268 475692 534324 475748
rect 4172 474236 4228 474292
rect 187068 471884 187124 471940
rect 4172 471212 4228 471268
rect 178892 471212 178948 471268
rect 590828 469644 590884 469700
rect 150332 469532 150388 469588
rect 4172 467852 4228 467908
rect 172172 467852 172228 467908
rect 4284 466172 4340 466228
rect 175532 466172 175588 466228
rect 187292 450380 187348 450436
rect 187404 443212 187460 443268
rect 532812 442764 532868 442820
rect 187628 436044 187684 436100
rect 167132 431900 167188 431956
rect 590940 430108 590996 430164
rect 168812 428876 168868 428932
rect 529228 428652 529284 428708
rect 189420 421708 189476 421764
rect 4172 417788 4228 417844
rect 540092 416780 540148 416836
rect 61852 413308 61908 413364
rect 355404 410060 355460 410116
rect 83916 409724 83972 409780
rect 444332 409388 444388 409444
rect 289772 409164 289828 409220
rect 295596 408940 295652 408996
rect 356748 408492 356804 408548
rect 466956 408492 467012 408548
rect 356524 408156 356580 408212
rect 208012 408044 208068 408100
rect 300636 408044 300692 408100
rect 352492 408044 352548 408100
rect 209468 407820 209524 407876
rect 208124 407708 208180 407764
rect 444892 407820 444948 407876
rect 496412 407596 496468 407652
rect 352604 407484 352660 407540
rect 522172 407484 522228 407540
rect 527324 407484 527380 407540
rect 356076 407372 356132 407428
rect 356412 407372 356468 407428
rect 357756 407148 357812 407204
rect 206668 406700 206724 406756
rect 490588 406700 490644 406756
rect 229964 406588 230020 406644
rect 280476 406588 280532 406644
rect 295596 406588 295652 406644
rect 352492 406588 352548 406644
rect 354396 406588 354452 406644
rect 581756 406588 581812 406644
rect 446012 406364 446068 406420
rect 92428 404908 92484 404964
rect 89964 403228 90020 403284
rect 355516 401548 355572 401604
rect 89852 400316 89908 400372
rect 208236 399084 208292 399140
rect 86492 397404 86548 397460
rect 546252 396844 546308 396900
rect 574028 396844 574084 396900
rect 580972 396732 581028 396788
rect 553196 396620 553252 396676
rect 567084 396508 567140 396564
rect 203196 395836 203252 395892
rect 201516 395724 201572 395780
rect 354956 395164 355012 395220
rect 355292 395164 355348 395220
rect 361228 395164 361284 395220
rect 356636 395052 356692 395108
rect 365148 395052 365204 395108
rect 379820 395052 379876 395108
rect 525532 394940 525588 394996
rect 476924 394716 476980 394772
rect 511644 394716 511700 394772
rect 463036 394604 463092 394660
rect 463708 394604 463764 394660
rect 590716 394604 590772 394660
rect 511644 394380 511700 394436
rect 476924 394156 476980 394212
rect 463036 394044 463092 394100
rect 361228 393820 361284 393876
rect 365148 393820 365204 393876
rect 364476 393260 364532 393316
rect 393148 393260 393204 393316
rect 393148 393036 393204 393092
rect 463708 393036 463764 393092
rect 206332 392812 206388 392868
rect 379820 392812 379876 392868
rect 466956 392812 467012 392868
rect 204652 392700 204708 392756
rect 189420 392476 189476 392532
rect 342860 392476 342916 392532
rect 355180 391356 355236 391412
rect 355292 391244 355348 391300
rect 355404 390796 355460 390852
rect 591164 390572 591220 390628
rect 355068 390460 355124 390516
rect 4284 389564 4340 389620
rect 355628 389452 355684 389508
rect 353612 387660 353668 387716
rect 353836 387548 353892 387604
rect 235116 385980 235172 386036
rect 354956 385980 355012 386036
rect 100156 385196 100212 385252
rect 352044 384972 352100 385028
rect 238364 384860 238420 384916
rect 241836 384524 241892 384580
rect 238476 384412 238532 384468
rect 238588 384300 238644 384356
rect 348572 384188 348628 384244
rect 237804 383068 237860 383124
rect 355516 382956 355572 383012
rect 288092 382732 288148 382788
rect 291452 382732 291508 382788
rect 203196 382508 203252 382564
rect 204764 382508 204820 382564
rect 206556 382508 206612 382564
rect 209916 382508 209972 382564
rect 201404 382396 201460 382452
rect 203084 382396 203140 382452
rect 204876 382396 204932 382452
rect 206444 382396 206500 382452
rect 208124 382396 208180 382452
rect 209804 382396 209860 382452
rect 226716 382060 226772 382116
rect 301532 382060 301588 382116
rect 250236 381948 250292 382004
rect 260316 381948 260372 382004
rect 267036 381948 267092 382004
rect 281708 381948 281764 382004
rect 288876 381948 288932 382004
rect 290556 381948 290612 382004
rect 293916 381948 293972 382004
rect 312396 381948 312452 382004
rect 314076 381948 314132 382004
rect 315756 381948 315812 382004
rect 322588 381948 322644 382004
rect 232764 381388 232820 381444
rect 241500 381388 241556 381444
rect 240156 380828 240212 380884
rect 237692 380716 237748 380772
rect 170492 380604 170548 380660
rect 241724 380604 241780 380660
rect 201292 379708 201348 379764
rect 202860 379708 202916 379764
rect 315756 379708 315812 379764
rect 214172 379596 214228 379652
rect 214396 379596 214452 379652
rect 222012 379484 222068 379540
rect 224028 379484 224084 379540
rect 227612 379484 227668 379540
rect 230076 379484 230132 379540
rect 235452 379484 235508 379540
rect 225148 379260 225204 379316
rect 225820 379260 225876 379316
rect 227836 379260 227892 379316
rect 232540 379260 232596 379316
rect 214172 379148 214228 379204
rect 214396 379036 214452 379092
rect 4172 375676 4228 375732
rect 343196 373996 343252 374052
rect 344092 373100 344148 373156
rect 344204 371308 344260 371364
rect 340620 369516 340676 369572
rect 346892 368620 346948 368676
rect 190652 368060 190708 368116
rect 355292 367724 355348 367780
rect 190652 366940 190708 366996
rect 190652 366380 190708 366436
rect 352268 366156 352324 366212
rect 190652 364588 190708 364644
rect 352268 364588 352324 364644
rect 339500 363244 339556 363300
rect 186508 363020 186564 363076
rect 186620 361900 186676 361956
rect 91532 361228 91588 361284
rect 179788 360780 179844 360836
rect 353612 360556 353668 360612
rect 186508 359772 186564 359828
rect 186396 359660 186452 359716
rect 89964 358652 90020 358708
rect 93324 358652 93380 358708
rect 168924 358540 168980 358596
rect 186620 356412 186676 356468
rect 179788 352940 179844 352996
rect 591052 350924 591108 350980
rect 186396 349580 186452 349636
rect 4396 347228 4452 347284
rect 339276 347116 339332 347172
rect 352716 346444 352772 346500
rect 342860 344428 342916 344484
rect 351932 340396 351988 340452
rect 168028 339500 168084 339556
rect 590828 337596 590884 337652
rect 168140 336812 168196 336868
rect 346780 335468 346836 335524
rect 346556 334572 346612 334628
rect 350028 334348 350084 334404
rect 348684 333676 348740 333732
rect 168252 332780 168308 332836
rect 346108 332780 346164 332836
rect 346668 331884 346724 331940
rect 345548 330988 345604 331044
rect 168700 330876 168756 330932
rect 168364 329420 168420 329476
rect 168700 329420 168756 329476
rect 340060 329308 340116 329364
rect 353724 329196 353780 329252
rect 344988 328300 345044 328356
rect 355068 328300 355124 328356
rect 348908 327404 348964 327460
rect 342076 326508 342132 326564
rect 168924 326060 168980 326116
rect 341964 325612 342020 325668
rect 345324 324716 345380 324772
rect 350588 323820 350644 323876
rect 350364 322924 350420 322980
rect 354396 322252 354452 322308
rect 165900 322028 165956 322084
rect 349020 322028 349076 322084
rect 165900 321692 165956 321748
rect 341068 321132 341124 321188
rect 342412 320908 342468 320964
rect 354396 320908 354452 320964
rect 184492 320460 184548 320516
rect 344092 320236 344148 320292
rect 190652 319340 190708 319396
rect 341180 319340 341236 319396
rect 349132 318444 349188 318500
rect 344876 317548 344932 317604
rect 182812 317100 182868 317156
rect 339388 316988 339444 317044
rect 344652 316652 344708 316708
rect 181244 315980 181300 316036
rect 344540 315756 344596 315812
rect 186396 314860 186452 314916
rect 341292 313964 341348 314020
rect 177996 313740 178052 313796
rect 4284 313292 4340 313348
rect 168924 313292 168980 313348
rect 350812 313068 350868 313124
rect 179676 312620 179732 312676
rect 344764 312172 344820 312228
rect 184380 311500 184436 311556
rect 340396 311276 340452 311332
rect 590716 311276 590772 311332
rect 190428 310380 190484 310436
rect 341404 310380 341460 310436
rect 339276 309484 339332 309540
rect 181020 309260 181076 309316
rect 189532 308140 189588 308196
rect 344428 307692 344484 307748
rect 181132 307020 181188 307076
rect 354508 306796 354564 306852
rect 182700 305900 182756 305956
rect 354060 305900 354116 305956
rect 342300 305004 342356 305060
rect 165452 304892 165508 304948
rect 186172 304780 186228 304836
rect 354732 304220 354788 304276
rect 354844 304108 354900 304164
rect 187740 303660 187796 303716
rect 350476 303212 350532 303268
rect 187964 302540 188020 302596
rect 342188 302316 342244 302372
rect 177884 301420 177940 301476
rect 345436 301420 345492 301476
rect 353948 300524 354004 300580
rect 187180 300300 187236 300356
rect 345212 299628 345268 299684
rect 187516 299180 187572 299236
rect 344428 299068 344484 299124
rect 341404 298956 341460 299012
rect 341852 298732 341908 298788
rect 179564 298060 179620 298116
rect 339388 298060 339444 298116
rect 590604 298060 590660 298116
rect 351148 297836 351204 297892
rect 186956 296940 187012 296996
rect 339836 296940 339892 296996
rect 4396 296492 4452 296548
rect 177212 296492 177268 296548
rect 187068 296492 187124 296548
rect 340732 296044 340788 296100
rect 187852 295820 187908 295876
rect 339948 295596 340004 295652
rect 348012 295148 348068 295204
rect 186060 294700 186116 294756
rect 349580 294252 349636 294308
rect 60396 293916 60452 293972
rect 353388 293132 353444 293188
rect 190652 293020 190708 293076
rect 7532 292460 7588 292516
rect 71820 292348 71876 292404
rect 84588 292348 84644 292404
rect 349468 292348 349524 292404
rect 352044 292012 352100 292068
rect 355180 292012 355236 292068
rect 339612 291564 339668 291620
rect 347788 291564 347844 291620
rect 352828 291452 352884 291508
rect 10892 291340 10948 291396
rect 4284 291004 4340 291060
rect 26012 290556 26068 290612
rect 4284 290444 4340 290500
rect 92316 290444 92372 290500
rect 188076 289884 188132 289940
rect 342748 289772 342804 289828
rect 349692 289772 349748 289828
rect 27692 289100 27748 289156
rect 93996 288876 94052 288932
rect 339724 288876 339780 288932
rect 348572 288876 348628 288932
rect 188076 288092 188132 288148
rect 115052 287980 115108 288036
rect 187068 287308 187124 287364
rect 344316 287084 344372 287140
rect 173852 286860 173908 286916
rect 188076 286524 188132 286580
rect 93996 286412 94052 286468
rect 166348 286412 166404 286468
rect 187068 286412 187124 286468
rect 339276 286188 339332 286244
rect 92316 285740 92372 285796
rect 353500 285964 353556 286020
rect 182252 285628 182308 285684
rect 183932 285628 183988 285684
rect 355628 285628 355684 285684
rect 93996 285404 94052 285460
rect 168028 285404 168084 285460
rect 167468 285292 167524 285348
rect 188076 284732 188132 284788
rect 353388 284732 353444 284788
rect 165452 284620 165508 284676
rect 344764 283836 344820 283892
rect 177212 283500 177268 283556
rect 347900 283500 347956 283556
rect 344764 282604 344820 282660
rect 168924 282380 168980 282436
rect 185724 282156 185780 282212
rect 187292 282156 187348 282212
rect 344876 282156 344932 282212
rect 187068 282044 187124 282100
rect 182252 281932 182308 281988
rect 339724 281708 339780 281764
rect 355516 281708 355572 281764
rect 167132 281260 167188 281316
rect 344204 280812 344260 280868
rect 188076 280588 188132 280644
rect 167468 280476 167524 280532
rect 168140 280476 168196 280532
rect 185612 280476 185668 280532
rect 187628 280476 187684 280532
rect 341292 280476 341348 280532
rect 346108 280476 346164 280532
rect 93996 280364 94052 280420
rect 185948 280364 186004 280420
rect 187404 280364 187460 280420
rect 178892 280140 178948 280196
rect 341404 279916 341460 279972
rect 185948 279132 186004 279188
rect 175532 279020 175588 279076
rect 346220 279020 346276 279076
rect 168140 278908 168196 278964
rect 353836 278908 353892 278964
rect 172172 277900 172228 277956
rect 339948 277452 340004 277508
rect 341180 277228 341236 277284
rect 93996 276108 94052 276164
rect 351260 275436 351316 275492
rect 348012 272972 348068 273028
rect 174636 272076 174692 272132
rect 93996 271852 94052 271908
rect 590716 271404 590772 271460
rect 177996 269836 178052 269892
rect 339276 269164 339332 269220
rect 185724 268716 185780 268772
rect 352044 268716 352100 268772
rect 166348 268604 166404 268660
rect 166348 267820 166404 267876
rect 352044 267820 352100 267876
rect 181356 266700 181412 266756
rect 343084 266476 343140 266532
rect 168140 265804 168196 265860
rect 183036 265580 183092 265636
rect 342860 265580 342916 265636
rect 168028 265356 168084 265412
rect 185612 265356 185668 265412
rect 182924 264460 182980 264516
rect 168028 263788 168084 263844
rect 184604 263340 184660 263396
rect 4284 262780 4340 262836
rect 344652 262332 344708 262388
rect 186284 262220 186340 262276
rect 344092 262108 344148 262164
rect 345100 262108 345156 262164
rect 342972 261996 343028 262052
rect 168812 261772 168868 261828
rect 352268 261772 352324 261828
rect 351260 261212 351316 261268
rect 184716 261100 184772 261156
rect 339612 261100 339668 261156
rect 187068 259980 187124 260036
rect 190652 259756 190708 259812
rect 92428 259084 92484 259140
rect 339276 259308 339332 259364
rect 344540 258636 344596 258692
rect 339276 258412 339332 258468
rect 590492 258412 590548 258468
rect 187628 257740 187684 257796
rect 339276 257516 339332 257572
rect 342636 256956 342692 257012
rect 344988 256956 345044 257012
rect 345996 256956 346052 257012
rect 351820 256956 351876 257012
rect 352492 256956 352548 257012
rect 339388 256844 339444 256900
rect 340060 256844 340116 256900
rect 339388 256620 339444 256676
rect 341068 256172 341124 256228
rect 190652 255724 190708 255780
rect 187404 255500 187460 255556
rect 93324 254828 93380 254884
rect 187292 254380 187348 254436
rect 339388 253708 339444 253764
rect 340060 253708 340116 253764
rect 344428 253036 344484 253092
rect 345100 252924 345156 252980
rect 354172 252924 354228 252980
rect 345548 252700 345604 252756
rect 350140 252700 350196 252756
rect 190652 252364 190708 252420
rect 340172 252028 340228 252084
rect 349580 252028 349636 252084
rect 352828 252028 352884 252084
rect 344652 251244 344708 251300
rect 93660 250572 93716 250628
rect 340060 250012 340116 250068
rect 352604 249676 352660 249732
rect 349468 249452 349524 249508
rect 343196 248556 343252 248612
rect 339388 247884 339444 247940
rect 349692 247772 349748 247828
rect 339276 247660 339332 247716
rect 340396 246988 340452 247044
rect 342524 246988 342580 247044
rect 341292 246876 341348 246932
rect 347788 246876 347844 246932
rect 339276 246764 339332 246820
rect 350252 246764 350308 246820
rect 344540 246652 344596 246708
rect 350700 246652 350756 246708
rect 340284 246540 340340 246596
rect 348460 246540 348516 246596
rect 93436 246316 93492 246372
rect 346108 245868 346164 245924
rect 339388 245308 339444 245364
rect 344652 245196 344708 245252
rect 345884 245196 345940 245252
rect 351820 245196 351876 245252
rect 352492 245196 352548 245252
rect 339388 245084 339444 245140
rect 339388 244860 339444 244916
rect 341404 243628 341460 243684
rect 348796 243628 348852 243684
rect 352492 243628 352548 243684
rect 93436 241948 93492 242004
rect 339388 241948 339444 242004
rect 339948 241948 340004 242004
rect 340956 241948 341012 242004
rect 342524 241948 342580 242004
rect 80444 240940 80500 240996
rect 80444 240716 80500 240772
rect 339724 240604 339780 240660
rect 347900 240604 347956 240660
rect 232764 240492 232820 240548
rect 236124 240492 236180 240548
rect 347900 240268 347956 240324
rect 349244 240268 349300 240324
rect 339724 240156 339780 240212
rect 339948 240156 340004 240212
rect 340844 240156 340900 240212
rect 185948 239932 186004 239988
rect 341404 239932 341460 239988
rect 238476 239820 238532 239876
rect 241836 239708 241892 239764
rect 281372 239708 281428 239764
rect 187180 239596 187236 239652
rect 273980 239596 274036 239652
rect 343084 239596 343140 239652
rect 179564 239484 179620 239540
rect 272972 239484 273028 239540
rect 342636 239484 342692 239540
rect 230972 239372 231028 239428
rect 236796 239260 236852 239316
rect 185724 239148 185780 239204
rect 344540 239148 344596 239204
rect 288316 239036 288372 239092
rect 342972 239036 343028 239092
rect 344428 238700 344484 238756
rect 62636 238476 62692 238532
rect 64428 238476 64484 238532
rect 244188 238476 244244 238532
rect 245084 238476 245140 238532
rect 340060 238476 340116 238532
rect 270508 238252 270564 238308
rect 39676 237916 39732 237972
rect 236796 237020 236852 237076
rect 243404 237020 243460 237076
rect 268716 237020 268772 237076
rect 209916 236908 209972 236964
rect 225148 236908 225204 236964
rect 233436 236908 233492 236964
rect 236684 236908 236740 236964
rect 238476 236908 238532 236964
rect 240044 236908 240100 236964
rect 241836 236908 241892 236964
rect 243516 236908 243572 236964
rect 267036 236908 267092 236964
rect 268604 236908 268660 236964
rect 302316 236908 302372 236964
rect 303436 236908 303492 236964
rect 307356 236908 307412 236964
rect 309036 236908 309092 236964
rect 310716 236908 310772 236964
rect 319116 236908 319172 236964
rect 334236 236908 334292 236964
rect 335916 236908 335972 236964
rect 168812 236796 168868 236852
rect 339388 236796 339444 236852
rect 339948 236796 340004 236852
rect 354284 236796 354340 236852
rect 182252 236684 182308 236740
rect 185612 236572 185668 236628
rect 345660 236572 345716 236628
rect 352940 236572 352996 236628
rect 355404 236572 355460 236628
rect 239484 236460 239540 236516
rect 236012 236348 236068 236404
rect 236236 236236 236292 236292
rect 343196 236124 343252 236180
rect 33516 236012 33572 236068
rect 241500 235116 241556 235172
rect 240156 235004 240212 235060
rect 43484 234556 43540 234612
rect 241724 234556 241780 234612
rect 283052 234556 283108 234612
rect 266924 234444 266980 234500
rect 12572 234332 12628 234388
rect 239932 234332 239988 234388
rect 344316 234332 344372 234388
rect 270060 234220 270116 234276
rect 235228 233436 235284 233492
rect 270620 232876 270676 232932
rect 271068 232764 271124 232820
rect 339276 232652 339332 232708
rect 590940 231868 590996 231924
rect 267260 231756 267316 231812
rect 269500 231644 269556 231700
rect 267484 231532 267540 231588
rect 351820 231532 351876 231588
rect 269612 231420 269668 231476
rect 269388 230860 269444 230916
rect 43596 229516 43652 229572
rect 43372 225932 43428 225988
rect 190428 224924 190484 224980
rect 272860 224924 272916 224980
rect 187292 223020 187348 223076
rect 296604 223020 296660 223076
rect 217644 222684 217700 222740
rect 301532 222684 301588 222740
rect 4284 222572 4340 222628
rect 173852 222572 173908 222628
rect 187740 221340 187796 221396
rect 274428 221340 274484 221396
rect 41020 220892 41076 220948
rect 338380 220892 338436 220948
rect 4284 220444 4340 220500
rect 239372 219884 239428 219940
rect 301644 219884 301700 219940
rect 214284 219772 214340 219828
rect 187516 219660 187572 219716
rect 271180 219660 271236 219716
rect 187404 219212 187460 219268
rect 337036 219212 337092 219268
rect 592284 218764 592340 218820
rect 184380 218092 184436 218148
rect 272524 218092 272580 218148
rect 239708 216412 239764 216468
rect 274652 216412 274708 216468
rect 214172 216300 214228 216356
rect 210812 216188 210868 216244
rect 177884 216076 177940 216132
rect 272636 216076 272692 216132
rect 35196 215852 35252 215908
rect 181020 214844 181076 214900
rect 272300 214844 272356 214900
rect 203196 214620 203252 214676
rect 187628 214508 187684 214564
rect 337372 214508 337428 214564
rect 40908 214396 40964 214452
rect 228172 214172 228228 214228
rect 355404 213388 355460 213444
rect 217532 213164 217588 213220
rect 201404 213052 201460 213108
rect 276332 213052 276388 213108
rect 186060 212940 186116 212996
rect 272412 212940 272468 212996
rect 187852 212828 187908 212884
rect 277340 212828 277396 212884
rect 230076 212716 230132 212772
rect 227612 212604 227668 212660
rect 187964 211372 188020 211428
rect 271292 211372 271348 211428
rect 186172 211260 186228 211316
rect 272188 211260 272244 211316
rect 272412 211260 272468 211316
rect 186956 211148 187012 211204
rect 274316 211148 274372 211204
rect 181244 211036 181300 211092
rect 272748 211036 272804 211092
rect 182812 210924 182868 210980
rect 4284 210812 4340 210868
rect 115052 210812 115108 210868
rect 179676 210812 179732 210868
rect 296492 210700 296548 210756
rect 273196 210476 273252 210532
rect 264796 210028 264852 210084
rect 189532 209804 189588 209860
rect 272972 209804 273028 209860
rect 186396 209692 186452 209748
rect 182700 209580 182756 209636
rect 269276 209580 269332 209636
rect 272188 209580 272244 209636
rect 273420 209580 273476 209636
rect 181132 209468 181188 209524
rect 272636 209468 272692 209524
rect 177996 209356 178052 209412
rect 273084 209356 273140 209412
rect 264796 209020 264852 209076
rect 293132 209020 293188 209076
rect 41132 206108 41188 206164
rect 272748 204092 272804 204148
rect 272860 202524 272916 202580
rect 273196 202524 273252 202580
rect 272188 202412 272244 202468
rect 269276 201180 269332 201236
rect 339164 201180 339220 201236
rect 344204 200956 344260 201012
rect 272972 199836 273028 199892
rect 300636 199276 300692 199332
rect 273084 198268 273140 198324
rect 352380 198156 352436 198212
rect 298956 198044 299012 198100
rect 318556 197148 318612 197204
rect 325276 197148 325332 197204
rect 323820 196476 323876 196532
rect 323820 196252 323876 196308
rect 300524 195916 300580 195972
rect 318556 195804 318612 195860
rect 325276 195692 325332 195748
rect 272748 195356 272804 195412
rect 339948 194572 340004 194628
rect 339948 193228 340004 193284
rect 340396 193228 340452 193284
rect 272636 192444 272692 192500
rect 336364 192444 336420 192500
rect 590492 192108 590548 192164
rect 272860 189532 272916 189588
rect 345660 189196 345716 189252
rect 354844 189196 354900 189252
rect 272412 186620 272468 186676
rect 351820 183820 351876 183876
rect 273420 183708 273476 183764
rect 354508 183372 354564 183428
rect 351820 183260 351876 183316
rect 340396 183148 340452 183204
rect 355404 183148 355460 183204
rect 349356 181132 349412 181188
rect 585452 179116 585508 179172
rect 4284 177996 4340 178052
rect 274428 172060 274484 172116
rect 271292 169148 271348 169204
rect 351820 167692 351876 167748
rect 356076 166236 356132 166292
rect 345772 166124 345828 166180
rect 590940 166124 590996 166180
rect 337372 165676 337428 165732
rect 590716 165676 590772 165732
rect 339724 165004 339780 165060
rect 356748 164892 356804 164948
rect 457884 164780 457940 164836
rect 557900 164780 557956 164836
rect 586460 164668 586516 164724
rect 41132 163772 41188 163828
rect 553644 163772 553700 163828
rect 273980 163324 274036 163380
rect 462812 163212 462868 163268
rect 460012 163100 460068 163156
rect 553980 163100 554036 163156
rect 457772 162988 457828 163044
rect 556220 162988 556276 163044
rect 477036 162876 477092 162932
rect 497868 162876 497924 162932
rect 532364 162876 532420 162932
rect 539308 162876 539364 162932
rect 546476 162876 546532 162932
rect 586348 162652 586404 162708
rect 584780 162540 584836 162596
rect 462924 161644 462980 161700
rect 460124 161532 460180 161588
rect 554652 161532 554708 161588
rect 460236 161420 460292 161476
rect 346332 160972 346388 161028
rect 303996 160748 304052 160804
rect 300636 160524 300692 160580
rect 307356 160524 307412 160580
rect 271180 160412 271236 160468
rect 300524 160412 300580 160468
rect 303996 160412 304052 160468
rect 480396 159740 480452 159796
rect 346892 159516 346948 159572
rect 422492 159516 422548 159572
rect 302316 159068 302372 159124
rect 460460 158060 460516 158116
rect 306572 157836 306628 157892
rect 341068 157836 341124 157892
rect 346108 157836 346164 157892
rect 349132 157836 349188 157892
rect 468636 157836 468692 157892
rect 356524 156940 356580 156996
rect 460572 156268 460628 156324
rect 346668 156044 346724 156100
rect 460012 156044 460068 156100
rect 460684 154700 460740 154756
rect 274316 154588 274372 154644
rect 421596 154476 421652 154532
rect 468636 154476 468692 154532
rect 483756 154476 483812 154532
rect 487788 154476 487844 154532
rect 488908 154476 488964 154532
rect 489244 154476 489300 154532
rect 491820 154476 491876 154532
rect 493164 154476 493220 154532
rect 274204 154364 274260 154420
rect 497308 154252 497364 154308
rect 274092 154140 274148 154196
rect 581756 153916 581812 153972
rect 352156 153804 352212 153860
rect 272300 153580 272356 153636
rect 463708 153132 463764 153188
rect 558012 153132 558068 153188
rect 475692 152908 475748 152964
rect 485100 152908 485156 152964
rect 494508 152908 494564 152964
rect 498540 152908 498596 152964
rect 499884 152908 499940 152964
rect 557900 152796 557956 152852
rect 590156 152684 590212 152740
rect 350812 152460 350868 152516
rect 352268 152460 352324 152516
rect 303436 152012 303492 152068
rect 277340 151676 277396 151732
rect 461580 151340 461636 151396
rect 350812 151228 350868 151284
rect 463596 151228 463652 151284
rect 342076 151116 342132 151172
rect 352044 151116 352100 151172
rect 557788 151116 557844 151172
rect 461916 150444 461972 150500
rect 477036 149884 477092 149940
rect 463036 149772 463092 149828
rect 461692 149660 461748 149716
rect 494732 149660 494788 149716
rect 500108 149660 500164 149716
rect 349020 149324 349076 149380
rect 457884 149324 457940 149380
rect 494508 149324 494564 149380
rect 500108 149324 500164 149380
rect 494508 149100 494564 149156
rect 494732 149100 494788 149156
rect 461916 148764 461972 148820
rect 554092 148764 554148 148820
rect 457660 147868 457716 147924
rect 558236 147868 558292 147924
rect 342524 147756 342580 147812
rect 456988 147756 457044 147812
rect 348908 147420 348964 147476
rect 458444 147420 458500 147476
rect 354060 147308 354116 147364
rect 457660 147308 457716 147364
rect 351036 146188 351092 146244
rect 351932 146188 351988 146244
rect 366268 145852 366324 145908
rect 342300 145068 342356 145124
rect 422492 144620 422548 144676
rect 274652 144508 274708 144564
rect 421708 144508 421764 144564
rect 557788 143836 557844 143892
rect 558236 143836 558292 143892
rect 558124 143612 558180 143668
rect 557900 143500 557956 143556
rect 557788 143388 557844 143444
rect 558124 143388 558180 143444
rect 301644 142716 301700 142772
rect 457212 142716 457268 142772
rect 354732 142156 354788 142212
rect 338380 141036 338436 141092
rect 353724 140924 353780 140980
rect 457772 140924 457828 140980
rect 587356 139356 587412 139412
rect 350476 139244 350532 139300
rect 344092 139132 344148 139188
rect 342188 136332 342244 136388
rect 27692 135548 27748 135604
rect 345436 133420 345492 133476
rect 353948 130508 354004 130564
rect 352044 128492 352100 128548
rect 345212 127596 345268 127652
rect 293244 125468 293300 125524
rect 341852 124684 341908 124740
rect 423276 122668 423332 122724
rect 555212 122556 555268 122612
rect 350924 121772 350980 121828
rect 311612 119644 311668 119700
rect 339836 118860 339892 118916
rect 556332 117852 556388 117908
rect 555212 116844 555268 116900
rect 340732 115836 340788 115892
rect 337260 113820 337316 113876
rect 345884 113036 345940 113092
rect 590492 113036 590548 113092
rect 272188 110908 272244 110964
rect 355628 110012 355684 110068
rect 458108 110012 458164 110068
rect 272972 107996 273028 108052
rect 31052 107324 31108 107380
rect 352156 107100 352212 107156
rect 558236 106876 558292 106932
rect 298172 106764 298228 106820
rect 558124 105308 558180 105364
rect 353836 105084 353892 105140
rect 458220 105084 458276 105140
rect 396508 104076 396564 104132
rect 398188 104076 398244 104132
rect 554316 104076 554372 104132
rect 558012 103740 558068 103796
rect 392364 103292 392420 103348
rect 389228 103180 389284 103236
rect 554316 102172 554372 102228
rect 355516 101612 355572 101668
rect 457884 101612 457940 101668
rect 554316 100604 554372 100660
rect 301532 99932 301588 99988
rect 554316 99932 554372 99988
rect 587132 99820 587188 99876
rect 353948 99036 354004 99092
rect 354844 99036 354900 99092
rect 419356 99036 419412 99092
rect 557900 99036 557956 99092
rect 350700 98924 350756 98980
rect 457996 98924 458052 98980
rect 350252 98812 350308 98868
rect 457436 98812 457492 98868
rect 348572 98700 348628 98756
rect 349244 98588 349300 98644
rect 458332 98588 458388 98644
rect 348796 98476 348852 98532
rect 457772 98476 457828 98532
rect 345548 98364 345604 98420
rect 457660 98364 457716 98420
rect 344316 98252 344372 98308
rect 457324 98252 457380 98308
rect 355404 98140 355460 98196
rect 421708 98140 421764 98196
rect 559132 97468 559188 97524
rect 356636 97244 356692 97300
rect 457548 97244 457604 97300
rect 419356 97020 419412 97076
rect 425852 96572 425908 96628
rect 269276 96348 269332 96404
rect 556220 95900 556276 95956
rect 342524 95676 342580 95732
rect 457660 95452 457716 95508
rect 554316 94332 554372 94388
rect 26012 93212 26068 93268
rect 555100 92764 555156 92820
rect 351932 91532 351988 91588
rect 421708 91532 421764 91588
rect 424172 91532 424228 91588
rect 554764 91196 554820 91252
rect 457324 89740 457380 89796
rect 554652 89628 554708 89684
rect 457660 86828 457716 86884
rect 554988 85260 555044 85316
rect 458108 83916 458164 83972
rect 554316 82292 554372 82348
rect 554652 82236 554708 82292
rect 554876 81788 554932 81844
rect 457436 81004 457492 81060
rect 554540 80220 554596 80276
rect 458220 78092 458276 78148
rect 556108 77084 556164 77140
rect 458332 75180 458388 75236
rect 554316 73948 554372 74004
rect 554428 72380 554484 72436
rect 457884 69356 457940 69412
rect 554316 67676 554372 67732
rect 457996 66444 458052 66500
rect 425852 66332 425908 66388
rect 457548 66332 457604 66388
rect 29372 64988 29428 65044
rect 557788 64540 557844 64596
rect 457772 63532 457828 63588
rect 424172 61292 424228 61348
rect 457660 61292 457716 61348
rect 457548 60620 457604 60676
rect 457660 57708 457716 57764
rect 10892 51100 10948 51156
rect 338044 50316 338100 50372
rect 43484 49756 43540 49812
rect 271068 49644 271124 49700
rect 269724 49532 269780 49588
rect 266924 48524 266980 48580
rect 340956 48524 341012 48580
rect 557788 48524 557844 48580
rect 345996 48300 346052 48356
rect 43372 48076 43428 48132
rect 269388 48076 269444 48132
rect 269500 47964 269556 48020
rect 269612 47852 269668 47908
rect 267596 47740 267652 47796
rect 337148 46396 337204 46452
rect 336924 46172 336980 46228
rect 277228 44716 277284 44772
rect 270956 44604 271012 44660
rect 269948 44492 270004 44548
rect 338828 43036 338884 43092
rect 338604 42924 338660 42980
rect 270732 41916 270788 41972
rect 336812 41804 336868 41860
rect 270620 41692 270676 41748
rect 270844 41580 270900 41636
rect 338940 41468 338996 41524
rect 267372 38220 267428 38276
rect 275548 38108 275604 38164
rect 338492 37996 338548 38052
rect 339052 37884 339108 37940
rect 273868 37772 273924 37828
rect 270508 29372 270564 29428
rect 4172 22876 4228 22932
rect 592172 20524 592228 20580
rect 3724 14140 3780 14196
rect 7532 14140 7588 14196
rect 3724 8764 3780 8820
rect 276332 7084 276388 7140
rect 269836 5852 269892 5908
rect 584668 4956 584724 5012
rect 40908 4732 40964 4788
rect 43596 4620 43652 4676
rect 289772 4508 289828 4564
rect 267260 4284 267316 4340
rect 16716 4172 16772 4228
rect 18396 4172 18452 4228
rect 21756 4172 21812 4228
rect 26796 4172 26852 4228
rect 33404 4172 33460 4228
rect 41020 4172 41076 4228
rect 104076 4172 104132 4228
rect 110796 4172 110852 4228
rect 267148 4172 267204 4228
rect 75516 4060 75572 4116
rect 90636 4060 90692 4116
rect 154476 4060 154532 4116
rect 55132 3388 55188 3444
rect 57148 3388 57204 3444
rect 137228 3388 137284 3444
rect 148652 3388 148708 3444
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 5418 562350 6038 579922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect 4172 558964 4228 558974
rect 4172 478828 4228 558908
rect 5418 544350 6038 561922
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 568350 9758 585922
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect 4060 478772 4228 478828
rect 4284 516628 4340 516638
rect 4060 470998 4116 478772
rect 4172 474292 4228 474302
rect 4172 471268 4228 474236
rect 4172 471202 4228 471212
rect 4060 470942 4228 470998
rect 4172 467908 4228 470942
rect 4172 467842 4228 467852
rect 4284 466228 4340 516572
rect 4284 466162 4340 466172
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 5418 472350 6038 489922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect 5418 454350 6038 471922
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect 4172 417844 4228 417854
rect 4172 416818 4228 417788
rect 4172 416752 4228 416762
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect 5418 400350 6038 417922
rect 7532 544852 7588 544862
rect 7532 409078 7588 544796
rect 7532 409012 7588 409022
rect 9138 532350 9758 549922
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 9138 478350 9758 495922
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect 4284 389620 4340 389630
rect 4172 377218 4228 377228
rect 4060 377162 4172 377218
rect 4060 372988 4116 377162
rect 4172 377152 4228 377162
rect 4172 376318 4228 376328
rect 4172 375732 4228 376262
rect 4172 375666 4228 375676
rect 4060 372932 4228 372988
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect 4172 22932 4228 372932
rect 4284 313348 4340 389564
rect 5418 382350 6038 399922
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 5418 364350 6038 381922
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect 4284 313282 4340 313292
rect 4396 347284 4452 347294
rect 4396 296548 4452 347228
rect 4396 296482 4452 296492
rect 5418 346350 6038 363922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect 5418 328350 6038 345922
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect 4284 294778 4340 294788
rect 4284 291060 4340 294722
rect 4284 290994 4340 291004
rect 5418 292350 6038 309922
rect 9138 406350 9758 423922
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 9138 370350 9758 387922
rect 36138 597212 36758 598268
rect 36138 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 36758 597212
rect 36138 597088 36758 597156
rect 36138 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 36758 597088
rect 36138 596964 36758 597032
rect 36138 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 36758 596964
rect 36138 596840 36758 596908
rect 36138 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 36758 596840
rect 36138 580350 36758 596784
rect 36138 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 36758 580350
rect 36138 580226 36758 580294
rect 36138 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 36758 580226
rect 36138 580102 36758 580170
rect 36138 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 36758 580102
rect 36138 579978 36758 580046
rect 36138 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 36758 579978
rect 36138 562350 36758 579922
rect 36138 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 36758 562350
rect 36138 562226 36758 562294
rect 36138 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 36758 562226
rect 36138 562102 36758 562170
rect 36138 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 36758 562102
rect 36138 561978 36758 562046
rect 36138 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 36758 561978
rect 36138 544350 36758 561922
rect 36138 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 36758 544350
rect 36138 544226 36758 544294
rect 36138 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 36758 544226
rect 36138 544102 36758 544170
rect 36138 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 36758 544102
rect 36138 543978 36758 544046
rect 36138 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 36758 543978
rect 36138 526350 36758 543922
rect 36138 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 36758 526350
rect 36138 526226 36758 526294
rect 36138 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 36758 526226
rect 36138 526102 36758 526170
rect 36138 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 36758 526102
rect 36138 525978 36758 526046
rect 36138 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 36758 525978
rect 36138 508350 36758 525922
rect 36138 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 36758 508350
rect 36138 508226 36758 508294
rect 36138 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 36758 508226
rect 36138 508102 36758 508170
rect 36138 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 36758 508102
rect 36138 507978 36758 508046
rect 36138 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 36758 507978
rect 36138 490350 36758 507922
rect 36138 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 36758 490350
rect 36138 490226 36758 490294
rect 36138 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 36758 490226
rect 36138 490102 36758 490170
rect 36138 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 36758 490102
rect 36138 489978 36758 490046
rect 36138 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 36758 489978
rect 36138 472350 36758 489922
rect 36138 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 36758 472350
rect 36138 472226 36758 472294
rect 36138 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 36758 472226
rect 36138 472102 36758 472170
rect 36138 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 36758 472102
rect 36138 471978 36758 472046
rect 36138 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 36758 471978
rect 36138 454350 36758 471922
rect 36138 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 36758 454350
rect 36138 454226 36758 454294
rect 36138 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 36758 454226
rect 36138 454102 36758 454170
rect 36138 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 36758 454102
rect 36138 453978 36758 454046
rect 36138 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 36758 453978
rect 36138 436350 36758 453922
rect 36138 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 36758 436350
rect 36138 436226 36758 436294
rect 36138 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 36758 436226
rect 36138 436102 36758 436170
rect 36138 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 36758 436102
rect 36138 435978 36758 436046
rect 36138 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 36758 435978
rect 36138 418350 36758 435922
rect 36138 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 36758 418350
rect 36138 418226 36758 418294
rect 36138 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 36758 418226
rect 36138 418102 36758 418170
rect 36138 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 36758 418102
rect 36138 417978 36758 418046
rect 36138 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 36758 417978
rect 36138 400350 36758 417922
rect 36138 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 36758 400350
rect 36138 400226 36758 400294
rect 36138 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 36758 400226
rect 36138 400102 36758 400170
rect 36138 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 36758 400102
rect 36138 399978 36758 400046
rect 36138 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 36758 399978
rect 36138 382350 36758 399922
rect 36138 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 36758 382350
rect 36138 382226 36758 382294
rect 36138 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 36758 382226
rect 36138 382102 36758 382170
rect 36138 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 36758 382102
rect 36138 381978 36758 382046
rect 36138 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 36758 381978
rect 31052 378838 31108 378848
rect 29372 377398 29428 377408
rect 9138 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 9758 370350
rect 9138 370226 9758 370294
rect 9138 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 9758 370226
rect 9138 370102 9758 370170
rect 9138 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 9758 370102
rect 9138 369978 9758 370046
rect 9138 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 9758 369978
rect 9138 352350 9758 369922
rect 9138 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 9758 352350
rect 9138 352226 9758 352294
rect 9138 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 9758 352226
rect 9138 352102 9758 352170
rect 9138 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 9758 352102
rect 9138 351978 9758 352046
rect 9138 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 9758 351978
rect 9138 334350 9758 351922
rect 9138 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 9758 334350
rect 9138 334226 9758 334294
rect 9138 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 9758 334226
rect 9138 334102 9758 334170
rect 9138 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 9758 334102
rect 9138 333978 9758 334046
rect 9138 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 9758 333978
rect 9138 316350 9758 333922
rect 9138 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 9758 316350
rect 9138 316226 9758 316294
rect 9138 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 9758 316226
rect 9138 316102 9758 316170
rect 9138 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 9758 316102
rect 9138 315978 9758 316046
rect 9138 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 9758 315978
rect 9138 298350 9758 315922
rect 9138 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 9758 298350
rect 9138 298226 9758 298294
rect 9138 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 9758 298226
rect 9138 298102 9758 298170
rect 9138 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 9758 298102
rect 9138 297978 9758 298046
rect 9138 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 9758 297978
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 4284 290500 4340 290510
rect 4284 262836 4340 290444
rect 4284 262770 4340 262780
rect 5418 274350 6038 291922
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect 5418 256350 6038 273922
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 4284 222628 4340 222638
rect 4284 220500 4340 222572
rect 4284 220434 4340 220444
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 4284 210868 4340 210878
rect 4284 178052 4340 210812
rect 4284 177986 4340 177996
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 4172 22866 4228 22876
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 5418 148350 6038 165922
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect 3724 14196 3780 14206
rect 3724 8820 3780 14140
rect 3724 8754 3780 8764
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 4350 6038 21922
rect 7532 292516 7588 292526
rect 7532 14196 7588 292460
rect 7532 14130 7588 14140
rect 9138 280350 9758 297922
rect 12572 372178 12628 372188
rect 9138 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 9758 280350
rect 9138 280226 9758 280294
rect 9138 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 9758 280226
rect 9138 280102 9758 280170
rect 9138 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 9758 280102
rect 9138 279978 9758 280046
rect 9138 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 9758 279978
rect 9138 262350 9758 279922
rect 9138 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 9758 262350
rect 9138 262226 9758 262294
rect 9138 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 9758 262226
rect 9138 262102 9758 262170
rect 9138 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 9758 262102
rect 9138 261978 9758 262046
rect 9138 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 9758 261978
rect 9138 244350 9758 261922
rect 9138 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 9758 244350
rect 9138 244226 9758 244294
rect 9138 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 9758 244226
rect 9138 244102 9758 244170
rect 9138 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 9758 244102
rect 9138 243978 9758 244046
rect 9138 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 9758 243978
rect 9138 226350 9758 243922
rect 9138 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 9758 226350
rect 9138 226226 9758 226294
rect 9138 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 9758 226226
rect 9138 226102 9758 226170
rect 9138 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 9758 226102
rect 9138 225978 9758 226046
rect 9138 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 9758 225978
rect 9138 208350 9758 225922
rect 9138 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 9758 208350
rect 9138 208226 9758 208294
rect 9138 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 9758 208226
rect 9138 208102 9758 208170
rect 9138 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 9758 208102
rect 9138 207978 9758 208046
rect 9138 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 9758 207978
rect 9138 190350 9758 207922
rect 9138 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 9758 190350
rect 9138 190226 9758 190294
rect 9138 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 9758 190226
rect 9138 190102 9758 190170
rect 9138 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 9758 190102
rect 9138 189978 9758 190046
rect 9138 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 9758 189978
rect 9138 172350 9758 189922
rect 9138 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 9758 172350
rect 9138 172226 9758 172294
rect 9138 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 9758 172226
rect 9138 172102 9758 172170
rect 9138 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 9758 172102
rect 9138 171978 9758 172046
rect 9138 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 9758 171978
rect 9138 154350 9758 171922
rect 9138 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 9758 154350
rect 9138 154226 9758 154294
rect 9138 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 9758 154226
rect 9138 154102 9758 154170
rect 9138 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 9758 154102
rect 9138 153978 9758 154046
rect 9138 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 9758 153978
rect 9138 136350 9758 153922
rect 9138 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 9758 136350
rect 9138 136226 9758 136294
rect 9138 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 9758 136226
rect 9138 136102 9758 136170
rect 9138 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 9758 136102
rect 9138 135978 9758 136046
rect 9138 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 9758 135978
rect 9138 118350 9758 135922
rect 9138 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 9758 118350
rect 9138 118226 9758 118294
rect 9138 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 9758 118226
rect 9138 118102 9758 118170
rect 9138 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 9758 118102
rect 9138 117978 9758 118046
rect 9138 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 9758 117978
rect 9138 100350 9758 117922
rect 9138 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 9758 100350
rect 9138 100226 9758 100294
rect 9138 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 9758 100226
rect 9138 100102 9758 100170
rect 9138 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 9758 100102
rect 9138 99978 9758 100046
rect 9138 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 9758 99978
rect 9138 82350 9758 99922
rect 9138 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 9758 82350
rect 9138 82226 9758 82294
rect 9138 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 9758 82226
rect 9138 82102 9758 82170
rect 9138 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 9758 82102
rect 9138 81978 9758 82046
rect 9138 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 9758 81978
rect 9138 64350 9758 81922
rect 9138 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 9758 64350
rect 9138 64226 9758 64294
rect 9138 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 9758 64226
rect 9138 64102 9758 64170
rect 9138 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 9758 64102
rect 9138 63978 9758 64046
rect 9138 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 9758 63978
rect 9138 46350 9758 63922
rect 10892 291396 10948 291406
rect 10892 51156 10948 291340
rect 12572 234388 12628 372122
rect 26012 290612 26068 290622
rect 18396 238978 18452 238988
rect 12572 234322 12628 234332
rect 16716 238798 16772 238808
rect 10892 51090 10948 51100
rect 9138 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 9758 46350
rect 9138 46226 9758 46294
rect 9138 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 9758 46226
rect 9138 46102 9758 46170
rect 9138 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 9758 46102
rect 9138 45978 9758 46046
rect 9138 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 9758 45978
rect 9138 28350 9758 45922
rect 9138 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 9758 28350
rect 9138 28226 9758 28294
rect 9138 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 9758 28226
rect 9138 28102 9758 28170
rect 9138 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 9758 28102
rect 9138 27978 9758 28046
rect 9138 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 9758 27978
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 10350 9758 27922
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 9138 -1120 9758 9922
rect 16716 4228 16772 238742
rect 16716 4162 16772 4172
rect 18396 4228 18452 238922
rect 18396 4162 18452 4172
rect 21756 234478 21812 234488
rect 21756 4228 21812 234422
rect 26012 93268 26068 290556
rect 27692 289156 27748 289166
rect 26012 93202 26068 93212
rect 26796 234298 26852 234308
rect 21756 4162 21812 4172
rect 26796 4228 26852 234242
rect 27692 135604 27748 289100
rect 27692 135538 27748 135548
rect 29372 65044 29428 377342
rect 31052 107380 31108 378782
rect 36138 364350 36758 381922
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 568350 40478 585922
rect 39858 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 40478 568350
rect 39858 568226 40478 568294
rect 39858 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 40478 568226
rect 39858 568102 40478 568170
rect 39858 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 40478 568102
rect 39858 567978 40478 568046
rect 39858 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 40478 567978
rect 39858 550350 40478 567922
rect 39858 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 40478 550350
rect 39858 550226 40478 550294
rect 39858 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 40478 550226
rect 39858 550102 40478 550170
rect 39858 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 40478 550102
rect 39858 549978 40478 550046
rect 39858 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 40478 549978
rect 39858 532350 40478 549922
rect 66858 597212 67478 598268
rect 66858 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 67478 597212
rect 66858 597088 67478 597156
rect 66858 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 67478 597088
rect 66858 596964 67478 597032
rect 66858 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 67478 596964
rect 66858 596840 67478 596908
rect 66858 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 67478 596840
rect 66858 580350 67478 596784
rect 66858 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 67478 580350
rect 66858 580226 67478 580294
rect 66858 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 67478 580226
rect 66858 580102 67478 580170
rect 66858 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 67478 580102
rect 66858 579978 67478 580046
rect 66858 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 67478 579978
rect 66858 562350 67478 579922
rect 66858 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 67478 562350
rect 66858 562226 67478 562294
rect 66858 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 67478 562226
rect 66858 562102 67478 562170
rect 66858 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 67478 562102
rect 66858 561978 67478 562046
rect 66858 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 67478 561978
rect 66858 544350 67478 561922
rect 66858 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 67478 544350
rect 66858 544226 67478 544294
rect 66858 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 67478 544226
rect 66858 544102 67478 544170
rect 66858 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 67478 544102
rect 66858 543978 67478 544046
rect 66858 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 67478 543978
rect 66858 535792 67478 543922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 568350 71198 585922
rect 70578 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 71198 568350
rect 70578 568226 71198 568294
rect 70578 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 71198 568226
rect 70578 568102 71198 568170
rect 70578 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 71198 568102
rect 70578 567978 71198 568046
rect 70578 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 71198 567978
rect 70578 550350 71198 567922
rect 70578 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 71198 550350
rect 70578 550226 71198 550294
rect 70578 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 71198 550226
rect 70578 550102 71198 550170
rect 70578 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 71198 550102
rect 70578 549978 71198 550046
rect 70578 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 71198 549978
rect 70578 539752 71198 549922
rect 97578 597212 98198 598268
rect 97578 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 98198 597212
rect 97578 597088 98198 597156
rect 97578 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 98198 597088
rect 97578 596964 98198 597032
rect 97578 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 98198 596964
rect 97578 596840 98198 596908
rect 97578 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 98198 596840
rect 97578 580350 98198 596784
rect 97578 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 98198 580350
rect 97578 580226 98198 580294
rect 97578 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 98198 580226
rect 97578 580102 98198 580170
rect 97578 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 98198 580102
rect 97578 579978 98198 580046
rect 97578 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 98198 579978
rect 97578 562350 98198 579922
rect 97578 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 98198 562350
rect 97578 562226 98198 562294
rect 97578 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 98198 562226
rect 97578 562102 98198 562170
rect 97578 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 98198 562102
rect 97578 561978 98198 562046
rect 97578 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 98198 561978
rect 97578 549832 98198 561922
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 101298 586350 101918 597744
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 101298 568350 101918 585922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 159018 597212 159638 598268
rect 159018 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 159638 597212
rect 159018 597088 159638 597156
rect 159018 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 159638 597088
rect 159018 596964 159638 597032
rect 159018 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 159638 596964
rect 159018 596840 159638 596908
rect 159018 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 159638 596840
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 130324 580063 130796 580120
rect 130324 580007 130346 580063
rect 130402 580007 130470 580063
rect 130526 580007 130594 580063
rect 130650 580007 130718 580063
rect 130774 580007 130796 580063
rect 130324 579939 130796 580007
rect 130324 579883 130346 579939
rect 130402 579883 130470 579939
rect 130526 579883 130594 579939
rect 130650 579883 130718 579939
rect 130774 579883 130796 579939
rect 130324 579826 130796 579883
rect 132018 578452 132638 585922
rect 157052 587188 157108 587198
rect 101298 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 101918 568350
rect 101298 568226 101918 568294
rect 101298 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 101918 568226
rect 101298 568102 101918 568170
rect 101298 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 101918 568102
rect 101298 567978 101918 568046
rect 101298 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 101918 567978
rect 101298 550350 101918 567922
rect 116160 562272 132720 562300
rect 116160 562216 116228 562272
rect 116284 562216 116352 562272
rect 116408 562216 116476 562272
rect 116532 562216 116600 562272
rect 116656 562216 116724 562272
rect 116780 562216 116848 562272
rect 116904 562216 116972 562272
rect 117028 562216 117096 562272
rect 117152 562216 117220 562272
rect 117276 562216 117344 562272
rect 117400 562216 117468 562272
rect 117524 562216 117592 562272
rect 117648 562216 117716 562272
rect 117772 562216 117840 562272
rect 117896 562216 117964 562272
rect 118020 562216 118088 562272
rect 118144 562216 118212 562272
rect 118268 562216 118336 562272
rect 118392 562216 118460 562272
rect 118516 562216 118584 562272
rect 118640 562216 118708 562272
rect 118764 562216 118832 562272
rect 118888 562216 118956 562272
rect 119012 562216 119080 562272
rect 119136 562216 119204 562272
rect 119260 562216 119328 562272
rect 119384 562216 119452 562272
rect 119508 562216 119576 562272
rect 119632 562216 119700 562272
rect 119756 562216 119824 562272
rect 119880 562216 119948 562272
rect 120004 562216 120072 562272
rect 120128 562216 120196 562272
rect 120252 562216 120320 562272
rect 120376 562216 120444 562272
rect 120500 562216 120568 562272
rect 120624 562216 120692 562272
rect 120748 562216 120816 562272
rect 120872 562216 120940 562272
rect 120996 562216 121064 562272
rect 121120 562216 121188 562272
rect 121244 562216 121312 562272
rect 121368 562216 121436 562272
rect 121492 562216 121560 562272
rect 121616 562216 121684 562272
rect 121740 562216 121808 562272
rect 121864 562216 121932 562272
rect 121988 562216 122056 562272
rect 122112 562216 122180 562272
rect 122236 562216 122304 562272
rect 122360 562216 122428 562272
rect 122484 562216 122552 562272
rect 122608 562216 122676 562272
rect 122732 562216 122800 562272
rect 122856 562216 122924 562272
rect 122980 562216 123048 562272
rect 123104 562216 123172 562272
rect 123228 562216 123296 562272
rect 123352 562216 123420 562272
rect 123476 562216 123544 562272
rect 123600 562216 123668 562272
rect 123724 562216 123792 562272
rect 123848 562216 123916 562272
rect 123972 562216 124040 562272
rect 124096 562216 124164 562272
rect 124220 562216 124288 562272
rect 124344 562216 124412 562272
rect 124468 562216 124536 562272
rect 124592 562216 124660 562272
rect 124716 562216 124784 562272
rect 124840 562216 124908 562272
rect 124964 562216 125032 562272
rect 125088 562216 125156 562272
rect 125212 562216 125280 562272
rect 125336 562216 125404 562272
rect 125460 562216 125528 562272
rect 125584 562216 125652 562272
rect 125708 562216 125776 562272
rect 125832 562216 125900 562272
rect 125956 562216 126024 562272
rect 126080 562216 126148 562272
rect 126204 562216 126272 562272
rect 126328 562216 126396 562272
rect 126452 562216 126520 562272
rect 126576 562216 126644 562272
rect 126700 562216 126768 562272
rect 126824 562216 126892 562272
rect 126948 562216 127016 562272
rect 127072 562216 127140 562272
rect 127196 562216 127264 562272
rect 127320 562216 127388 562272
rect 127444 562216 127512 562272
rect 127568 562216 127636 562272
rect 127692 562216 127760 562272
rect 127816 562216 127884 562272
rect 127940 562216 128008 562272
rect 128064 562216 128132 562272
rect 128188 562216 128256 562272
rect 128312 562216 128380 562272
rect 128436 562216 128504 562272
rect 128560 562216 128628 562272
rect 128684 562216 128752 562272
rect 128808 562216 128876 562272
rect 128932 562216 129000 562272
rect 129056 562216 129124 562272
rect 129180 562216 129248 562272
rect 129304 562216 129372 562272
rect 129428 562216 129496 562272
rect 129552 562216 129620 562272
rect 129676 562216 129744 562272
rect 129800 562216 129868 562272
rect 129924 562216 129992 562272
rect 130048 562216 130116 562272
rect 130172 562216 130240 562272
rect 130296 562216 130364 562272
rect 130420 562216 130488 562272
rect 130544 562216 130612 562272
rect 130668 562216 130736 562272
rect 130792 562216 130860 562272
rect 130916 562216 130984 562272
rect 131040 562216 131108 562272
rect 131164 562216 131232 562272
rect 131288 562216 131356 562272
rect 131412 562216 131480 562272
rect 131536 562216 131604 562272
rect 131660 562216 131728 562272
rect 131784 562216 131852 562272
rect 131908 562216 131976 562272
rect 132032 562216 132100 562272
rect 132156 562216 132224 562272
rect 132280 562216 132348 562272
rect 132404 562216 132472 562272
rect 132528 562216 132596 562272
rect 132652 562216 132720 562272
rect 116160 562148 132720 562216
rect 116160 562092 116228 562148
rect 116284 562092 116352 562148
rect 116408 562092 116476 562148
rect 116532 562092 116600 562148
rect 116656 562092 116724 562148
rect 116780 562092 116848 562148
rect 116904 562092 116972 562148
rect 117028 562092 117096 562148
rect 117152 562092 117220 562148
rect 117276 562092 117344 562148
rect 117400 562092 117468 562148
rect 117524 562092 117592 562148
rect 117648 562092 117716 562148
rect 117772 562092 117840 562148
rect 117896 562092 117964 562148
rect 118020 562092 118088 562148
rect 118144 562092 118212 562148
rect 118268 562092 118336 562148
rect 118392 562092 118460 562148
rect 118516 562092 118584 562148
rect 118640 562092 118708 562148
rect 118764 562092 118832 562148
rect 118888 562092 118956 562148
rect 119012 562092 119080 562148
rect 119136 562092 119204 562148
rect 119260 562092 119328 562148
rect 119384 562092 119452 562148
rect 119508 562092 119576 562148
rect 119632 562092 119700 562148
rect 119756 562092 119824 562148
rect 119880 562092 119948 562148
rect 120004 562092 120072 562148
rect 120128 562092 120196 562148
rect 120252 562092 120320 562148
rect 120376 562092 120444 562148
rect 120500 562092 120568 562148
rect 120624 562092 120692 562148
rect 120748 562092 120816 562148
rect 120872 562092 120940 562148
rect 120996 562092 121064 562148
rect 121120 562092 121188 562148
rect 121244 562092 121312 562148
rect 121368 562092 121436 562148
rect 121492 562092 121560 562148
rect 121616 562092 121684 562148
rect 121740 562092 121808 562148
rect 121864 562092 121932 562148
rect 121988 562092 122056 562148
rect 122112 562092 122180 562148
rect 122236 562092 122304 562148
rect 122360 562092 122428 562148
rect 122484 562092 122552 562148
rect 122608 562092 122676 562148
rect 122732 562092 122800 562148
rect 122856 562092 122924 562148
rect 122980 562092 123048 562148
rect 123104 562092 123172 562148
rect 123228 562092 123296 562148
rect 123352 562092 123420 562148
rect 123476 562092 123544 562148
rect 123600 562092 123668 562148
rect 123724 562092 123792 562148
rect 123848 562092 123916 562148
rect 123972 562092 124040 562148
rect 124096 562092 124164 562148
rect 124220 562092 124288 562148
rect 124344 562092 124412 562148
rect 124468 562092 124536 562148
rect 124592 562092 124660 562148
rect 124716 562092 124784 562148
rect 124840 562092 124908 562148
rect 124964 562092 125032 562148
rect 125088 562092 125156 562148
rect 125212 562092 125280 562148
rect 125336 562092 125404 562148
rect 125460 562092 125528 562148
rect 125584 562092 125652 562148
rect 125708 562092 125776 562148
rect 125832 562092 125900 562148
rect 125956 562092 126024 562148
rect 126080 562092 126148 562148
rect 126204 562092 126272 562148
rect 126328 562092 126396 562148
rect 126452 562092 126520 562148
rect 126576 562092 126644 562148
rect 126700 562092 126768 562148
rect 126824 562092 126892 562148
rect 126948 562092 127016 562148
rect 127072 562092 127140 562148
rect 127196 562092 127264 562148
rect 127320 562092 127388 562148
rect 127444 562092 127512 562148
rect 127568 562092 127636 562148
rect 127692 562092 127760 562148
rect 127816 562092 127884 562148
rect 127940 562092 128008 562148
rect 128064 562092 128132 562148
rect 128188 562092 128256 562148
rect 128312 562092 128380 562148
rect 128436 562092 128504 562148
rect 128560 562092 128628 562148
rect 128684 562092 128752 562148
rect 128808 562092 128876 562148
rect 128932 562092 129000 562148
rect 129056 562092 129124 562148
rect 129180 562092 129248 562148
rect 129304 562092 129372 562148
rect 129428 562092 129496 562148
rect 129552 562092 129620 562148
rect 129676 562092 129744 562148
rect 129800 562092 129868 562148
rect 129924 562092 129992 562148
rect 130048 562092 130116 562148
rect 130172 562092 130240 562148
rect 130296 562092 130364 562148
rect 130420 562092 130488 562148
rect 130544 562092 130612 562148
rect 130668 562092 130736 562148
rect 130792 562092 130860 562148
rect 130916 562092 130984 562148
rect 131040 562092 131108 562148
rect 131164 562092 131232 562148
rect 131288 562092 131356 562148
rect 131412 562092 131480 562148
rect 131536 562092 131604 562148
rect 131660 562092 131728 562148
rect 131784 562092 131852 562148
rect 131908 562092 131976 562148
rect 132032 562092 132100 562148
rect 132156 562092 132224 562148
rect 132280 562092 132348 562148
rect 132404 562092 132472 562148
rect 132528 562092 132596 562148
rect 132652 562092 132720 562148
rect 116160 562024 132720 562092
rect 116160 561968 116228 562024
rect 116284 561968 116352 562024
rect 116408 561968 116476 562024
rect 116532 561968 116600 562024
rect 116656 561968 116724 562024
rect 116780 561968 116848 562024
rect 116904 561968 116972 562024
rect 117028 561968 117096 562024
rect 117152 561968 117220 562024
rect 117276 561968 117344 562024
rect 117400 561968 117468 562024
rect 117524 561968 117592 562024
rect 117648 561968 117716 562024
rect 117772 561968 117840 562024
rect 117896 561968 117964 562024
rect 118020 561968 118088 562024
rect 118144 561968 118212 562024
rect 118268 561968 118336 562024
rect 118392 561968 118460 562024
rect 118516 561968 118584 562024
rect 118640 561968 118708 562024
rect 118764 561968 118832 562024
rect 118888 561968 118956 562024
rect 119012 561968 119080 562024
rect 119136 561968 119204 562024
rect 119260 561968 119328 562024
rect 119384 561968 119452 562024
rect 119508 561968 119576 562024
rect 119632 561968 119700 562024
rect 119756 561968 119824 562024
rect 119880 561968 119948 562024
rect 120004 561968 120072 562024
rect 120128 561968 120196 562024
rect 120252 561968 120320 562024
rect 120376 561968 120444 562024
rect 120500 561968 120568 562024
rect 120624 561968 120692 562024
rect 120748 561968 120816 562024
rect 120872 561968 120940 562024
rect 120996 561968 121064 562024
rect 121120 561968 121188 562024
rect 121244 561968 121312 562024
rect 121368 561968 121436 562024
rect 121492 561968 121560 562024
rect 121616 561968 121684 562024
rect 121740 561968 121808 562024
rect 121864 561968 121932 562024
rect 121988 561968 122056 562024
rect 122112 561968 122180 562024
rect 122236 561968 122304 562024
rect 122360 561968 122428 562024
rect 122484 561968 122552 562024
rect 122608 561968 122676 562024
rect 122732 561968 122800 562024
rect 122856 561968 122924 562024
rect 122980 561968 123048 562024
rect 123104 561968 123172 562024
rect 123228 561968 123296 562024
rect 123352 561968 123420 562024
rect 123476 561968 123544 562024
rect 123600 561968 123668 562024
rect 123724 561968 123792 562024
rect 123848 561968 123916 562024
rect 123972 561968 124040 562024
rect 124096 561968 124164 562024
rect 124220 561968 124288 562024
rect 124344 561968 124412 562024
rect 124468 561968 124536 562024
rect 124592 561968 124660 562024
rect 124716 561968 124784 562024
rect 124840 561968 124908 562024
rect 124964 561968 125032 562024
rect 125088 561968 125156 562024
rect 125212 561968 125280 562024
rect 125336 561968 125404 562024
rect 125460 561968 125528 562024
rect 125584 561968 125652 562024
rect 125708 561968 125776 562024
rect 125832 561968 125900 562024
rect 125956 561968 126024 562024
rect 126080 561968 126148 562024
rect 126204 561968 126272 562024
rect 126328 561968 126396 562024
rect 126452 561968 126520 562024
rect 126576 561968 126644 562024
rect 126700 561968 126768 562024
rect 126824 561968 126892 562024
rect 126948 561968 127016 562024
rect 127072 561968 127140 562024
rect 127196 561968 127264 562024
rect 127320 561968 127388 562024
rect 127444 561968 127512 562024
rect 127568 561968 127636 562024
rect 127692 561968 127760 562024
rect 127816 561968 127884 562024
rect 127940 561968 128008 562024
rect 128064 561968 128132 562024
rect 128188 561968 128256 562024
rect 128312 561968 128380 562024
rect 128436 561968 128504 562024
rect 128560 561968 128628 562024
rect 128684 561968 128752 562024
rect 128808 561968 128876 562024
rect 128932 561968 129000 562024
rect 129056 561968 129124 562024
rect 129180 561968 129248 562024
rect 129304 561968 129372 562024
rect 129428 561968 129496 562024
rect 129552 561968 129620 562024
rect 129676 561968 129744 562024
rect 129800 561968 129868 562024
rect 129924 561968 129992 562024
rect 130048 561968 130116 562024
rect 130172 561968 130240 562024
rect 130296 561968 130364 562024
rect 130420 561968 130488 562024
rect 130544 561968 130612 562024
rect 130668 561968 130736 562024
rect 130792 561968 130860 562024
rect 130916 561968 130984 562024
rect 131040 561968 131108 562024
rect 131164 561968 131232 562024
rect 131288 561968 131356 562024
rect 131412 561968 131480 562024
rect 131536 561968 131604 562024
rect 131660 561968 131728 562024
rect 131784 561968 131852 562024
rect 131908 561968 131976 562024
rect 132032 561968 132100 562024
rect 132156 561968 132224 562024
rect 132280 561968 132348 562024
rect 132404 561968 132472 562024
rect 132528 561968 132596 562024
rect 132652 561968 132720 562024
rect 116160 561940 132720 561968
rect 101298 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 101918 550350
rect 101298 550226 101918 550294
rect 101298 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 101918 550226
rect 101298 550102 101918 550170
rect 101298 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 101918 550102
rect 101298 549978 101918 550046
rect 101298 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 101918 549978
rect 101298 549472 101918 549922
rect 104280 544058 126420 544120
rect 104280 544002 104348 544058
rect 104404 544002 104472 544058
rect 104528 544002 104596 544058
rect 104652 544002 104720 544058
rect 104776 544002 104844 544058
rect 104900 544002 104968 544058
rect 105024 544002 105092 544058
rect 105148 544002 105216 544058
rect 105272 544002 105340 544058
rect 105396 544002 105464 544058
rect 105520 544002 105588 544058
rect 105644 544002 105712 544058
rect 105768 544002 105836 544058
rect 105892 544002 105960 544058
rect 106016 544002 106084 544058
rect 106140 544002 106208 544058
rect 106264 544002 106332 544058
rect 106388 544002 106456 544058
rect 106512 544002 106580 544058
rect 106636 544002 106704 544058
rect 106760 544002 106828 544058
rect 106884 544002 106952 544058
rect 107008 544002 107076 544058
rect 107132 544002 107200 544058
rect 107256 544002 107324 544058
rect 107380 544002 107448 544058
rect 107504 544002 107572 544058
rect 107628 544002 107696 544058
rect 107752 544002 107820 544058
rect 107876 544002 107944 544058
rect 108000 544002 108068 544058
rect 108124 544002 108192 544058
rect 108248 544002 108316 544058
rect 108372 544002 108440 544058
rect 108496 544002 108564 544058
rect 108620 544002 108688 544058
rect 108744 544002 108812 544058
rect 108868 544002 108936 544058
rect 108992 544002 109060 544058
rect 109116 544002 109184 544058
rect 109240 544002 109308 544058
rect 109364 544002 109432 544058
rect 109488 544002 109556 544058
rect 109612 544002 109680 544058
rect 109736 544002 109804 544058
rect 109860 544002 109928 544058
rect 109984 544002 110052 544058
rect 110108 544002 110176 544058
rect 110232 544002 110300 544058
rect 110356 544002 110424 544058
rect 110480 544002 110548 544058
rect 110604 544002 110672 544058
rect 110728 544002 110796 544058
rect 110852 544002 110920 544058
rect 110976 544002 111044 544058
rect 111100 544002 111168 544058
rect 111224 544002 111292 544058
rect 111348 544002 111416 544058
rect 111472 544002 111540 544058
rect 111596 544002 111664 544058
rect 111720 544002 111788 544058
rect 111844 544002 111912 544058
rect 111968 544002 112036 544058
rect 112092 544002 112160 544058
rect 112216 544002 112284 544058
rect 112340 544002 112408 544058
rect 112464 544002 112532 544058
rect 112588 544002 112656 544058
rect 112712 544002 112780 544058
rect 112836 544002 112904 544058
rect 112960 544002 113028 544058
rect 113084 544002 113152 544058
rect 113208 544002 113276 544058
rect 113332 544002 113400 544058
rect 113456 544002 113524 544058
rect 113580 544002 113648 544058
rect 113704 544002 113772 544058
rect 113828 544002 113896 544058
rect 113952 544002 114020 544058
rect 114076 544002 114144 544058
rect 114200 544002 114268 544058
rect 114324 544002 114392 544058
rect 114448 544002 114516 544058
rect 114572 544002 114640 544058
rect 114696 544002 114764 544058
rect 114820 544002 114888 544058
rect 114944 544002 115012 544058
rect 115068 544002 115136 544058
rect 115192 544002 115260 544058
rect 115316 544002 115384 544058
rect 115440 544002 115508 544058
rect 115564 544002 115632 544058
rect 115688 544002 115756 544058
rect 115812 544002 115880 544058
rect 115936 544002 116004 544058
rect 116060 544002 116128 544058
rect 116184 544002 116252 544058
rect 116308 544002 116376 544058
rect 116432 544002 116500 544058
rect 116556 544002 116624 544058
rect 116680 544002 116748 544058
rect 116804 544002 116872 544058
rect 116928 544002 116996 544058
rect 117052 544002 117120 544058
rect 117176 544002 117244 544058
rect 117300 544002 117368 544058
rect 117424 544002 117492 544058
rect 117548 544002 117616 544058
rect 117672 544002 117740 544058
rect 117796 544002 117864 544058
rect 117920 544002 117988 544058
rect 118044 544002 118112 544058
rect 118168 544002 118236 544058
rect 118292 544002 118360 544058
rect 118416 544002 118484 544058
rect 118540 544002 118608 544058
rect 118664 544002 118732 544058
rect 118788 544002 118856 544058
rect 118912 544002 118980 544058
rect 119036 544002 119104 544058
rect 119160 544002 119228 544058
rect 119284 544002 119352 544058
rect 119408 544002 119476 544058
rect 119532 544002 119600 544058
rect 119656 544002 119724 544058
rect 119780 544002 119848 544058
rect 119904 544002 119972 544058
rect 120028 544002 120096 544058
rect 120152 544002 120220 544058
rect 120276 544002 120344 544058
rect 120400 544002 120468 544058
rect 120524 544002 120592 544058
rect 120648 544002 120716 544058
rect 120772 544002 120840 544058
rect 120896 544002 120964 544058
rect 121020 544002 121088 544058
rect 121144 544002 121212 544058
rect 121268 544002 121336 544058
rect 121392 544002 121460 544058
rect 121516 544002 121584 544058
rect 121640 544002 121708 544058
rect 121764 544002 121832 544058
rect 121888 544002 121956 544058
rect 122012 544002 122080 544058
rect 122136 544002 122204 544058
rect 122260 544002 122328 544058
rect 122384 544002 122452 544058
rect 122508 544002 122576 544058
rect 122632 544002 122700 544058
rect 122756 544002 122824 544058
rect 122880 544002 122948 544058
rect 123004 544002 123072 544058
rect 123128 544002 123196 544058
rect 123252 544002 123320 544058
rect 123376 544002 123444 544058
rect 123500 544002 123568 544058
rect 123624 544002 123692 544058
rect 123748 544002 123816 544058
rect 123872 544002 123940 544058
rect 123996 544002 124064 544058
rect 124120 544002 124188 544058
rect 124244 544002 124312 544058
rect 124368 544002 124436 544058
rect 124492 544002 124560 544058
rect 124616 544002 124684 544058
rect 124740 544002 124808 544058
rect 124864 544002 124932 544058
rect 124988 544002 125056 544058
rect 125112 544002 125180 544058
rect 125236 544002 125304 544058
rect 125360 544002 125428 544058
rect 125484 544002 125552 544058
rect 125608 544002 125676 544058
rect 125732 544002 125800 544058
rect 125856 544002 125924 544058
rect 125980 544002 126048 544058
rect 126104 544002 126172 544058
rect 126228 544002 126296 544058
rect 126352 544002 126420 544058
rect 104280 543940 126420 544002
rect 39858 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532294 40478 532350
rect 39858 532226 40478 532294
rect 66660 532358 74760 532420
rect 66660 532302 66714 532358
rect 66770 532302 66838 532358
rect 66894 532302 66962 532358
rect 67018 532302 67086 532358
rect 67142 532302 67210 532358
rect 67266 532302 67334 532358
rect 67390 532302 67458 532358
rect 67514 532302 67582 532358
rect 67638 532302 67706 532358
rect 67762 532302 67830 532358
rect 67886 532302 67954 532358
rect 68010 532302 68078 532358
rect 68134 532302 68202 532358
rect 68258 532302 68326 532358
rect 68382 532302 68450 532358
rect 68506 532302 68574 532358
rect 68630 532302 68698 532358
rect 68754 532302 68822 532358
rect 68878 532302 68946 532358
rect 69002 532302 69070 532358
rect 69126 532302 69194 532358
rect 69250 532302 69318 532358
rect 69374 532302 69442 532358
rect 69498 532302 69566 532358
rect 69622 532302 69690 532358
rect 69746 532302 69814 532358
rect 69870 532302 69938 532358
rect 69994 532302 70062 532358
rect 70118 532302 70186 532358
rect 70242 532302 70310 532358
rect 70366 532302 70434 532358
rect 70490 532302 70558 532358
rect 70614 532302 70682 532358
rect 70738 532302 70806 532358
rect 70862 532302 70930 532358
rect 70986 532302 71054 532358
rect 71110 532302 71178 532358
rect 71234 532302 71302 532358
rect 71358 532302 71426 532358
rect 71482 532302 71550 532358
rect 71606 532302 71674 532358
rect 71730 532302 71798 532358
rect 71854 532302 71922 532358
rect 71978 532302 72046 532358
rect 72102 532302 72170 532358
rect 72226 532302 72294 532358
rect 72350 532302 72418 532358
rect 72474 532302 72542 532358
rect 72598 532302 72666 532358
rect 72722 532302 72790 532358
rect 72846 532302 72914 532358
rect 72970 532302 73038 532358
rect 73094 532302 73162 532358
rect 73218 532302 73286 532358
rect 73342 532302 73410 532358
rect 73466 532302 73534 532358
rect 73590 532302 73658 532358
rect 73714 532302 73782 532358
rect 73838 532302 73906 532358
rect 73962 532302 74030 532358
rect 74086 532302 74154 532358
rect 74210 532302 74278 532358
rect 74334 532302 74402 532358
rect 74458 532302 74526 532358
rect 74582 532302 74650 532358
rect 74706 532302 74760 532358
rect 66660 532240 74760 532302
rect 39858 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 40478 532226
rect 39858 532102 40478 532170
rect 39858 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 40478 532102
rect 39858 531978 40478 532046
rect 39858 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 40478 531978
rect 39858 514350 40478 531922
rect 66480 531998 66960 532060
rect 66480 531942 66506 531998
rect 66562 531942 66630 531998
rect 66686 531942 66754 531998
rect 66810 531942 66878 531998
rect 66934 531942 66960 531998
rect 66480 531880 66960 531942
rect 66976 531998 67456 532060
rect 66976 531942 67002 531998
rect 67058 531942 67126 531998
rect 67182 531942 67250 531998
rect 67306 531942 67374 531998
rect 67430 531942 67456 531998
rect 66976 531880 67456 531942
rect 67472 531998 67952 532060
rect 67472 531942 67498 531998
rect 67554 531942 67622 531998
rect 67678 531942 67746 531998
rect 67802 531942 67870 531998
rect 67926 531942 67952 531998
rect 67472 531880 67952 531942
rect 67968 531998 68448 532060
rect 67968 531942 67994 531998
rect 68050 531942 68118 531998
rect 68174 531942 68242 531998
rect 68298 531942 68366 531998
rect 68422 531942 68448 531998
rect 67968 531880 68448 531942
rect 68464 531998 68944 532060
rect 68464 531942 68490 531998
rect 68546 531942 68614 531998
rect 68670 531942 68738 531998
rect 68794 531942 68862 531998
rect 68918 531942 68944 531998
rect 68464 531880 68944 531942
rect 68960 531998 69440 532060
rect 68960 531942 68986 531998
rect 69042 531942 69110 531998
rect 69166 531942 69234 531998
rect 69290 531942 69358 531998
rect 69414 531942 69440 531998
rect 68960 531880 69440 531942
rect 69456 531998 69936 532060
rect 69456 531942 69482 531998
rect 69538 531942 69606 531998
rect 69662 531942 69730 531998
rect 69786 531942 69854 531998
rect 69910 531942 69936 531998
rect 69456 531880 69936 531942
rect 69952 531998 70432 532060
rect 69952 531942 69978 531998
rect 70034 531942 70102 531998
rect 70158 531942 70226 531998
rect 70282 531942 70350 531998
rect 70406 531942 70432 531998
rect 69952 531880 70432 531942
rect 70448 531998 70928 532060
rect 70448 531942 70474 531998
rect 70530 531942 70598 531998
rect 70654 531942 70722 531998
rect 70778 531942 70846 531998
rect 70902 531942 70928 531998
rect 70448 531880 70928 531942
rect 70944 531998 71424 532060
rect 70944 531942 70970 531998
rect 71026 531942 71094 531998
rect 71150 531942 71218 531998
rect 71274 531942 71342 531998
rect 71398 531942 71424 531998
rect 70944 531880 71424 531942
rect 71440 531998 71920 532060
rect 71440 531942 71466 531998
rect 71522 531942 71590 531998
rect 71646 531942 71714 531998
rect 71770 531942 71838 531998
rect 71894 531942 71920 531998
rect 71440 531880 71920 531942
rect 71936 531998 72416 532060
rect 71936 531942 71962 531998
rect 72018 531942 72086 531998
rect 72142 531942 72210 531998
rect 72266 531942 72334 531998
rect 72390 531942 72416 531998
rect 71936 531880 72416 531942
rect 72432 531998 72912 532060
rect 72432 531942 72458 531998
rect 72514 531942 72582 531998
rect 72638 531942 72706 531998
rect 72762 531942 72830 531998
rect 72886 531942 72912 531998
rect 72432 531880 72912 531942
rect 72928 531998 73408 532060
rect 72928 531942 72954 531998
rect 73010 531942 73078 531998
rect 73134 531942 73202 531998
rect 73258 531942 73326 531998
rect 73382 531942 73408 531998
rect 72928 531880 73408 531942
rect 73424 531998 73904 532060
rect 73424 531942 73450 531998
rect 73506 531942 73574 531998
rect 73630 531942 73698 531998
rect 73754 531942 73822 531998
rect 73878 531942 73904 531998
rect 73424 531880 73904 531942
rect 73920 531998 74400 532060
rect 73920 531942 73946 531998
rect 74002 531942 74070 531998
rect 74126 531942 74194 531998
rect 74250 531942 74318 531998
rect 74374 531942 74400 531998
rect 73920 531880 74400 531942
rect 96000 526238 96232 526300
rect 96000 526182 96026 526238
rect 96082 526182 96150 526238
rect 96206 526182 96232 526238
rect 96000 526120 96232 526182
rect 96248 526238 96728 526300
rect 96248 526182 96274 526238
rect 96330 526182 96398 526238
rect 96454 526182 96522 526238
rect 96578 526182 96646 526238
rect 96702 526182 96728 526238
rect 96248 526120 96728 526182
rect 96744 526238 97224 526300
rect 96744 526182 96770 526238
rect 96826 526182 96894 526238
rect 96950 526182 97018 526238
rect 97074 526182 97142 526238
rect 97198 526182 97224 526238
rect 96744 526120 97224 526182
rect 97240 526238 97720 526300
rect 97240 526182 97266 526238
rect 97322 526182 97390 526238
rect 97446 526182 97514 526238
rect 97570 526182 97638 526238
rect 97694 526182 97720 526238
rect 97240 526120 97720 526182
rect 97736 526238 98216 526300
rect 97736 526182 97762 526238
rect 97818 526182 97886 526238
rect 97942 526182 98010 526238
rect 98066 526182 98134 526238
rect 98190 526182 98216 526238
rect 97736 526120 98216 526182
rect 98232 526238 98712 526300
rect 98232 526182 98258 526238
rect 98314 526182 98382 526238
rect 98438 526182 98506 526238
rect 98562 526182 98630 526238
rect 98686 526182 98712 526238
rect 98232 526120 98712 526182
rect 98728 526238 99208 526300
rect 98728 526182 98754 526238
rect 98810 526182 98878 526238
rect 98934 526182 99002 526238
rect 99058 526182 99126 526238
rect 99182 526182 99208 526238
rect 98728 526120 99208 526182
rect 99224 526238 99704 526300
rect 99224 526182 99250 526238
rect 99306 526182 99374 526238
rect 99430 526182 99498 526238
rect 99554 526182 99622 526238
rect 99678 526182 99704 526238
rect 99224 526120 99704 526182
rect 99720 526238 100200 526300
rect 99720 526182 99746 526238
rect 99802 526182 99870 526238
rect 99926 526182 99994 526238
rect 100050 526182 100118 526238
rect 100174 526182 100200 526238
rect 99720 526120 100200 526182
rect 100216 526238 100696 526300
rect 100216 526182 100242 526238
rect 100298 526182 100366 526238
rect 100422 526182 100490 526238
rect 100546 526182 100614 526238
rect 100670 526182 100696 526238
rect 100216 526120 100696 526182
rect 100712 526238 101192 526300
rect 100712 526182 100738 526238
rect 100794 526182 100862 526238
rect 100918 526182 100986 526238
rect 101042 526182 101110 526238
rect 101166 526182 101192 526238
rect 100712 526120 101192 526182
rect 101208 526238 101688 526300
rect 101208 526182 101234 526238
rect 101290 526182 101358 526238
rect 101414 526182 101482 526238
rect 101538 526182 101606 526238
rect 101662 526182 101688 526238
rect 101208 526120 101688 526182
rect 101704 526238 102184 526300
rect 101704 526182 101730 526238
rect 101786 526182 101854 526238
rect 101910 526182 101978 526238
rect 102034 526182 102102 526238
rect 102158 526182 102184 526238
rect 101704 526120 102184 526182
rect 102200 526238 102680 526300
rect 102200 526182 102226 526238
rect 102282 526182 102350 526238
rect 102406 526182 102474 526238
rect 102530 526182 102598 526238
rect 102654 526182 102680 526238
rect 102200 526120 102680 526182
rect 102696 526238 103176 526300
rect 102696 526182 102722 526238
rect 102778 526182 102846 526238
rect 102902 526182 102970 526238
rect 103026 526182 103094 526238
rect 103150 526182 103176 526238
rect 102696 526120 103176 526182
rect 103192 526238 103672 526300
rect 103192 526182 103218 526238
rect 103274 526182 103342 526238
rect 103398 526182 103466 526238
rect 103522 526182 103590 526238
rect 103646 526182 103672 526238
rect 103192 526120 103672 526182
rect 103688 526238 104168 526300
rect 103688 526182 103714 526238
rect 103770 526182 103838 526238
rect 103894 526182 103962 526238
rect 104018 526182 104086 526238
rect 104142 526182 104168 526238
rect 103688 526120 104168 526182
rect 104184 526238 104664 526300
rect 104184 526182 104210 526238
rect 104266 526182 104334 526238
rect 104390 526182 104458 526238
rect 104514 526182 104582 526238
rect 104638 526182 104664 526238
rect 104184 526120 104664 526182
rect 104680 526238 105160 526300
rect 104680 526182 104706 526238
rect 104762 526182 104830 526238
rect 104886 526182 104954 526238
rect 105010 526182 105078 526238
rect 105134 526182 105160 526238
rect 104680 526120 105160 526182
rect 105176 526238 105656 526300
rect 105176 526182 105202 526238
rect 105258 526182 105326 526238
rect 105382 526182 105450 526238
rect 105506 526182 105574 526238
rect 105630 526182 105656 526238
rect 105176 526120 105656 526182
rect 105672 526238 106152 526300
rect 105672 526182 105698 526238
rect 105754 526182 105822 526238
rect 105878 526182 105946 526238
rect 106002 526182 106070 526238
rect 106126 526182 106152 526238
rect 105672 526120 106152 526182
rect 106168 526238 106648 526300
rect 106168 526182 106194 526238
rect 106250 526182 106318 526238
rect 106374 526182 106442 526238
rect 106498 526182 106566 526238
rect 106622 526182 106648 526238
rect 106168 526120 106648 526182
rect 106664 526238 107144 526300
rect 106664 526182 106690 526238
rect 106746 526182 106814 526238
rect 106870 526182 106938 526238
rect 106994 526182 107062 526238
rect 107118 526182 107144 526238
rect 106664 526120 107144 526182
rect 107160 526238 107640 526300
rect 107160 526182 107186 526238
rect 107242 526182 107310 526238
rect 107366 526182 107434 526238
rect 107490 526182 107558 526238
rect 107614 526182 107640 526238
rect 107160 526120 107640 526182
rect 107656 526238 108136 526300
rect 107656 526182 107682 526238
rect 107738 526182 107806 526238
rect 107862 526182 107930 526238
rect 107986 526182 108054 526238
rect 108110 526182 108136 526238
rect 107656 526120 108136 526182
rect 108152 526238 108632 526300
rect 108152 526182 108178 526238
rect 108234 526182 108302 526238
rect 108358 526182 108426 526238
rect 108482 526182 108550 526238
rect 108606 526182 108632 526238
rect 108152 526120 108632 526182
rect 108648 526238 109128 526300
rect 108648 526182 108674 526238
rect 108730 526182 108798 526238
rect 108854 526182 108922 526238
rect 108978 526182 109046 526238
rect 109102 526182 109128 526238
rect 108648 526120 109128 526182
rect 109144 526238 109624 526300
rect 109144 526182 109170 526238
rect 109226 526182 109294 526238
rect 109350 526182 109418 526238
rect 109474 526182 109542 526238
rect 109598 526182 109624 526238
rect 109144 526120 109624 526182
rect 109640 526238 110120 526300
rect 109640 526182 109666 526238
rect 109722 526182 109790 526238
rect 109846 526182 109914 526238
rect 109970 526182 110038 526238
rect 110094 526182 110120 526238
rect 109640 526120 110120 526182
rect 110136 526238 110616 526300
rect 110136 526182 110162 526238
rect 110218 526182 110286 526238
rect 110342 526182 110410 526238
rect 110466 526182 110534 526238
rect 110590 526182 110616 526238
rect 110136 526120 110616 526182
rect 110632 526238 111112 526300
rect 110632 526182 110658 526238
rect 110714 526182 110782 526238
rect 110838 526182 110906 526238
rect 110962 526182 111030 526238
rect 111086 526182 111112 526238
rect 110632 526120 111112 526182
rect 111128 526238 111608 526300
rect 111128 526182 111154 526238
rect 111210 526182 111278 526238
rect 111334 526182 111402 526238
rect 111458 526182 111526 526238
rect 111582 526182 111608 526238
rect 111128 526120 111608 526182
rect 111624 526238 112104 526300
rect 111624 526182 111650 526238
rect 111706 526182 111774 526238
rect 111830 526182 111898 526238
rect 111954 526182 112022 526238
rect 112078 526182 112104 526238
rect 111624 526120 112104 526182
rect 112120 526238 112600 526300
rect 112120 526182 112146 526238
rect 112202 526182 112270 526238
rect 112326 526182 112394 526238
rect 112450 526182 112518 526238
rect 112574 526182 112600 526238
rect 112120 526120 112600 526182
rect 112616 526238 113096 526300
rect 112616 526182 112642 526238
rect 112698 526182 112766 526238
rect 112822 526182 112890 526238
rect 112946 526182 113014 526238
rect 113070 526182 113096 526238
rect 112616 526120 113096 526182
rect 113112 526238 113592 526300
rect 113112 526182 113138 526238
rect 113194 526182 113262 526238
rect 113318 526182 113386 526238
rect 113442 526182 113510 526238
rect 113566 526182 113592 526238
rect 113112 526120 113592 526182
rect 113608 526238 114088 526300
rect 113608 526182 113634 526238
rect 113690 526182 113758 526238
rect 113814 526182 113882 526238
rect 113938 526182 114006 526238
rect 114062 526182 114088 526238
rect 113608 526120 114088 526182
rect 114104 526238 114584 526300
rect 114104 526182 114130 526238
rect 114186 526182 114254 526238
rect 114310 526182 114378 526238
rect 114434 526182 114502 526238
rect 114558 526182 114584 526238
rect 114104 526120 114584 526182
rect 114600 526238 115080 526300
rect 114600 526182 114626 526238
rect 114682 526182 114750 526238
rect 114806 526182 114874 526238
rect 114930 526182 114998 526238
rect 115054 526182 115080 526238
rect 114600 526120 115080 526182
rect 95820 525911 114720 525940
rect 95820 525855 95880 525911
rect 95936 525855 96004 525911
rect 96060 525855 96128 525911
rect 96184 525855 96252 525911
rect 96308 525855 96376 525911
rect 96432 525855 96500 525911
rect 96556 525855 96624 525911
rect 96680 525855 96748 525911
rect 96804 525855 96872 525911
rect 96928 525855 96996 525911
rect 97052 525855 97120 525911
rect 97176 525855 97244 525911
rect 97300 525855 97368 525911
rect 97424 525855 97492 525911
rect 97548 525855 97616 525911
rect 97672 525855 97740 525911
rect 97796 525855 97864 525911
rect 97920 525855 97988 525911
rect 98044 525855 98112 525911
rect 98168 525855 98236 525911
rect 98292 525855 98360 525911
rect 98416 525855 98484 525911
rect 98540 525855 98608 525911
rect 98664 525855 98732 525911
rect 98788 525855 98856 525911
rect 98912 525855 98980 525911
rect 99036 525855 99104 525911
rect 99160 525855 99228 525911
rect 99284 525855 99352 525911
rect 99408 525855 99476 525911
rect 99532 525855 99600 525911
rect 99656 525855 99724 525911
rect 99780 525855 99848 525911
rect 99904 525855 99972 525911
rect 100028 525855 100096 525911
rect 100152 525855 100220 525911
rect 100276 525855 100344 525911
rect 100400 525855 100468 525911
rect 100524 525855 100592 525911
rect 100648 525855 100716 525911
rect 100772 525855 100840 525911
rect 100896 525855 100964 525911
rect 101020 525855 101088 525911
rect 101144 525855 101212 525911
rect 101268 525855 101336 525911
rect 101392 525855 101460 525911
rect 101516 525855 101584 525911
rect 101640 525855 101708 525911
rect 101764 525855 101832 525911
rect 101888 525855 101956 525911
rect 102012 525855 102080 525911
rect 102136 525855 102204 525911
rect 102260 525855 102328 525911
rect 102384 525855 102452 525911
rect 102508 525855 102576 525911
rect 102632 525855 102700 525911
rect 102756 525855 102824 525911
rect 102880 525855 102948 525911
rect 103004 525855 103072 525911
rect 103128 525855 103196 525911
rect 103252 525855 103320 525911
rect 103376 525855 103444 525911
rect 103500 525855 103568 525911
rect 103624 525855 103692 525911
rect 103748 525855 103816 525911
rect 103872 525855 103940 525911
rect 103996 525855 104064 525911
rect 104120 525855 104188 525911
rect 104244 525855 104312 525911
rect 104368 525855 104436 525911
rect 104492 525855 104560 525911
rect 104616 525855 104684 525911
rect 104740 525855 104808 525911
rect 104864 525855 104932 525911
rect 104988 525855 105056 525911
rect 105112 525855 105180 525911
rect 105236 525855 105304 525911
rect 105360 525855 105428 525911
rect 105484 525855 105552 525911
rect 105608 525855 105676 525911
rect 105732 525855 105800 525911
rect 105856 525855 105924 525911
rect 105980 525855 106048 525911
rect 106104 525855 106172 525911
rect 106228 525855 106296 525911
rect 106352 525855 106420 525911
rect 106476 525855 106544 525911
rect 106600 525855 106668 525911
rect 106724 525855 106792 525911
rect 106848 525855 106916 525911
rect 106972 525855 107040 525911
rect 107096 525855 107164 525911
rect 107220 525855 107288 525911
rect 107344 525855 107412 525911
rect 107468 525855 107536 525911
rect 107592 525855 107660 525911
rect 107716 525855 107784 525911
rect 107840 525855 107908 525911
rect 107964 525855 108032 525911
rect 108088 525855 108156 525911
rect 108212 525855 108280 525911
rect 108336 525855 108404 525911
rect 108460 525855 108528 525911
rect 108584 525855 108652 525911
rect 108708 525855 108776 525911
rect 108832 525855 108900 525911
rect 108956 525855 109024 525911
rect 109080 525855 109148 525911
rect 109204 525855 109272 525911
rect 109328 525855 109396 525911
rect 109452 525855 109520 525911
rect 109576 525855 109644 525911
rect 109700 525855 109768 525911
rect 109824 525855 109892 525911
rect 109948 525855 110016 525911
rect 110072 525855 110140 525911
rect 110196 525855 110264 525911
rect 110320 525855 110388 525911
rect 110444 525855 110512 525911
rect 110568 525855 110636 525911
rect 110692 525855 110760 525911
rect 110816 525855 110884 525911
rect 110940 525855 111008 525911
rect 111064 525855 111132 525911
rect 111188 525855 111256 525911
rect 111312 525855 111380 525911
rect 111436 525855 111504 525911
rect 111560 525855 111628 525911
rect 111684 525855 111752 525911
rect 111808 525855 111876 525911
rect 111932 525855 112000 525911
rect 112056 525855 112124 525911
rect 112180 525855 112248 525911
rect 112304 525855 112372 525911
rect 112428 525855 112496 525911
rect 112552 525855 112620 525911
rect 112676 525855 112744 525911
rect 112800 525855 112868 525911
rect 112924 525855 112992 525911
rect 113048 525855 113116 525911
rect 113172 525855 113240 525911
rect 113296 525855 113364 525911
rect 113420 525855 113488 525911
rect 113544 525855 113612 525911
rect 113668 525855 113736 525911
rect 113792 525855 113860 525911
rect 113916 525855 113984 525911
rect 114040 525855 114108 525911
rect 114164 525855 114232 525911
rect 114288 525855 114356 525911
rect 114412 525855 114480 525911
rect 114536 525855 114604 525911
rect 114660 525855 114720 525911
rect 95820 525826 114720 525855
rect 39858 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 40478 514350
rect 39858 514226 40478 514294
rect 39858 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 40478 514226
rect 39858 514102 40478 514170
rect 39858 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 40478 514102
rect 39858 513978 40478 514046
rect 39858 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 40478 513978
rect 39858 496350 40478 513922
rect 60180 514412 60528 514446
rect 60180 514356 60202 514412
rect 60258 514356 60326 514412
rect 60382 514356 60450 514412
rect 60506 514356 60528 514412
rect 60180 514288 60528 514356
rect 60180 514232 60202 514288
rect 60258 514232 60326 514288
rect 60382 514232 60450 514288
rect 60506 514232 60528 514288
rect 60180 514164 60528 514232
rect 60180 514108 60202 514164
rect 60258 514108 60326 514164
rect 60382 514108 60450 514164
rect 60506 514108 60528 514164
rect 60180 514040 60528 514108
rect 60180 513984 60202 514040
rect 60258 513984 60326 514040
rect 60382 513984 60450 514040
rect 60506 513984 60528 514040
rect 60180 513916 60528 513984
rect 60180 513860 60202 513916
rect 60258 513860 60326 513916
rect 60382 513860 60450 513916
rect 60506 513860 60528 513916
rect 60180 513826 60528 513860
rect 60552 514412 61024 514446
rect 60552 514356 60574 514412
rect 60630 514356 60698 514412
rect 60754 514356 60822 514412
rect 60878 514356 60946 514412
rect 61002 514356 61024 514412
rect 60552 514288 61024 514356
rect 60552 514232 60574 514288
rect 60630 514232 60698 514288
rect 60754 514232 60822 514288
rect 60878 514232 60946 514288
rect 61002 514232 61024 514288
rect 60552 514164 61024 514232
rect 60552 514108 60574 514164
rect 60630 514108 60698 514164
rect 60754 514108 60822 514164
rect 60878 514108 60946 514164
rect 61002 514108 61024 514164
rect 60552 514040 61024 514108
rect 60552 513984 60574 514040
rect 60630 513984 60698 514040
rect 60754 513984 60822 514040
rect 60878 513984 60946 514040
rect 61002 513984 61024 514040
rect 60552 513916 61024 513984
rect 60552 513860 60574 513916
rect 60630 513860 60698 513916
rect 60754 513860 60822 513916
rect 60878 513860 60946 513916
rect 61002 513860 61024 513916
rect 60552 513826 61024 513860
rect 61048 514412 61520 514446
rect 61048 514356 61070 514412
rect 61126 514356 61194 514412
rect 61250 514356 61318 514412
rect 61374 514356 61442 514412
rect 61498 514356 61520 514412
rect 61048 514288 61520 514356
rect 61048 514232 61070 514288
rect 61126 514232 61194 514288
rect 61250 514232 61318 514288
rect 61374 514232 61442 514288
rect 61498 514232 61520 514288
rect 61048 514164 61520 514232
rect 61048 514108 61070 514164
rect 61126 514108 61194 514164
rect 61250 514108 61318 514164
rect 61374 514108 61442 514164
rect 61498 514108 61520 514164
rect 61048 514040 61520 514108
rect 61048 513984 61070 514040
rect 61126 513984 61194 514040
rect 61250 513984 61318 514040
rect 61374 513984 61442 514040
rect 61498 513984 61520 514040
rect 61048 513916 61520 513984
rect 61048 513860 61070 513916
rect 61126 513860 61194 513916
rect 61250 513860 61318 513916
rect 61374 513860 61442 513916
rect 61498 513860 61520 513916
rect 61048 513826 61520 513860
rect 61544 514412 62016 514446
rect 61544 514356 61566 514412
rect 61622 514356 61690 514412
rect 61746 514356 61814 514412
rect 61870 514356 61938 514412
rect 61994 514356 62016 514412
rect 61544 514288 62016 514356
rect 61544 514232 61566 514288
rect 61622 514232 61690 514288
rect 61746 514232 61814 514288
rect 61870 514232 61938 514288
rect 61994 514232 62016 514288
rect 61544 514164 62016 514232
rect 61544 514108 61566 514164
rect 61622 514108 61690 514164
rect 61746 514108 61814 514164
rect 61870 514108 61938 514164
rect 61994 514108 62016 514164
rect 61544 514040 62016 514108
rect 61544 513984 61566 514040
rect 61622 513984 61690 514040
rect 61746 513984 61814 514040
rect 61870 513984 61938 514040
rect 61994 513984 62016 514040
rect 61544 513916 62016 513984
rect 61544 513860 61566 513916
rect 61622 513860 61690 513916
rect 61746 513860 61814 513916
rect 61870 513860 61938 513916
rect 61994 513860 62016 513916
rect 61544 513826 62016 513860
rect 62040 514412 62512 514446
rect 62040 514356 62062 514412
rect 62118 514356 62186 514412
rect 62242 514356 62310 514412
rect 62366 514356 62434 514412
rect 62490 514356 62512 514412
rect 62040 514288 62512 514356
rect 62040 514232 62062 514288
rect 62118 514232 62186 514288
rect 62242 514232 62310 514288
rect 62366 514232 62434 514288
rect 62490 514232 62512 514288
rect 62040 514164 62512 514232
rect 62040 514108 62062 514164
rect 62118 514108 62186 514164
rect 62242 514108 62310 514164
rect 62366 514108 62434 514164
rect 62490 514108 62512 514164
rect 62040 514040 62512 514108
rect 62040 513984 62062 514040
rect 62118 513984 62186 514040
rect 62242 513984 62310 514040
rect 62366 513984 62434 514040
rect 62490 513984 62512 514040
rect 62040 513916 62512 513984
rect 62040 513860 62062 513916
rect 62118 513860 62186 513916
rect 62242 513860 62310 513916
rect 62366 513860 62434 513916
rect 62490 513860 62512 513916
rect 62040 513826 62512 513860
rect 62536 514412 63008 514446
rect 62536 514356 62558 514412
rect 62614 514356 62682 514412
rect 62738 514356 62806 514412
rect 62862 514356 62930 514412
rect 62986 514356 63008 514412
rect 62536 514288 63008 514356
rect 62536 514232 62558 514288
rect 62614 514232 62682 514288
rect 62738 514232 62806 514288
rect 62862 514232 62930 514288
rect 62986 514232 63008 514288
rect 62536 514164 63008 514232
rect 62536 514108 62558 514164
rect 62614 514108 62682 514164
rect 62738 514108 62806 514164
rect 62862 514108 62930 514164
rect 62986 514108 63008 514164
rect 62536 514040 63008 514108
rect 62536 513984 62558 514040
rect 62614 513984 62682 514040
rect 62738 513984 62806 514040
rect 62862 513984 62930 514040
rect 62986 513984 63008 514040
rect 62536 513916 63008 513984
rect 62536 513860 62558 513916
rect 62614 513860 62682 513916
rect 62738 513860 62806 513916
rect 62862 513860 62930 513916
rect 62986 513860 63008 513916
rect 62536 513826 63008 513860
rect 63032 514412 63504 514446
rect 63032 514356 63054 514412
rect 63110 514356 63178 514412
rect 63234 514356 63302 514412
rect 63358 514356 63426 514412
rect 63482 514356 63504 514412
rect 63032 514288 63504 514356
rect 63032 514232 63054 514288
rect 63110 514232 63178 514288
rect 63234 514232 63302 514288
rect 63358 514232 63426 514288
rect 63482 514232 63504 514288
rect 63032 514164 63504 514232
rect 63032 514108 63054 514164
rect 63110 514108 63178 514164
rect 63234 514108 63302 514164
rect 63358 514108 63426 514164
rect 63482 514108 63504 514164
rect 63032 514040 63504 514108
rect 63032 513984 63054 514040
rect 63110 513984 63178 514040
rect 63234 513984 63302 514040
rect 63358 513984 63426 514040
rect 63482 513984 63504 514040
rect 63032 513916 63504 513984
rect 63032 513860 63054 513916
rect 63110 513860 63178 513916
rect 63234 513860 63302 513916
rect 63358 513860 63426 513916
rect 63482 513860 63504 513916
rect 63032 513826 63504 513860
rect 63528 514412 64000 514446
rect 63528 514356 63550 514412
rect 63606 514356 63674 514412
rect 63730 514356 63798 514412
rect 63854 514356 63922 514412
rect 63978 514356 64000 514412
rect 63528 514288 64000 514356
rect 63528 514232 63550 514288
rect 63606 514232 63674 514288
rect 63730 514232 63798 514288
rect 63854 514232 63922 514288
rect 63978 514232 64000 514288
rect 63528 514164 64000 514232
rect 63528 514108 63550 514164
rect 63606 514108 63674 514164
rect 63730 514108 63798 514164
rect 63854 514108 63922 514164
rect 63978 514108 64000 514164
rect 63528 514040 64000 514108
rect 63528 513984 63550 514040
rect 63606 513984 63674 514040
rect 63730 513984 63798 514040
rect 63854 513984 63922 514040
rect 63978 513984 64000 514040
rect 63528 513916 64000 513984
rect 63528 513860 63550 513916
rect 63606 513860 63674 513916
rect 63730 513860 63798 513916
rect 63854 513860 63922 513916
rect 63978 513860 64000 513916
rect 63528 513826 64000 513860
rect 64024 514412 64496 514446
rect 64024 514356 64046 514412
rect 64102 514356 64170 514412
rect 64226 514356 64294 514412
rect 64350 514356 64418 514412
rect 64474 514356 64496 514412
rect 64024 514288 64496 514356
rect 64024 514232 64046 514288
rect 64102 514232 64170 514288
rect 64226 514232 64294 514288
rect 64350 514232 64418 514288
rect 64474 514232 64496 514288
rect 64024 514164 64496 514232
rect 64024 514108 64046 514164
rect 64102 514108 64170 514164
rect 64226 514108 64294 514164
rect 64350 514108 64418 514164
rect 64474 514108 64496 514164
rect 64024 514040 64496 514108
rect 64024 513984 64046 514040
rect 64102 513984 64170 514040
rect 64226 513984 64294 514040
rect 64350 513984 64418 514040
rect 64474 513984 64496 514040
rect 64024 513916 64496 513984
rect 64024 513860 64046 513916
rect 64102 513860 64170 513916
rect 64226 513860 64294 513916
rect 64350 513860 64418 513916
rect 64474 513860 64496 513916
rect 64024 513826 64496 513860
rect 64520 514412 64992 514446
rect 64520 514356 64542 514412
rect 64598 514356 64666 514412
rect 64722 514356 64790 514412
rect 64846 514356 64914 514412
rect 64970 514356 64992 514412
rect 64520 514288 64992 514356
rect 64520 514232 64542 514288
rect 64598 514232 64666 514288
rect 64722 514232 64790 514288
rect 64846 514232 64914 514288
rect 64970 514232 64992 514288
rect 64520 514164 64992 514232
rect 64520 514108 64542 514164
rect 64598 514108 64666 514164
rect 64722 514108 64790 514164
rect 64846 514108 64914 514164
rect 64970 514108 64992 514164
rect 64520 514040 64992 514108
rect 64520 513984 64542 514040
rect 64598 513984 64666 514040
rect 64722 513984 64790 514040
rect 64846 513984 64914 514040
rect 64970 513984 64992 514040
rect 64520 513916 64992 513984
rect 64520 513860 64542 513916
rect 64598 513860 64666 513916
rect 64722 513860 64790 513916
rect 64846 513860 64914 513916
rect 64970 513860 64992 513916
rect 64520 513826 64992 513860
rect 65016 514412 65488 514446
rect 65016 514356 65038 514412
rect 65094 514356 65162 514412
rect 65218 514356 65286 514412
rect 65342 514356 65410 514412
rect 65466 514356 65488 514412
rect 65016 514288 65488 514356
rect 65016 514232 65038 514288
rect 65094 514232 65162 514288
rect 65218 514232 65286 514288
rect 65342 514232 65410 514288
rect 65466 514232 65488 514288
rect 65016 514164 65488 514232
rect 65016 514108 65038 514164
rect 65094 514108 65162 514164
rect 65218 514108 65286 514164
rect 65342 514108 65410 514164
rect 65466 514108 65488 514164
rect 65016 514040 65488 514108
rect 65016 513984 65038 514040
rect 65094 513984 65162 514040
rect 65218 513984 65286 514040
rect 65342 513984 65410 514040
rect 65466 513984 65488 514040
rect 65016 513916 65488 513984
rect 65016 513860 65038 513916
rect 65094 513860 65162 513916
rect 65218 513860 65286 513916
rect 65342 513860 65410 513916
rect 65466 513860 65488 513916
rect 65016 513826 65488 513860
rect 65512 514412 65984 514446
rect 65512 514356 65534 514412
rect 65590 514356 65658 514412
rect 65714 514356 65782 514412
rect 65838 514356 65906 514412
rect 65962 514356 65984 514412
rect 65512 514288 65984 514356
rect 65512 514232 65534 514288
rect 65590 514232 65658 514288
rect 65714 514232 65782 514288
rect 65838 514232 65906 514288
rect 65962 514232 65984 514288
rect 65512 514164 65984 514232
rect 65512 514108 65534 514164
rect 65590 514108 65658 514164
rect 65714 514108 65782 514164
rect 65838 514108 65906 514164
rect 65962 514108 65984 514164
rect 65512 514040 65984 514108
rect 65512 513984 65534 514040
rect 65590 513984 65658 514040
rect 65714 513984 65782 514040
rect 65838 513984 65906 514040
rect 65962 513984 65984 514040
rect 65512 513916 65984 513984
rect 65512 513860 65534 513916
rect 65590 513860 65658 513916
rect 65714 513860 65782 513916
rect 65838 513860 65906 513916
rect 65962 513860 65984 513916
rect 65512 513826 65984 513860
rect 66008 514412 66480 514446
rect 66008 514356 66030 514412
rect 66086 514356 66154 514412
rect 66210 514356 66278 514412
rect 66334 514356 66402 514412
rect 66458 514356 66480 514412
rect 66008 514288 66480 514356
rect 66008 514232 66030 514288
rect 66086 514232 66154 514288
rect 66210 514232 66278 514288
rect 66334 514232 66402 514288
rect 66458 514232 66480 514288
rect 66008 514164 66480 514232
rect 66008 514108 66030 514164
rect 66086 514108 66154 514164
rect 66210 514108 66278 514164
rect 66334 514108 66402 514164
rect 66458 514108 66480 514164
rect 66008 514040 66480 514108
rect 66008 513984 66030 514040
rect 66086 513984 66154 514040
rect 66210 513984 66278 514040
rect 66334 513984 66402 514040
rect 66458 513984 66480 514040
rect 66008 513916 66480 513984
rect 66008 513860 66030 513916
rect 66086 513860 66154 513916
rect 66210 513860 66278 513916
rect 66334 513860 66402 513916
rect 66458 513860 66480 513916
rect 66008 513826 66480 513860
rect 90060 508435 100140 508446
rect 90060 508379 90112 508435
rect 90168 508379 90236 508435
rect 90292 508379 90360 508435
rect 90416 508379 90484 508435
rect 90540 508379 90608 508435
rect 90664 508379 90732 508435
rect 90788 508379 90856 508435
rect 90912 508379 90980 508435
rect 91036 508379 91104 508435
rect 91160 508379 91228 508435
rect 91284 508379 91352 508435
rect 91408 508379 91476 508435
rect 91532 508379 91600 508435
rect 91656 508379 91724 508435
rect 91780 508379 91848 508435
rect 91904 508379 91972 508435
rect 92028 508379 92096 508435
rect 92152 508379 92220 508435
rect 92276 508379 92344 508435
rect 92400 508379 92468 508435
rect 92524 508379 92592 508435
rect 92648 508379 92716 508435
rect 92772 508379 92840 508435
rect 92896 508379 92964 508435
rect 93020 508379 93088 508435
rect 93144 508379 93212 508435
rect 93268 508379 93336 508435
rect 93392 508379 93460 508435
rect 93516 508379 93584 508435
rect 93640 508379 93708 508435
rect 93764 508379 93832 508435
rect 93888 508379 93956 508435
rect 94012 508379 94080 508435
rect 94136 508379 94204 508435
rect 94260 508379 94328 508435
rect 94384 508379 94452 508435
rect 94508 508379 94576 508435
rect 94632 508379 94700 508435
rect 94756 508379 94824 508435
rect 94880 508379 94948 508435
rect 95004 508379 95072 508435
rect 95128 508379 95196 508435
rect 95252 508379 95320 508435
rect 95376 508379 95444 508435
rect 95500 508379 95568 508435
rect 95624 508379 95692 508435
rect 95748 508379 95816 508435
rect 95872 508379 95940 508435
rect 95996 508379 96064 508435
rect 96120 508379 96188 508435
rect 96244 508379 96312 508435
rect 96368 508379 96436 508435
rect 96492 508379 96560 508435
rect 96616 508379 96684 508435
rect 96740 508379 96808 508435
rect 96864 508379 96932 508435
rect 96988 508379 97056 508435
rect 97112 508379 97180 508435
rect 97236 508379 97304 508435
rect 97360 508379 97428 508435
rect 97484 508379 97552 508435
rect 97608 508379 97676 508435
rect 97732 508379 97800 508435
rect 97856 508379 97924 508435
rect 97980 508379 98048 508435
rect 98104 508379 98172 508435
rect 98228 508379 98296 508435
rect 98352 508379 98420 508435
rect 98476 508379 98544 508435
rect 98600 508379 98668 508435
rect 98724 508379 98792 508435
rect 98848 508379 98916 508435
rect 98972 508379 99040 508435
rect 99096 508379 99164 508435
rect 99220 508379 99288 508435
rect 99344 508379 99412 508435
rect 99468 508379 99536 508435
rect 99592 508379 99660 508435
rect 99716 508379 99784 508435
rect 99840 508379 99908 508435
rect 99964 508379 100032 508435
rect 100088 508379 100140 508435
rect 90060 508311 100140 508379
rect 90060 508255 90112 508311
rect 90168 508255 90236 508311
rect 90292 508255 90360 508311
rect 90416 508255 90484 508311
rect 90540 508255 90608 508311
rect 90664 508255 90732 508311
rect 90788 508255 90856 508311
rect 90912 508255 90980 508311
rect 91036 508255 91104 508311
rect 91160 508255 91228 508311
rect 91284 508255 91352 508311
rect 91408 508255 91476 508311
rect 91532 508255 91600 508311
rect 91656 508255 91724 508311
rect 91780 508255 91848 508311
rect 91904 508255 91972 508311
rect 92028 508255 92096 508311
rect 92152 508255 92220 508311
rect 92276 508255 92344 508311
rect 92400 508255 92468 508311
rect 92524 508255 92592 508311
rect 92648 508255 92716 508311
rect 92772 508255 92840 508311
rect 92896 508255 92964 508311
rect 93020 508255 93088 508311
rect 93144 508255 93212 508311
rect 93268 508255 93336 508311
rect 93392 508255 93460 508311
rect 93516 508255 93584 508311
rect 93640 508255 93708 508311
rect 93764 508255 93832 508311
rect 93888 508255 93956 508311
rect 94012 508255 94080 508311
rect 94136 508255 94204 508311
rect 94260 508255 94328 508311
rect 94384 508255 94452 508311
rect 94508 508255 94576 508311
rect 94632 508255 94700 508311
rect 94756 508255 94824 508311
rect 94880 508255 94948 508311
rect 95004 508255 95072 508311
rect 95128 508255 95196 508311
rect 95252 508255 95320 508311
rect 95376 508255 95444 508311
rect 95500 508255 95568 508311
rect 95624 508255 95692 508311
rect 95748 508255 95816 508311
rect 95872 508255 95940 508311
rect 95996 508255 96064 508311
rect 96120 508255 96188 508311
rect 96244 508255 96312 508311
rect 96368 508255 96436 508311
rect 96492 508255 96560 508311
rect 96616 508255 96684 508311
rect 96740 508255 96808 508311
rect 96864 508255 96932 508311
rect 96988 508255 97056 508311
rect 97112 508255 97180 508311
rect 97236 508255 97304 508311
rect 97360 508255 97428 508311
rect 97484 508255 97552 508311
rect 97608 508255 97676 508311
rect 97732 508255 97800 508311
rect 97856 508255 97924 508311
rect 97980 508255 98048 508311
rect 98104 508255 98172 508311
rect 98228 508255 98296 508311
rect 98352 508255 98420 508311
rect 98476 508255 98544 508311
rect 98600 508255 98668 508311
rect 98724 508255 98792 508311
rect 98848 508255 98916 508311
rect 98972 508255 99040 508311
rect 99096 508255 99164 508311
rect 99220 508255 99288 508311
rect 99344 508255 99412 508311
rect 99468 508255 99536 508311
rect 99592 508255 99660 508311
rect 99716 508255 99784 508311
rect 99840 508255 99908 508311
rect 99964 508255 100032 508311
rect 100088 508255 100140 508311
rect 90060 508187 100140 508255
rect 90060 508131 90112 508187
rect 90168 508131 90236 508187
rect 90292 508131 90360 508187
rect 90416 508131 90484 508187
rect 90540 508131 90608 508187
rect 90664 508131 90732 508187
rect 90788 508131 90856 508187
rect 90912 508131 90980 508187
rect 91036 508131 91104 508187
rect 91160 508131 91228 508187
rect 91284 508131 91352 508187
rect 91408 508131 91476 508187
rect 91532 508131 91600 508187
rect 91656 508131 91724 508187
rect 91780 508131 91848 508187
rect 91904 508131 91972 508187
rect 92028 508131 92096 508187
rect 92152 508131 92220 508187
rect 92276 508131 92344 508187
rect 92400 508131 92468 508187
rect 92524 508131 92592 508187
rect 92648 508131 92716 508187
rect 92772 508131 92840 508187
rect 92896 508131 92964 508187
rect 93020 508131 93088 508187
rect 93144 508131 93212 508187
rect 93268 508131 93336 508187
rect 93392 508131 93460 508187
rect 93516 508131 93584 508187
rect 93640 508131 93708 508187
rect 93764 508131 93832 508187
rect 93888 508131 93956 508187
rect 94012 508131 94080 508187
rect 94136 508131 94204 508187
rect 94260 508131 94328 508187
rect 94384 508131 94452 508187
rect 94508 508131 94576 508187
rect 94632 508131 94700 508187
rect 94756 508131 94824 508187
rect 94880 508131 94948 508187
rect 95004 508131 95072 508187
rect 95128 508131 95196 508187
rect 95252 508131 95320 508187
rect 95376 508131 95444 508187
rect 95500 508131 95568 508187
rect 95624 508131 95692 508187
rect 95748 508131 95816 508187
rect 95872 508131 95940 508187
rect 95996 508131 96064 508187
rect 96120 508131 96188 508187
rect 96244 508131 96312 508187
rect 96368 508131 96436 508187
rect 96492 508131 96560 508187
rect 96616 508131 96684 508187
rect 96740 508131 96808 508187
rect 96864 508131 96932 508187
rect 96988 508131 97056 508187
rect 97112 508131 97180 508187
rect 97236 508131 97304 508187
rect 97360 508131 97428 508187
rect 97484 508131 97552 508187
rect 97608 508131 97676 508187
rect 97732 508131 97800 508187
rect 97856 508131 97924 508187
rect 97980 508131 98048 508187
rect 98104 508131 98172 508187
rect 98228 508131 98296 508187
rect 98352 508131 98420 508187
rect 98476 508131 98544 508187
rect 98600 508131 98668 508187
rect 98724 508131 98792 508187
rect 98848 508131 98916 508187
rect 98972 508131 99040 508187
rect 99096 508131 99164 508187
rect 99220 508131 99288 508187
rect 99344 508131 99412 508187
rect 99468 508131 99536 508187
rect 99592 508131 99660 508187
rect 99716 508131 99784 508187
rect 99840 508131 99908 508187
rect 99964 508131 100032 508187
rect 100088 508131 100140 508187
rect 90060 508120 100140 508131
rect 39858 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 40478 496350
rect 39858 496226 40478 496294
rect 39858 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 40478 496226
rect 39858 496102 40478 496170
rect 39858 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 40478 496102
rect 39858 495978 40478 496046
rect 39858 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 40478 495978
rect 39858 478350 40478 495922
rect 63420 496212 63496 496240
rect 63420 496156 63430 496212
rect 63486 496156 63496 496212
rect 63420 496088 63496 496156
rect 63420 496032 63430 496088
rect 63486 496032 63496 496088
rect 63420 495964 63496 496032
rect 63420 495908 63430 495964
rect 63486 495908 63496 495964
rect 63420 495880 63496 495908
rect 63544 496212 63992 496240
rect 63544 496156 63554 496212
rect 63610 496156 63678 496212
rect 63734 496156 63802 496212
rect 63858 496156 63926 496212
rect 63982 496156 63992 496212
rect 63544 496088 63992 496156
rect 63544 496032 63554 496088
rect 63610 496032 63678 496088
rect 63734 496032 63802 496088
rect 63858 496032 63926 496088
rect 63982 496032 63992 496088
rect 63544 495964 63992 496032
rect 63544 495908 63554 495964
rect 63610 495908 63678 495964
rect 63734 495908 63802 495964
rect 63858 495908 63926 495964
rect 63982 495908 63992 495964
rect 63544 495880 63992 495908
rect 64040 496212 64488 496240
rect 64040 496156 64050 496212
rect 64106 496156 64174 496212
rect 64230 496156 64298 496212
rect 64354 496156 64422 496212
rect 64478 496156 64488 496212
rect 64040 496088 64488 496156
rect 64040 496032 64050 496088
rect 64106 496032 64174 496088
rect 64230 496032 64298 496088
rect 64354 496032 64422 496088
rect 64478 496032 64488 496088
rect 64040 495964 64488 496032
rect 64040 495908 64050 495964
rect 64106 495908 64174 495964
rect 64230 495908 64298 495964
rect 64354 495908 64422 495964
rect 64478 495908 64488 495964
rect 64040 495880 64488 495908
rect 64536 496212 64984 496240
rect 64536 496156 64546 496212
rect 64602 496156 64670 496212
rect 64726 496156 64794 496212
rect 64850 496156 64918 496212
rect 64974 496156 64984 496212
rect 64536 496088 64984 496156
rect 64536 496032 64546 496088
rect 64602 496032 64670 496088
rect 64726 496032 64794 496088
rect 64850 496032 64918 496088
rect 64974 496032 64984 496088
rect 64536 495964 64984 496032
rect 64536 495908 64546 495964
rect 64602 495908 64670 495964
rect 64726 495908 64794 495964
rect 64850 495908 64918 495964
rect 64974 495908 64984 495964
rect 64536 495880 64984 495908
rect 65032 496212 65480 496240
rect 65032 496156 65042 496212
rect 65098 496156 65166 496212
rect 65222 496156 65290 496212
rect 65346 496156 65414 496212
rect 65470 496156 65480 496212
rect 65032 496088 65480 496156
rect 65032 496032 65042 496088
rect 65098 496032 65166 496088
rect 65222 496032 65290 496088
rect 65346 496032 65414 496088
rect 65470 496032 65480 496088
rect 65032 495964 65480 496032
rect 65032 495908 65042 495964
rect 65098 495908 65166 495964
rect 65222 495908 65290 495964
rect 65346 495908 65414 495964
rect 65470 495908 65480 495964
rect 65032 495880 65480 495908
rect 65528 496212 65976 496240
rect 65528 496156 65538 496212
rect 65594 496156 65662 496212
rect 65718 496156 65786 496212
rect 65842 496156 65910 496212
rect 65966 496156 65976 496212
rect 65528 496088 65976 496156
rect 65528 496032 65538 496088
rect 65594 496032 65662 496088
rect 65718 496032 65786 496088
rect 65842 496032 65910 496088
rect 65966 496032 65976 496088
rect 65528 495964 65976 496032
rect 65528 495908 65538 495964
rect 65594 495908 65662 495964
rect 65718 495908 65786 495964
rect 65842 495908 65910 495964
rect 65966 495908 65976 495964
rect 65528 495880 65976 495908
rect 66024 496212 66472 496240
rect 66024 496156 66034 496212
rect 66090 496156 66158 496212
rect 66214 496156 66282 496212
rect 66338 496156 66406 496212
rect 66462 496156 66472 496212
rect 66024 496088 66472 496156
rect 66024 496032 66034 496088
rect 66090 496032 66158 496088
rect 66214 496032 66282 496088
rect 66338 496032 66406 496088
rect 66462 496032 66472 496088
rect 66024 495964 66472 496032
rect 66024 495908 66034 495964
rect 66090 495908 66158 495964
rect 66214 495908 66282 495964
rect 66338 495908 66406 495964
rect 66462 495908 66472 495964
rect 66024 495880 66472 495908
rect 66520 496212 66968 496240
rect 66520 496156 66530 496212
rect 66586 496156 66654 496212
rect 66710 496156 66778 496212
rect 66834 496156 66902 496212
rect 66958 496156 66968 496212
rect 66520 496088 66968 496156
rect 66520 496032 66530 496088
rect 66586 496032 66654 496088
rect 66710 496032 66778 496088
rect 66834 496032 66902 496088
rect 66958 496032 66968 496088
rect 66520 495964 66968 496032
rect 66520 495908 66530 495964
rect 66586 495908 66654 495964
rect 66710 495908 66778 495964
rect 66834 495908 66902 495964
rect 66958 495908 66968 495964
rect 66520 495880 66968 495908
rect 67016 496212 67464 496240
rect 67016 496156 67026 496212
rect 67082 496156 67150 496212
rect 67206 496156 67274 496212
rect 67330 496156 67398 496212
rect 67454 496156 67464 496212
rect 67016 496088 67464 496156
rect 67016 496032 67026 496088
rect 67082 496032 67150 496088
rect 67206 496032 67274 496088
rect 67330 496032 67398 496088
rect 67454 496032 67464 496088
rect 67016 495964 67464 496032
rect 67016 495908 67026 495964
rect 67082 495908 67150 495964
rect 67206 495908 67274 495964
rect 67330 495908 67398 495964
rect 67454 495908 67464 495964
rect 67016 495880 67464 495908
rect 67512 496212 67960 496240
rect 67512 496156 67522 496212
rect 67578 496156 67646 496212
rect 67702 496156 67770 496212
rect 67826 496156 67894 496212
rect 67950 496156 67960 496212
rect 67512 496088 67960 496156
rect 67512 496032 67522 496088
rect 67578 496032 67646 496088
rect 67702 496032 67770 496088
rect 67826 496032 67894 496088
rect 67950 496032 67960 496088
rect 67512 495964 67960 496032
rect 67512 495908 67522 495964
rect 67578 495908 67646 495964
rect 67702 495908 67770 495964
rect 67826 495908 67894 495964
rect 67950 495908 67960 495964
rect 67512 495880 67960 495908
rect 68008 496212 68456 496240
rect 68008 496156 68018 496212
rect 68074 496156 68142 496212
rect 68198 496156 68266 496212
rect 68322 496156 68390 496212
rect 68446 496156 68456 496212
rect 68008 496088 68456 496156
rect 68008 496032 68018 496088
rect 68074 496032 68142 496088
rect 68198 496032 68266 496088
rect 68322 496032 68390 496088
rect 68446 496032 68456 496088
rect 68008 495964 68456 496032
rect 68008 495908 68018 495964
rect 68074 495908 68142 495964
rect 68198 495908 68266 495964
rect 68322 495908 68390 495964
rect 68446 495908 68456 495964
rect 68008 495880 68456 495908
rect 68504 496212 68952 496240
rect 68504 496156 68514 496212
rect 68570 496156 68638 496212
rect 68694 496156 68762 496212
rect 68818 496156 68886 496212
rect 68942 496156 68952 496212
rect 68504 496088 68952 496156
rect 68504 496032 68514 496088
rect 68570 496032 68638 496088
rect 68694 496032 68762 496088
rect 68818 496032 68886 496088
rect 68942 496032 68952 496088
rect 68504 495964 68952 496032
rect 68504 495908 68514 495964
rect 68570 495908 68638 495964
rect 68694 495908 68762 495964
rect 68818 495908 68886 495964
rect 68942 495908 68952 495964
rect 68504 495880 68952 495908
rect 69000 496212 69448 496240
rect 69000 496156 69010 496212
rect 69066 496156 69134 496212
rect 69190 496156 69258 496212
rect 69314 496156 69382 496212
rect 69438 496156 69448 496212
rect 69000 496088 69448 496156
rect 69000 496032 69010 496088
rect 69066 496032 69134 496088
rect 69190 496032 69258 496088
rect 69314 496032 69382 496088
rect 69438 496032 69448 496088
rect 69000 495964 69448 496032
rect 69000 495908 69010 495964
rect 69066 495908 69134 495964
rect 69190 495908 69258 495964
rect 69314 495908 69382 495964
rect 69438 495908 69448 495964
rect 69000 495880 69448 495908
rect 69496 496212 69944 496240
rect 69496 496156 69506 496212
rect 69562 496156 69630 496212
rect 69686 496156 69754 496212
rect 69810 496156 69878 496212
rect 69934 496156 69944 496212
rect 69496 496088 69944 496156
rect 69496 496032 69506 496088
rect 69562 496032 69630 496088
rect 69686 496032 69754 496088
rect 69810 496032 69878 496088
rect 69934 496032 69944 496088
rect 69496 495964 69944 496032
rect 69496 495908 69506 495964
rect 69562 495908 69630 495964
rect 69686 495908 69754 495964
rect 69810 495908 69878 495964
rect 69934 495908 69944 495964
rect 69496 495880 69944 495908
rect 69992 496212 70440 496240
rect 69992 496156 70002 496212
rect 70058 496156 70126 496212
rect 70182 496156 70250 496212
rect 70306 496156 70374 496212
rect 70430 496156 70440 496212
rect 69992 496088 70440 496156
rect 69992 496032 70002 496088
rect 70058 496032 70126 496088
rect 70182 496032 70250 496088
rect 70306 496032 70374 496088
rect 70430 496032 70440 496088
rect 69992 495964 70440 496032
rect 69992 495908 70002 495964
rect 70058 495908 70126 495964
rect 70182 495908 70250 495964
rect 70306 495908 70374 495964
rect 70430 495908 70440 495964
rect 69992 495880 70440 495908
rect 85200 490272 88800 490300
rect 85200 490216 85236 490272
rect 85292 490216 85360 490272
rect 85416 490216 85484 490272
rect 85540 490216 85608 490272
rect 85664 490216 85732 490272
rect 85788 490216 85856 490272
rect 85912 490216 85980 490272
rect 86036 490216 86104 490272
rect 86160 490216 86228 490272
rect 86284 490216 86352 490272
rect 86408 490216 86476 490272
rect 86532 490216 86600 490272
rect 86656 490216 86724 490272
rect 86780 490216 86848 490272
rect 86904 490216 86972 490272
rect 87028 490216 87096 490272
rect 87152 490216 87220 490272
rect 87276 490216 87344 490272
rect 87400 490216 87468 490272
rect 87524 490216 87592 490272
rect 87648 490216 87716 490272
rect 87772 490216 87840 490272
rect 87896 490216 87964 490272
rect 88020 490216 88088 490272
rect 88144 490216 88212 490272
rect 88268 490216 88336 490272
rect 88392 490216 88460 490272
rect 88516 490216 88584 490272
rect 88640 490216 88708 490272
rect 88764 490216 88800 490272
rect 85200 490148 88800 490216
rect 85200 490092 85236 490148
rect 85292 490092 85360 490148
rect 85416 490092 85484 490148
rect 85540 490092 85608 490148
rect 85664 490092 85732 490148
rect 85788 490092 85856 490148
rect 85912 490092 85980 490148
rect 86036 490092 86104 490148
rect 86160 490092 86228 490148
rect 86284 490092 86352 490148
rect 86408 490092 86476 490148
rect 86532 490092 86600 490148
rect 86656 490092 86724 490148
rect 86780 490092 86848 490148
rect 86904 490092 86972 490148
rect 87028 490092 87096 490148
rect 87152 490092 87220 490148
rect 87276 490092 87344 490148
rect 87400 490092 87468 490148
rect 87524 490092 87592 490148
rect 87648 490092 87716 490148
rect 87772 490092 87840 490148
rect 87896 490092 87964 490148
rect 88020 490092 88088 490148
rect 88144 490092 88212 490148
rect 88268 490092 88336 490148
rect 88392 490092 88460 490148
rect 88516 490092 88584 490148
rect 88640 490092 88708 490148
rect 88764 490092 88800 490148
rect 85200 490024 88800 490092
rect 85200 489968 85236 490024
rect 85292 489968 85360 490024
rect 85416 489968 85484 490024
rect 85540 489968 85608 490024
rect 85664 489968 85732 490024
rect 85788 489968 85856 490024
rect 85912 489968 85980 490024
rect 86036 489968 86104 490024
rect 86160 489968 86228 490024
rect 86284 489968 86352 490024
rect 86408 489968 86476 490024
rect 86532 489968 86600 490024
rect 86656 489968 86724 490024
rect 86780 489968 86848 490024
rect 86904 489968 86972 490024
rect 87028 489968 87096 490024
rect 87152 489968 87220 490024
rect 87276 489968 87344 490024
rect 87400 489968 87468 490024
rect 87524 489968 87592 490024
rect 87648 489968 87716 490024
rect 87772 489968 87840 490024
rect 87896 489968 87964 490024
rect 88020 489968 88088 490024
rect 88144 489968 88212 490024
rect 88268 489968 88336 490024
rect 88392 489968 88460 490024
rect 88516 489968 88584 490024
rect 88640 489968 88708 490024
rect 88764 489968 88800 490024
rect 85200 489940 88800 489968
rect 39858 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 40478 478350
rect 39858 478226 40478 478294
rect 39858 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 40478 478226
rect 39858 478102 40478 478170
rect 39858 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 40478 478102
rect 39858 477978 40478 478046
rect 39858 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 40478 477978
rect 39858 460350 40478 477922
rect 39858 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 40478 460350
rect 39858 460226 40478 460294
rect 39858 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 40478 460226
rect 39858 460102 40478 460170
rect 39858 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 40478 460102
rect 39858 459978 40478 460046
rect 39858 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 40478 459978
rect 39858 442350 40478 459922
rect 39858 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 40478 442350
rect 39858 442226 40478 442294
rect 39858 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 40478 442226
rect 39858 442102 40478 442170
rect 39858 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 40478 442102
rect 39858 441978 40478 442046
rect 39858 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 40478 441978
rect 39858 424350 40478 441922
rect 39858 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 40478 424350
rect 39858 424226 40478 424294
rect 39858 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 40478 424226
rect 39858 424102 40478 424170
rect 39858 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 40478 424102
rect 39858 423978 40478 424046
rect 39858 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 40478 423978
rect 39858 406350 40478 423922
rect 66858 472350 67478 486928
rect 66858 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 67478 472350
rect 66858 472226 67478 472294
rect 66858 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 67478 472226
rect 66858 472102 67478 472170
rect 66858 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 67478 472102
rect 66858 471978 67478 472046
rect 66858 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 67478 471978
rect 66858 454350 67478 471922
rect 66858 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 67478 454350
rect 66858 454226 67478 454294
rect 66858 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 67478 454226
rect 66858 454102 67478 454170
rect 66858 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 67478 454102
rect 66858 453978 67478 454046
rect 66858 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 67478 453978
rect 66858 436350 67478 453922
rect 66858 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 67478 436350
rect 66858 436226 67478 436294
rect 66858 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 67478 436226
rect 66858 436102 67478 436170
rect 66858 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 67478 436102
rect 66858 435978 67478 436046
rect 66858 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 67478 435978
rect 66858 418350 67478 435922
rect 66858 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 67478 418350
rect 66858 418226 67478 418294
rect 66858 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 67478 418226
rect 66858 418102 67478 418170
rect 66858 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 67478 418102
rect 66858 417978 67478 418046
rect 66858 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 67478 417978
rect 61852 413364 61908 413374
rect 61852 408268 61908 413308
rect 66858 412556 67478 417922
rect 70578 478350 71198 482968
rect 70578 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 71198 478350
rect 70578 478226 71198 478294
rect 80880 478358 81420 478420
rect 80880 478302 80936 478358
rect 80992 478302 81060 478358
rect 81116 478302 81184 478358
rect 81240 478302 81308 478358
rect 81364 478302 81420 478358
rect 80880 478240 81420 478302
rect 70578 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 71198 478226
rect 70578 478102 71198 478170
rect 70578 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 71198 478102
rect 70578 477978 71198 478046
rect 70578 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 71198 477978
rect 70578 460350 71198 477922
rect 70578 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 71198 460350
rect 70578 460226 71198 460294
rect 70578 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 71198 460226
rect 70578 460102 71198 460170
rect 70578 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 71198 460102
rect 70578 459978 71198 460046
rect 70578 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 71198 459978
rect 70578 442350 71198 459922
rect 70578 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 71198 442350
rect 70578 442226 71198 442294
rect 70578 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 71198 442226
rect 70578 442102 71198 442170
rect 70578 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 71198 442102
rect 70578 441978 71198 442046
rect 70578 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 71198 441978
rect 70578 424350 71198 441922
rect 70578 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 71198 424350
rect 70578 424226 71198 424294
rect 70578 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 71198 424226
rect 70578 424102 71198 424170
rect 70578 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 71198 424102
rect 70578 423978 71198 424046
rect 70578 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 71198 423978
rect 70578 410574 71198 423922
rect 97578 472350 98198 472888
rect 97578 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 98198 472350
rect 97578 472226 98198 472294
rect 97578 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 98198 472226
rect 97578 472102 98198 472170
rect 97578 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 98198 472102
rect 97578 471978 98198 472046
rect 97578 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 98198 471978
rect 97578 454350 98198 471922
rect 97578 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 98198 454350
rect 97578 454226 98198 454294
rect 97578 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 98198 454226
rect 97578 454102 98198 454170
rect 97578 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 98198 454102
rect 97578 453978 98198 454046
rect 97578 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 98198 453978
rect 97578 436350 98198 453922
rect 97578 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 98198 436350
rect 97578 436226 98198 436294
rect 97578 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 98198 436226
rect 97578 436102 98198 436170
rect 97578 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 98198 436102
rect 97578 435978 98198 436046
rect 97578 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 98198 435978
rect 97578 418350 98198 435922
rect 97578 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 98198 418350
rect 97578 418226 98198 418294
rect 97578 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 98198 418226
rect 97578 418102 98198 418170
rect 97578 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 98198 418102
rect 97578 417978 98198 418046
rect 97578 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 98198 417978
rect 83916 416818 83972 416828
rect 83916 409780 83972 416762
rect 83916 409714 83972 409724
rect 61852 408212 62132 408268
rect 39858 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 40478 406350
rect 39858 406226 40478 406294
rect 39858 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 40478 406226
rect 39858 406102 40478 406170
rect 39858 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 40478 406102
rect 39858 405978 40478 406046
rect 39858 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 40478 405978
rect 39858 388350 40478 405922
rect 62076 390538 62132 408212
rect 66504 406350 66824 406384
rect 66504 406294 66574 406350
rect 66630 406294 66698 406350
rect 66754 406294 66824 406350
rect 66504 406226 66824 406294
rect 66504 406170 66574 406226
rect 66630 406170 66698 406226
rect 66754 406170 66824 406226
rect 66504 406102 66824 406170
rect 66504 406046 66574 406102
rect 66630 406046 66698 406102
rect 66754 406046 66824 406102
rect 66504 405978 66824 406046
rect 66504 405922 66574 405978
rect 66630 405922 66698 405978
rect 66754 405922 66824 405978
rect 66504 405888 66824 405922
rect 71824 406350 72144 406384
rect 71824 406294 71894 406350
rect 71950 406294 72018 406350
rect 72074 406294 72144 406350
rect 71824 406226 72144 406294
rect 71824 406170 71894 406226
rect 71950 406170 72018 406226
rect 72074 406170 72144 406226
rect 71824 406102 72144 406170
rect 71824 406046 71894 406102
rect 71950 406046 72018 406102
rect 72074 406046 72144 406102
rect 71824 405978 72144 406046
rect 71824 405922 71894 405978
rect 71950 405922 72018 405978
rect 72074 405922 72144 405978
rect 71824 405888 72144 405922
rect 77144 406350 77464 406384
rect 77144 406294 77214 406350
rect 77270 406294 77338 406350
rect 77394 406294 77464 406350
rect 77144 406226 77464 406294
rect 77144 406170 77214 406226
rect 77270 406170 77338 406226
rect 77394 406170 77464 406226
rect 77144 406102 77464 406170
rect 77144 406046 77214 406102
rect 77270 406046 77338 406102
rect 77394 406046 77464 406102
rect 77144 405978 77464 406046
rect 77144 405922 77214 405978
rect 77270 405922 77338 405978
rect 77394 405922 77464 405978
rect 77144 405888 77464 405922
rect 82464 406350 82784 406384
rect 82464 406294 82534 406350
rect 82590 406294 82658 406350
rect 82714 406294 82784 406350
rect 82464 406226 82784 406294
rect 82464 406170 82534 406226
rect 82590 406170 82658 406226
rect 82714 406170 82784 406226
rect 82464 406102 82784 406170
rect 82464 406046 82534 406102
rect 82590 406046 82658 406102
rect 82714 406046 82784 406102
rect 82464 405978 82784 406046
rect 82464 405922 82534 405978
rect 82590 405922 82658 405978
rect 82714 405922 82784 405978
rect 82464 405888 82784 405922
rect 92428 404964 92484 404974
rect 89964 403284 90020 403294
rect 63844 400350 64164 400384
rect 63844 400294 63914 400350
rect 63970 400294 64038 400350
rect 64094 400294 64164 400350
rect 63844 400226 64164 400294
rect 63844 400170 63914 400226
rect 63970 400170 64038 400226
rect 64094 400170 64164 400226
rect 63844 400102 64164 400170
rect 63844 400046 63914 400102
rect 63970 400046 64038 400102
rect 64094 400046 64164 400102
rect 63844 399978 64164 400046
rect 63844 399922 63914 399978
rect 63970 399922 64038 399978
rect 64094 399922 64164 399978
rect 63844 399888 64164 399922
rect 69164 400350 69484 400384
rect 69164 400294 69234 400350
rect 69290 400294 69358 400350
rect 69414 400294 69484 400350
rect 69164 400226 69484 400294
rect 69164 400170 69234 400226
rect 69290 400170 69358 400226
rect 69414 400170 69484 400226
rect 69164 400102 69484 400170
rect 69164 400046 69234 400102
rect 69290 400046 69358 400102
rect 69414 400046 69484 400102
rect 69164 399978 69484 400046
rect 69164 399922 69234 399978
rect 69290 399922 69358 399978
rect 69414 399922 69484 399978
rect 69164 399888 69484 399922
rect 74484 400350 74804 400384
rect 74484 400294 74554 400350
rect 74610 400294 74678 400350
rect 74734 400294 74804 400350
rect 74484 400226 74804 400294
rect 74484 400170 74554 400226
rect 74610 400170 74678 400226
rect 74734 400170 74804 400226
rect 74484 400102 74804 400170
rect 74484 400046 74554 400102
rect 74610 400046 74678 400102
rect 74734 400046 74804 400102
rect 74484 399978 74804 400046
rect 74484 399922 74554 399978
rect 74610 399922 74678 399978
rect 74734 399922 74804 399978
rect 74484 399888 74804 399922
rect 79804 400350 80124 400384
rect 79804 400294 79874 400350
rect 79930 400294 79998 400350
rect 80054 400294 80124 400350
rect 79804 400226 80124 400294
rect 79804 400170 79874 400226
rect 79930 400170 79998 400226
rect 80054 400170 80124 400226
rect 79804 400102 80124 400170
rect 79804 400046 79874 400102
rect 79930 400046 79998 400102
rect 80054 400046 80124 400102
rect 79804 399978 80124 400046
rect 79804 399922 79874 399978
rect 79930 399922 79998 399978
rect 80054 399922 80124 399978
rect 79804 399888 80124 399922
rect 89852 400372 89908 400382
rect 62076 390472 62132 390482
rect 39858 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 40478 388350
rect 39858 388226 40478 388294
rect 39858 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 40478 388226
rect 39858 388102 40478 388170
rect 39858 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 40478 388102
rect 39858 387978 40478 388046
rect 39858 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 40478 387978
rect 36138 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 36758 364350
rect 36138 364226 36758 364294
rect 36138 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 36758 364226
rect 36138 364102 36758 364170
rect 36138 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 36758 364102
rect 36138 363978 36758 364046
rect 36138 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 36758 363978
rect 36138 346350 36758 363922
rect 36138 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 36758 346350
rect 36138 346226 36758 346294
rect 36138 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 36758 346226
rect 36138 346102 36758 346170
rect 36138 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 36758 346102
rect 36138 345978 36758 346046
rect 36138 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 36758 345978
rect 36138 328350 36758 345922
rect 36138 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 36758 328350
rect 36138 328226 36758 328294
rect 36138 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 36758 328226
rect 36138 328102 36758 328170
rect 36138 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 36758 328102
rect 36138 327978 36758 328046
rect 36138 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 36758 327978
rect 36138 310350 36758 327922
rect 36138 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 36758 310350
rect 36138 310226 36758 310294
rect 36138 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 36758 310226
rect 36138 310102 36758 310170
rect 36138 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 36758 310102
rect 36138 309978 36758 310046
rect 36138 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 36758 309978
rect 36138 292350 36758 309922
rect 36138 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 36758 292350
rect 36138 292226 36758 292294
rect 36138 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 36758 292226
rect 36138 292102 36758 292170
rect 36138 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 36758 292102
rect 36138 291978 36758 292046
rect 36138 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 36758 291978
rect 36138 274350 36758 291922
rect 36138 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 36758 274350
rect 36138 274226 36758 274294
rect 36138 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 36758 274226
rect 36138 274102 36758 274170
rect 36138 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 36758 274102
rect 36138 273978 36758 274046
rect 36138 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 36758 273978
rect 36138 256350 36758 273922
rect 36138 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 36758 256350
rect 36138 256226 36758 256294
rect 36138 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 36758 256226
rect 36138 256102 36758 256170
rect 36138 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 36758 256102
rect 36138 255978 36758 256046
rect 36138 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 36758 255978
rect 36138 238350 36758 255922
rect 36138 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 36758 238350
rect 36138 238226 36758 238294
rect 36138 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 36758 238226
rect 36138 238102 36758 238170
rect 36138 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 36758 238102
rect 36138 237978 36758 238046
rect 36138 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 36758 237978
rect 33516 236068 33572 236078
rect 31052 107314 31108 107324
rect 33404 224218 33460 224228
rect 29372 64978 29428 64988
rect 26796 4162 26852 4172
rect 33404 4228 33460 224162
rect 33516 4978 33572 236012
rect 36138 220350 36758 237922
rect 39676 373798 39732 373808
rect 39676 237972 39732 373742
rect 39676 237906 39732 237916
rect 39858 370350 40478 387922
rect 39858 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 40478 370350
rect 39858 370226 40478 370294
rect 39858 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 40478 370226
rect 39858 370102 40478 370170
rect 39858 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 40478 370102
rect 39858 369978 40478 370046
rect 39858 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 40478 369978
rect 39858 352350 40478 369922
rect 66858 382350 67478 390964
rect 66858 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 67478 382350
rect 66858 382226 67478 382294
rect 66858 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 67478 382226
rect 66858 382102 67478 382170
rect 66858 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 67478 382102
rect 66858 381978 67478 382046
rect 66858 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 67478 381978
rect 66858 364350 67478 381922
rect 66858 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 67478 364350
rect 66858 364226 67478 364294
rect 66858 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 67478 364226
rect 66858 364102 67478 364170
rect 66858 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 67478 364102
rect 66858 363978 67478 364046
rect 66858 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 67478 363978
rect 66858 355174 67478 363922
rect 70578 388350 71198 399778
rect 70578 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 71198 388350
rect 70578 388226 71198 388294
rect 70578 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 71198 388226
rect 70578 388102 71198 388170
rect 70578 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 71198 388102
rect 70578 387978 71198 388046
rect 70578 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 71198 387978
rect 70578 370350 71198 387922
rect 70578 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 71198 370350
rect 70578 370226 71198 370294
rect 70578 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 71198 370226
rect 70578 370102 71198 370170
rect 70578 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 71198 370102
rect 70578 369978 71198 370046
rect 70578 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 71198 369978
rect 70578 355174 71198 369922
rect 86492 397460 86548 397470
rect 86492 356158 86548 397404
rect 86492 356092 86548 356102
rect 89852 354358 89908 400316
rect 89964 358708 90020 403228
rect 89964 358642 90020 358652
rect 91532 361284 91588 361294
rect 89852 354292 89908 354302
rect 39858 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 40478 352350
rect 39858 352226 40478 352294
rect 39858 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 40478 352226
rect 39858 352102 40478 352170
rect 39858 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 40478 352102
rect 39858 351978 40478 352046
rect 39858 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 40478 351978
rect 39858 334350 40478 351922
rect 69808 352350 70128 352384
rect 69808 352294 69878 352350
rect 69934 352294 70002 352350
rect 70058 352294 70128 352350
rect 69808 352226 70128 352294
rect 69808 352170 69878 352226
rect 69934 352170 70002 352226
rect 70058 352170 70128 352226
rect 69808 352102 70128 352170
rect 69808 352046 69878 352102
rect 69934 352046 70002 352102
rect 70058 352046 70128 352102
rect 69808 351978 70128 352046
rect 69808 351922 69878 351978
rect 69934 351922 70002 351978
rect 70058 351922 70128 351978
rect 69808 351888 70128 351922
rect 54448 346350 54768 346384
rect 54448 346294 54518 346350
rect 54574 346294 54642 346350
rect 54698 346294 54768 346350
rect 54448 346226 54768 346294
rect 54448 346170 54518 346226
rect 54574 346170 54642 346226
rect 54698 346170 54768 346226
rect 54448 346102 54768 346170
rect 54448 346046 54518 346102
rect 54574 346046 54642 346102
rect 54698 346046 54768 346102
rect 54448 345978 54768 346046
rect 54448 345922 54518 345978
rect 54574 345922 54642 345978
rect 54698 345922 54768 345978
rect 54448 345888 54768 345922
rect 85168 346350 85488 346384
rect 85168 346294 85238 346350
rect 85294 346294 85362 346350
rect 85418 346294 85488 346350
rect 85168 346226 85488 346294
rect 85168 346170 85238 346226
rect 85294 346170 85362 346226
rect 85418 346170 85488 346226
rect 85168 346102 85488 346170
rect 85168 346046 85238 346102
rect 85294 346046 85362 346102
rect 85418 346046 85488 346102
rect 85168 345978 85488 346046
rect 85168 345922 85238 345978
rect 85294 345922 85362 345978
rect 85418 345922 85488 345978
rect 85168 345888 85488 345922
rect 39858 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 40478 334350
rect 39858 334226 40478 334294
rect 39858 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 40478 334226
rect 39858 334102 40478 334170
rect 39858 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 40478 334102
rect 39858 333978 40478 334046
rect 39858 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 40478 333978
rect 39858 316350 40478 333922
rect 54448 328350 54768 328384
rect 54448 328294 54518 328350
rect 54574 328294 54642 328350
rect 54698 328294 54768 328350
rect 54448 328226 54768 328294
rect 54448 328170 54518 328226
rect 54574 328170 54642 328226
rect 54698 328170 54768 328226
rect 54448 328102 54768 328170
rect 54448 328046 54518 328102
rect 54574 328046 54642 328102
rect 54698 328046 54768 328102
rect 54448 327978 54768 328046
rect 54448 327922 54518 327978
rect 54574 327922 54642 327978
rect 54698 327922 54768 327978
rect 54448 327888 54768 327922
rect 66858 328350 67478 337658
rect 69808 334350 70128 334384
rect 69808 334294 69878 334350
rect 69934 334294 70002 334350
rect 70058 334294 70128 334350
rect 69808 334226 70128 334294
rect 69808 334170 69878 334226
rect 69934 334170 70002 334226
rect 70058 334170 70128 334226
rect 69808 334102 70128 334170
rect 69808 334046 69878 334102
rect 69934 334046 70002 334102
rect 70058 334046 70128 334102
rect 69808 333978 70128 334046
rect 69808 333922 69878 333978
rect 69934 333922 70002 333978
rect 70058 333922 70128 333978
rect 69808 333888 70128 333922
rect 70578 334350 71198 337658
rect 70578 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 71198 334350
rect 70578 334226 71198 334294
rect 70578 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 71198 334226
rect 70578 334102 71198 334170
rect 70578 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 71198 334102
rect 70578 333978 71198 334046
rect 70578 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 71198 333978
rect 66858 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 67478 328350
rect 66858 328226 67478 328294
rect 66858 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 67478 328226
rect 66858 328102 67478 328170
rect 66858 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 67478 328102
rect 66858 327978 67478 328046
rect 66858 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 67478 327978
rect 39858 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 40478 316350
rect 39858 316226 40478 316294
rect 39858 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 40478 316226
rect 39858 316102 40478 316170
rect 39858 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 40478 316102
rect 39858 315978 40478 316046
rect 39858 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 40478 315978
rect 39858 298350 40478 315922
rect 39858 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 40478 298350
rect 39858 298226 40478 298294
rect 39858 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 40478 298226
rect 39858 298102 40478 298170
rect 39858 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 40478 298102
rect 39858 297978 40478 298046
rect 39858 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 40478 297978
rect 39858 280350 40478 297922
rect 60396 311698 60452 311708
rect 60396 293972 60452 311642
rect 60396 293906 60452 293916
rect 66858 310350 67478 327922
rect 66858 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 67478 310350
rect 66858 310226 67478 310294
rect 66858 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 67478 310226
rect 66858 310102 67478 310170
rect 66858 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 67478 310102
rect 66858 309978 67478 310046
rect 66858 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 67478 309978
rect 66858 292350 67478 309922
rect 66858 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 67478 292350
rect 66858 292226 67478 292294
rect 66858 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 67478 292226
rect 66858 292102 67478 292170
rect 66858 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 67478 292102
rect 66858 291978 67478 292046
rect 66858 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 67478 291978
rect 66858 289134 67478 291922
rect 70578 316350 71198 333922
rect 91532 330958 91588 361228
rect 91644 356158 91700 356168
rect 91644 332758 91700 356102
rect 91644 332692 91700 332702
rect 91532 330892 91588 330902
rect 85168 328350 85488 328384
rect 85168 328294 85238 328350
rect 85294 328294 85362 328350
rect 85418 328294 85488 328350
rect 85168 328226 85488 328294
rect 85168 328170 85238 328226
rect 85294 328170 85362 328226
rect 85418 328170 85488 328226
rect 85168 328102 85488 328170
rect 85168 328046 85238 328102
rect 85294 328046 85362 328102
rect 85418 328046 85488 328102
rect 85168 327978 85488 328046
rect 85168 327922 85238 327978
rect 85294 327922 85362 327978
rect 85418 327922 85488 327978
rect 85168 327888 85488 327922
rect 70578 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 71198 316350
rect 70578 316226 71198 316294
rect 70578 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 71198 316226
rect 70578 316102 71198 316170
rect 70578 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 71198 316102
rect 70578 315978 71198 316046
rect 70578 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 71198 315978
rect 70578 298350 71198 315922
rect 70578 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 71198 298350
rect 70578 298226 71198 298294
rect 70578 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 71198 298226
rect 70578 298102 71198 298170
rect 70578 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 71198 298102
rect 70578 297978 71198 298046
rect 70578 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 71198 297978
rect 70578 289134 71198 297922
rect 71820 294058 71876 294068
rect 71820 292404 71876 294002
rect 71820 292338 71876 292348
rect 84588 293878 84644 293888
rect 84588 292404 84644 293822
rect 84588 292338 84644 292348
rect 92316 290500 92372 290510
rect 92316 285796 92372 290444
rect 92316 285730 92372 285740
rect 39858 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 40478 280350
rect 39858 280226 40478 280294
rect 39858 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 40478 280226
rect 39858 280102 40478 280170
rect 39858 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 40478 280102
rect 39858 279978 40478 280046
rect 39858 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 40478 279978
rect 39858 262350 40478 279922
rect 59808 280350 60128 280384
rect 59808 280294 59878 280350
rect 59934 280294 60002 280350
rect 60058 280294 60128 280350
rect 59808 280226 60128 280294
rect 59808 280170 59878 280226
rect 59934 280170 60002 280226
rect 60058 280170 60128 280226
rect 59808 280102 60128 280170
rect 59808 280046 59878 280102
rect 59934 280046 60002 280102
rect 60058 280046 60128 280102
rect 59808 279978 60128 280046
rect 59808 279922 59878 279978
rect 59934 279922 60002 279978
rect 60058 279922 60128 279978
rect 59808 279888 60128 279922
rect 44448 274350 44768 274384
rect 44448 274294 44518 274350
rect 44574 274294 44642 274350
rect 44698 274294 44768 274350
rect 44448 274226 44768 274294
rect 44448 274170 44518 274226
rect 44574 274170 44642 274226
rect 44698 274170 44768 274226
rect 44448 274102 44768 274170
rect 44448 274046 44518 274102
rect 44574 274046 44642 274102
rect 44698 274046 44768 274102
rect 44448 273978 44768 274046
rect 44448 273922 44518 273978
rect 44574 273922 44642 273978
rect 44698 273922 44768 273978
rect 44448 273888 44768 273922
rect 75168 274350 75488 274384
rect 75168 274294 75238 274350
rect 75294 274294 75362 274350
rect 75418 274294 75488 274350
rect 75168 274226 75488 274294
rect 75168 274170 75238 274226
rect 75294 274170 75362 274226
rect 75418 274170 75488 274226
rect 75168 274102 75488 274170
rect 75168 274046 75238 274102
rect 75294 274046 75362 274102
rect 75418 274046 75488 274102
rect 75168 273978 75488 274046
rect 75168 273922 75238 273978
rect 75294 273922 75362 273978
rect 75418 273922 75488 273978
rect 75168 273888 75488 273922
rect 39858 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 40478 262350
rect 39858 262226 40478 262294
rect 39858 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 40478 262226
rect 39858 262102 40478 262170
rect 39858 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 40478 262102
rect 39858 261978 40478 262046
rect 39858 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 40478 261978
rect 39858 244350 40478 261922
rect 59808 262350 60128 262384
rect 59808 262294 59878 262350
rect 59934 262294 60002 262350
rect 60058 262294 60128 262350
rect 59808 262226 60128 262294
rect 59808 262170 59878 262226
rect 59934 262170 60002 262226
rect 60058 262170 60128 262226
rect 59808 262102 60128 262170
rect 59808 262046 59878 262102
rect 59934 262046 60002 262102
rect 60058 262046 60128 262102
rect 59808 261978 60128 262046
rect 59808 261922 59878 261978
rect 59934 261922 60002 261978
rect 60058 261922 60128 261978
rect 59808 261888 60128 261922
rect 92428 259140 92484 404908
rect 97578 400350 98198 417922
rect 97578 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 98198 400350
rect 97578 400226 98198 400294
rect 97578 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 98198 400226
rect 97578 400102 98198 400170
rect 97578 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 98198 400102
rect 97578 399978 98198 400046
rect 97578 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 98198 399978
rect 97578 382350 98198 399922
rect 101298 460350 101918 473068
rect 101298 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 101918 460350
rect 101298 460226 101918 460294
rect 101298 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 101918 460226
rect 101298 460102 101918 460170
rect 101298 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 101918 460102
rect 101298 459978 101918 460046
rect 101298 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 101918 459978
rect 101298 442350 101918 459922
rect 101298 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 101918 442350
rect 101298 442226 101918 442294
rect 101298 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 101918 442226
rect 101298 442102 101918 442170
rect 101298 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 101918 442102
rect 101298 441978 101918 442046
rect 101298 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 101918 441978
rect 101298 424350 101918 441922
rect 101298 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 101918 424350
rect 101298 424226 101918 424294
rect 101298 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 101918 424226
rect 101298 424102 101918 424170
rect 101298 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 101918 424102
rect 101298 423978 101918 424046
rect 101298 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 101918 423978
rect 101298 406350 101918 423922
rect 101298 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 101918 406350
rect 101298 406226 101918 406294
rect 101298 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 101918 406226
rect 101298 406102 101918 406170
rect 101298 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 101918 406102
rect 101298 405978 101918 406046
rect 101298 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 101918 405978
rect 101298 388350 101918 405922
rect 101298 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 101918 388350
rect 101298 388226 101918 388294
rect 101298 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 101918 388226
rect 101298 388102 101918 388170
rect 101298 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 101918 388102
rect 101298 387978 101918 388046
rect 101298 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 101918 387978
rect 97578 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 98198 382350
rect 97578 382226 98198 382294
rect 97578 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 98198 382226
rect 97578 382102 98198 382170
rect 97578 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 98198 382102
rect 97578 381978 98198 382046
rect 97578 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 98198 381978
rect 97578 364350 98198 381922
rect 97578 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 98198 364350
rect 97578 364226 98198 364294
rect 97578 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 98198 364226
rect 97578 364102 98198 364170
rect 97578 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 98198 364102
rect 97578 363978 98198 364046
rect 97578 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 98198 363978
rect 93324 358708 93380 358718
rect 92428 259074 92484 259084
rect 93212 330958 93268 330968
rect 93212 320878 93268 330902
rect 44448 256350 44768 256384
rect 44448 256294 44518 256350
rect 44574 256294 44642 256350
rect 44698 256294 44768 256350
rect 44448 256226 44768 256294
rect 44448 256170 44518 256226
rect 44574 256170 44642 256226
rect 44698 256170 44768 256226
rect 44448 256102 44768 256170
rect 44448 256046 44518 256102
rect 44574 256046 44642 256102
rect 44698 256046 44768 256102
rect 44448 255978 44768 256046
rect 44448 255922 44518 255978
rect 44574 255922 44642 255978
rect 44698 255922 44768 255978
rect 44448 255888 44768 255922
rect 75168 256350 75488 256384
rect 75168 256294 75238 256350
rect 75294 256294 75362 256350
rect 75418 256294 75488 256350
rect 75168 256226 75488 256294
rect 75168 256170 75238 256226
rect 75294 256170 75362 256226
rect 75418 256170 75488 256226
rect 75168 256102 75488 256170
rect 75168 256046 75238 256102
rect 75294 256046 75362 256102
rect 75418 256046 75488 256102
rect 75168 255978 75488 256046
rect 75168 255922 75238 255978
rect 75294 255922 75362 255978
rect 75418 255922 75488 255978
rect 75168 255888 75488 255922
rect 39858 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 40478 244350
rect 39858 244226 40478 244294
rect 39858 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 40478 244226
rect 39858 244102 40478 244170
rect 39858 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 40478 244102
rect 39858 243978 40478 244046
rect 39858 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 40478 243978
rect 36138 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 36758 220350
rect 36138 220226 36758 220294
rect 36138 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 36758 220226
rect 36138 220102 36758 220170
rect 36138 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 36758 220102
rect 36138 219978 36758 220046
rect 36138 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 36758 219978
rect 33516 4912 33572 4922
rect 35196 215908 35252 215918
rect 35196 4798 35252 215852
rect 35196 4732 35252 4742
rect 36138 202350 36758 219922
rect 36138 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 36758 202350
rect 36138 202226 36758 202294
rect 36138 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 36758 202226
rect 36138 202102 36758 202170
rect 36138 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 36758 202102
rect 36138 201978 36758 202046
rect 36138 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 36758 201978
rect 36138 184350 36758 201922
rect 36138 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 36758 184350
rect 36138 184226 36758 184294
rect 36138 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 36758 184226
rect 36138 184102 36758 184170
rect 36138 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 36758 184102
rect 36138 183978 36758 184046
rect 36138 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 36758 183978
rect 36138 166350 36758 183922
rect 36138 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 36758 166350
rect 36138 166226 36758 166294
rect 36138 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 36758 166226
rect 36138 166102 36758 166170
rect 36138 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 36758 166102
rect 36138 165978 36758 166046
rect 36138 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 36758 165978
rect 36138 148350 36758 165922
rect 36138 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 36758 148350
rect 36138 148226 36758 148294
rect 36138 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 36758 148226
rect 36138 148102 36758 148170
rect 36138 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 36758 148102
rect 36138 147978 36758 148046
rect 36138 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 36758 147978
rect 36138 130350 36758 147922
rect 36138 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 36758 130350
rect 36138 130226 36758 130294
rect 36138 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 36758 130226
rect 36138 130102 36758 130170
rect 36138 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 36758 130102
rect 36138 129978 36758 130046
rect 36138 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 36758 129978
rect 36138 112350 36758 129922
rect 36138 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 36758 112350
rect 36138 112226 36758 112294
rect 36138 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 36758 112226
rect 36138 112102 36758 112170
rect 36138 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 36758 112102
rect 36138 111978 36758 112046
rect 36138 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 36758 111978
rect 36138 94350 36758 111922
rect 36138 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 36758 94350
rect 36138 94226 36758 94294
rect 36138 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 36758 94226
rect 36138 94102 36758 94170
rect 36138 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 36758 94102
rect 36138 93978 36758 94046
rect 36138 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 36758 93978
rect 36138 76350 36758 93922
rect 36138 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 36758 76350
rect 36138 76226 36758 76294
rect 36138 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 36758 76226
rect 36138 76102 36758 76170
rect 36138 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 36758 76102
rect 36138 75978 36758 76046
rect 36138 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 36758 75978
rect 36138 58350 36758 75922
rect 36138 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 36758 58350
rect 36138 58226 36758 58294
rect 36138 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 36758 58226
rect 36138 58102 36758 58170
rect 36138 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 36758 58102
rect 36138 57978 36758 58046
rect 36138 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 36758 57978
rect 36138 40350 36758 57922
rect 36138 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 36758 40350
rect 36138 40226 36758 40294
rect 36138 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 36758 40226
rect 36138 40102 36758 40170
rect 36138 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 36758 40102
rect 36138 39978 36758 40046
rect 36138 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 36758 39978
rect 36138 22350 36758 39922
rect 36138 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 36758 22350
rect 36138 22226 36758 22294
rect 36138 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 36758 22226
rect 36138 22102 36758 22170
rect 36138 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 36758 22102
rect 36138 21978 36758 22046
rect 36138 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 36758 21978
rect 33404 4162 33460 4172
rect 36138 4350 36758 21922
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 226350 40478 243922
rect 59808 244350 60128 244384
rect 59808 244294 59878 244350
rect 59934 244294 60002 244350
rect 60058 244294 60128 244350
rect 59808 244226 60128 244294
rect 59808 244170 59878 244226
rect 59934 244170 60002 244226
rect 60058 244170 60128 244226
rect 59808 244102 60128 244170
rect 59808 244046 59878 244102
rect 59934 244046 60002 244102
rect 60058 244046 60128 244102
rect 59808 243978 60128 244046
rect 59808 243922 59878 243978
rect 59934 243922 60002 243978
rect 60058 243922 60128 243978
rect 59808 243888 60128 243922
rect 93212 243628 93268 320822
rect 93324 322498 93380 358652
rect 93660 354358 93716 354368
rect 93324 254884 93380 322442
rect 93324 254818 93380 254828
rect 93436 332758 93492 332768
rect 93436 320698 93492 332702
rect 93436 246372 93492 320642
rect 93660 320518 93716 354302
rect 93660 250628 93716 320462
rect 97578 346350 98198 363922
rect 97578 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 98198 346350
rect 97578 346226 98198 346294
rect 97578 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 98198 346226
rect 97578 346102 98198 346170
rect 97578 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 98198 346102
rect 97578 345978 98198 346046
rect 97578 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 98198 345978
rect 97578 328350 98198 345922
rect 97578 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 98198 328350
rect 97578 328226 98198 328294
rect 97578 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 98198 328226
rect 97578 328102 98198 328170
rect 97578 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 98198 328102
rect 97578 327978 98198 328046
rect 97578 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 98198 327978
rect 97578 310350 98198 327922
rect 97578 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 98198 310350
rect 97578 310226 98198 310294
rect 97578 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 98198 310226
rect 97578 310102 98198 310170
rect 97578 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 98198 310102
rect 97578 309978 98198 310046
rect 97578 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 98198 309978
rect 97578 292350 98198 309922
rect 97578 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 98198 292350
rect 97578 292226 98198 292294
rect 97578 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 98198 292226
rect 97578 292102 98198 292170
rect 97578 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 98198 292102
rect 97578 291978 98198 292046
rect 97578 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 98198 291978
rect 93996 288932 94052 288942
rect 93996 286468 94052 288876
rect 93996 286402 94052 286412
rect 93996 285460 94052 285470
rect 93996 280420 94052 285404
rect 93996 280354 94052 280364
rect 93996 276164 94052 276174
rect 93996 275698 94052 276108
rect 93996 275632 94052 275642
rect 97578 274350 98198 291922
rect 97578 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 98198 274350
rect 97578 274226 98198 274294
rect 97578 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 98198 274226
rect 97578 274102 98198 274170
rect 97578 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 98198 274102
rect 97578 273978 98198 274046
rect 97578 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 98198 273978
rect 93996 271908 94052 271918
rect 93996 270658 94052 271852
rect 93996 270592 94052 270602
rect 93660 250562 93716 250572
rect 97578 256350 98198 273922
rect 97578 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 98198 256350
rect 97578 256226 98198 256294
rect 97578 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 98198 256226
rect 97578 256102 98198 256170
rect 97578 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 98198 256102
rect 97578 255978 98198 256046
rect 97578 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 98198 255978
rect 93436 246306 93492 246316
rect 93212 243572 93492 243628
rect 93436 242004 93492 243572
rect 93436 241938 93492 241948
rect 62636 238532 62692 238542
rect 62636 237718 62692 238476
rect 62636 237652 62692 237662
rect 64428 238532 64484 238542
rect 64428 237538 64484 238476
rect 64428 237472 64484 237482
rect 66858 238350 67478 241266
rect 80444 240996 80500 241006
rect 80444 240772 80500 240940
rect 80444 240706 80500 240716
rect 66858 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 67478 238350
rect 66858 238226 67478 238294
rect 66858 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 67478 238226
rect 66858 238102 67478 238170
rect 66858 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 67478 238102
rect 66858 237978 67478 238046
rect 66858 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 67478 237978
rect 39858 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 40478 226350
rect 39858 226226 40478 226294
rect 39858 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 40478 226226
rect 39858 226102 40478 226170
rect 39858 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 40478 226102
rect 39858 225978 40478 226046
rect 43484 234612 43540 234622
rect 39858 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 40478 225978
rect 39858 208350 40478 225922
rect 43372 225988 43428 225998
rect 41020 220948 41076 220958
rect 39858 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 40478 208350
rect 39858 208226 40478 208294
rect 39858 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 40478 208226
rect 39858 208102 40478 208170
rect 39858 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 40478 208102
rect 39858 207978 40478 208046
rect 39858 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 40478 207978
rect 39858 190350 40478 207922
rect 39858 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 40478 190350
rect 39858 190226 40478 190294
rect 39858 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 40478 190226
rect 39858 190102 40478 190170
rect 39858 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 40478 190102
rect 39858 189978 40478 190046
rect 39858 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 40478 189978
rect 39858 172350 40478 189922
rect 39858 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 40478 172350
rect 39858 172226 40478 172294
rect 39858 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 40478 172226
rect 39858 172102 40478 172170
rect 39858 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 40478 172102
rect 39858 171978 40478 172046
rect 39858 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 40478 171978
rect 39858 154350 40478 171922
rect 39858 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 40478 154350
rect 39858 154226 40478 154294
rect 39858 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 40478 154226
rect 39858 154102 40478 154170
rect 39858 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 40478 154102
rect 39858 153978 40478 154046
rect 39858 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 40478 153978
rect 39858 136350 40478 153922
rect 39858 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 40478 136350
rect 39858 136226 40478 136294
rect 39858 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 40478 136226
rect 39858 136102 40478 136170
rect 39858 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 40478 136102
rect 39858 135978 40478 136046
rect 39858 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 40478 135978
rect 39858 118350 40478 135922
rect 39858 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 40478 118350
rect 39858 118226 40478 118294
rect 39858 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 40478 118226
rect 39858 118102 40478 118170
rect 39858 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 40478 118102
rect 39858 117978 40478 118046
rect 39858 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 40478 117978
rect 39858 100350 40478 117922
rect 39858 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 40478 100350
rect 39858 100226 40478 100294
rect 39858 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 40478 100226
rect 39858 100102 40478 100170
rect 39858 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 40478 100102
rect 39858 99978 40478 100046
rect 39858 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 40478 99978
rect 39858 82350 40478 99922
rect 39858 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 40478 82350
rect 39858 82226 40478 82294
rect 39858 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 40478 82226
rect 39858 82102 40478 82170
rect 39858 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 40478 82102
rect 39858 81978 40478 82046
rect 39858 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 40478 81978
rect 39858 64350 40478 81922
rect 39858 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 40478 64350
rect 39858 64226 40478 64294
rect 39858 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 40478 64226
rect 39858 64102 40478 64170
rect 39858 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 40478 64102
rect 39858 63978 40478 64046
rect 39858 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 40478 63978
rect 39858 46350 40478 63922
rect 39858 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 40478 46350
rect 39858 46226 40478 46294
rect 39858 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 40478 46226
rect 39858 46102 40478 46170
rect 39858 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 40478 46102
rect 39858 45978 40478 46046
rect 39858 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 40478 45978
rect 39858 28350 40478 45922
rect 39858 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 40478 28350
rect 39858 28226 40478 28294
rect 39858 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 40478 28226
rect 39858 28102 40478 28170
rect 39858 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 40478 28102
rect 39858 27978 40478 28046
rect 39858 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 40478 27978
rect 39858 10350 40478 27922
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 39858 -1120 40478 9922
rect 40908 214452 40964 214462
rect 40908 4788 40964 214396
rect 40908 4722 40964 4732
rect 41020 4228 41076 220892
rect 41132 210178 41188 210188
rect 41132 206164 41188 210122
rect 41132 206098 41188 206108
rect 41468 208738 41524 208748
rect 41468 196588 41524 208682
rect 41132 196532 41524 196588
rect 41132 163828 41188 196532
rect 41132 163762 41188 163772
rect 43372 48132 43428 225932
rect 43484 49812 43540 234556
rect 43484 49746 43540 49756
rect 43596 229572 43652 229582
rect 43372 48066 43428 48076
rect 43596 4676 43652 229516
rect 66858 220350 67478 237922
rect 66858 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 67478 220350
rect 66858 220226 67478 220294
rect 66858 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 67478 220226
rect 66858 220102 67478 220170
rect 66858 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 67478 220102
rect 66858 219978 67478 220046
rect 66858 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 67478 219978
rect 66858 210574 67478 219922
rect 97578 238350 98198 255922
rect 97578 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 98198 238350
rect 97578 238226 98198 238294
rect 97578 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 98198 238226
rect 97578 238102 98198 238170
rect 97578 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 98198 238102
rect 97578 237978 98198 238046
rect 97578 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 98198 237978
rect 97578 220350 98198 237922
rect 100156 385252 100212 385262
rect 100156 237538 100212 385196
rect 100156 237472 100212 237482
rect 101298 370350 101918 387922
rect 101298 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 101918 370350
rect 101298 370226 101918 370294
rect 101298 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 101918 370226
rect 101298 370102 101918 370170
rect 101298 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 101918 370102
rect 101298 369978 101918 370046
rect 101298 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 101918 369978
rect 101298 352350 101918 369922
rect 101298 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 101918 352350
rect 101298 352226 101918 352294
rect 101298 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 101918 352226
rect 101298 352102 101918 352170
rect 101298 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 101918 352102
rect 101298 351978 101918 352046
rect 101298 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 101918 351978
rect 101298 334350 101918 351922
rect 128298 472350 128918 488368
rect 128298 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 128918 472350
rect 128298 472226 128918 472294
rect 128298 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 128918 472226
rect 128298 472102 128918 472170
rect 128298 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 128918 472102
rect 128298 471978 128918 472046
rect 128298 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 128918 471978
rect 128298 454350 128918 471922
rect 128298 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 128918 454350
rect 128298 454226 128918 454294
rect 128298 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 128918 454226
rect 128298 454102 128918 454170
rect 128298 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 128918 454102
rect 128298 453978 128918 454046
rect 128298 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 128918 453978
rect 128298 436350 128918 453922
rect 128298 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 128918 436350
rect 128298 436226 128918 436294
rect 128298 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 128918 436226
rect 128298 436102 128918 436170
rect 128298 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 128918 436102
rect 128298 435978 128918 436046
rect 128298 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 128918 435978
rect 128298 418350 128918 435922
rect 128298 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 128918 418350
rect 128298 418226 128918 418294
rect 128298 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 128918 418226
rect 128298 418102 128918 418170
rect 128298 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 128918 418102
rect 128298 417978 128918 418046
rect 128298 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 128918 417978
rect 128298 400350 128918 417922
rect 128298 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 128918 400350
rect 128298 400226 128918 400294
rect 128298 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 128918 400226
rect 128298 400102 128918 400170
rect 128298 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 128918 400102
rect 128298 399978 128918 400046
rect 128298 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 128918 399978
rect 128298 382350 128918 399922
rect 128298 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 128918 382350
rect 128298 382226 128918 382294
rect 128298 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 128918 382226
rect 128298 382102 128918 382170
rect 128298 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 128918 382102
rect 128298 381978 128918 382046
rect 128298 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 128918 381978
rect 128298 364350 128918 381922
rect 128298 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 128918 364350
rect 128298 364226 128918 364294
rect 128298 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 128918 364226
rect 128298 364102 128918 364170
rect 128298 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 128918 364102
rect 128298 363978 128918 364046
rect 128298 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 128918 363978
rect 124448 346350 124768 346384
rect 124448 346294 124518 346350
rect 124574 346294 124642 346350
rect 124698 346294 124768 346350
rect 124448 346226 124768 346294
rect 124448 346170 124518 346226
rect 124574 346170 124642 346226
rect 124698 346170 124768 346226
rect 124448 346102 124768 346170
rect 124448 346046 124518 346102
rect 124574 346046 124642 346102
rect 124698 346046 124768 346102
rect 124448 345978 124768 346046
rect 124448 345922 124518 345978
rect 124574 345922 124642 345978
rect 124698 345922 124768 345978
rect 124448 345888 124768 345922
rect 128298 346350 128918 363922
rect 128298 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 128918 346350
rect 128298 346226 128918 346294
rect 128298 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 128918 346226
rect 128298 346102 128918 346170
rect 128298 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 128918 346102
rect 128298 345978 128918 346046
rect 128298 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 128918 345978
rect 101298 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 101918 334350
rect 101298 334226 101918 334294
rect 101298 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 101918 334226
rect 101298 334102 101918 334170
rect 101298 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 101918 334102
rect 101298 333978 101918 334046
rect 101298 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 101918 333978
rect 101298 316350 101918 333922
rect 124448 328350 124768 328384
rect 124448 328294 124518 328350
rect 124574 328294 124642 328350
rect 124698 328294 124768 328350
rect 124448 328226 124768 328294
rect 124448 328170 124518 328226
rect 124574 328170 124642 328226
rect 124698 328170 124768 328226
rect 124448 328102 124768 328170
rect 124448 328046 124518 328102
rect 124574 328046 124642 328102
rect 124698 328046 124768 328102
rect 124448 327978 124768 328046
rect 124448 327922 124518 327978
rect 124574 327922 124642 327978
rect 124698 327922 124768 327978
rect 124448 327888 124768 327922
rect 128298 328350 128918 345922
rect 128298 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 128918 328350
rect 128298 328226 128918 328294
rect 128298 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 128918 328226
rect 128298 328102 128918 328170
rect 128298 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 128918 328102
rect 128298 327978 128918 328046
rect 128298 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 128918 327978
rect 101298 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 101918 316350
rect 101298 316226 101918 316294
rect 101298 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 101918 316226
rect 101298 316102 101918 316170
rect 101298 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 101918 316102
rect 101298 315978 101918 316046
rect 101298 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 101918 315978
rect 101298 298350 101918 315922
rect 101298 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 101918 298350
rect 101298 298226 101918 298294
rect 101298 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 101918 298226
rect 101298 298102 101918 298170
rect 101298 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 101918 298102
rect 101298 297978 101918 298046
rect 101298 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 101918 297978
rect 101298 280350 101918 297922
rect 128298 310350 128918 327922
rect 128298 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 128918 310350
rect 128298 310226 128918 310294
rect 128298 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 128918 310226
rect 128298 310102 128918 310170
rect 128298 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 128918 310102
rect 128298 309978 128918 310046
rect 128298 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 128918 309978
rect 128298 292350 128918 309922
rect 128298 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 128918 292350
rect 128298 292226 128918 292294
rect 128298 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 128918 292226
rect 128298 292102 128918 292170
rect 128298 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 128918 292102
rect 128298 291978 128918 292046
rect 128298 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 128918 291978
rect 101298 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 101918 280350
rect 101298 280226 101918 280294
rect 101298 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 101918 280226
rect 101298 280102 101918 280170
rect 101298 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 101918 280102
rect 101298 279978 101918 280046
rect 101298 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 101918 279978
rect 101298 262350 101918 279922
rect 101298 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 101918 262350
rect 101298 262226 101918 262294
rect 101298 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 101918 262226
rect 101298 262102 101918 262170
rect 101298 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 101918 262102
rect 101298 261978 101918 262046
rect 101298 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 101918 261978
rect 101298 244350 101918 261922
rect 101298 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 101918 244350
rect 101298 244226 101918 244294
rect 101298 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 101918 244226
rect 101298 244102 101918 244170
rect 101298 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 101918 244102
rect 101298 243978 101918 244046
rect 101298 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 101918 243978
rect 97578 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 98198 220350
rect 97578 220226 98198 220294
rect 97578 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 98198 220226
rect 97578 220102 98198 220170
rect 97578 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 98198 220102
rect 97578 219978 98198 220046
rect 97578 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 98198 219978
rect 97578 210574 98198 219922
rect 101298 226350 101918 243922
rect 101298 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 101918 226350
rect 101298 226226 101918 226294
rect 101298 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 101918 226226
rect 101298 226102 101918 226170
rect 101298 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 101918 226102
rect 101298 225978 101918 226046
rect 101298 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 101918 225978
rect 101298 210574 101918 225922
rect 115052 288036 115108 288046
rect 115052 210868 115108 287980
rect 115052 210802 115108 210812
rect 128298 274350 128918 291922
rect 128298 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 128918 274350
rect 128298 274226 128918 274294
rect 128298 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 128918 274226
rect 128298 274102 128918 274170
rect 128298 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 128918 274102
rect 128298 273978 128918 274046
rect 128298 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 128918 273978
rect 128298 256350 128918 273922
rect 128298 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 128918 256350
rect 128298 256226 128918 256294
rect 128298 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 128918 256226
rect 128298 256102 128918 256170
rect 128298 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 128918 256102
rect 128298 255978 128918 256046
rect 128298 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 128918 255978
rect 128298 238350 128918 255922
rect 128298 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 128918 238350
rect 128298 238226 128918 238294
rect 128298 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 128918 238226
rect 128298 238102 128918 238170
rect 128298 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 128918 238102
rect 128298 237978 128918 238046
rect 128298 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 128918 237978
rect 128298 220350 128918 237922
rect 128298 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 128918 220350
rect 128298 220226 128918 220294
rect 128298 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 128918 220226
rect 128298 220102 128918 220170
rect 128298 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 128918 220102
rect 128298 219978 128918 220046
rect 128298 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 128918 219978
rect 128298 210574 128918 219922
rect 132018 478350 132638 490708
rect 132018 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 132638 478350
rect 132018 478226 132638 478294
rect 132018 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 132638 478226
rect 132018 478102 132638 478170
rect 132018 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 132638 478102
rect 132018 477978 132638 478046
rect 132018 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 132638 477978
rect 132018 460350 132638 477922
rect 132018 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 132638 460350
rect 132018 460226 132638 460294
rect 132018 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 132638 460226
rect 132018 460102 132638 460170
rect 132018 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 132638 460102
rect 132018 459978 132638 460046
rect 132018 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 132638 459978
rect 132018 442350 132638 459922
rect 132018 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 132638 442350
rect 132018 442226 132638 442294
rect 132018 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 132638 442226
rect 132018 442102 132638 442170
rect 132018 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 132638 442102
rect 132018 441978 132638 442046
rect 132018 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 132638 441978
rect 132018 424350 132638 441922
rect 132018 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 132638 424350
rect 132018 424226 132638 424294
rect 132018 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 132638 424226
rect 132018 424102 132638 424170
rect 132018 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 132638 424102
rect 132018 423978 132638 424046
rect 132018 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 132638 423978
rect 132018 406350 132638 423922
rect 150332 469588 150388 469598
rect 150332 407998 150388 469532
rect 157052 409438 157108 587132
rect 157052 409372 157108 409382
rect 159018 580350 159638 596784
rect 159018 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 159638 580350
rect 159018 580226 159638 580294
rect 159018 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 159638 580226
rect 159018 580102 159638 580170
rect 159018 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 159638 580102
rect 159018 579978 159638 580046
rect 159018 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 159638 579978
rect 159018 562350 159638 579922
rect 159018 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 159638 562350
rect 159018 562226 159638 562294
rect 159018 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 159638 562226
rect 159018 562102 159638 562170
rect 159018 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 159638 562102
rect 159018 561978 159638 562046
rect 159018 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 159638 561978
rect 159018 544350 159638 561922
rect 159018 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 159638 544350
rect 159018 544226 159638 544294
rect 159018 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 159638 544226
rect 159018 544102 159638 544170
rect 159018 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 159638 544102
rect 159018 543978 159638 544046
rect 159018 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 159638 543978
rect 159018 526350 159638 543922
rect 159018 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 159638 526350
rect 159018 526226 159638 526294
rect 159018 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 159638 526226
rect 159018 526102 159638 526170
rect 159018 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 159638 526102
rect 159018 525978 159638 526046
rect 159018 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 159638 525978
rect 159018 508350 159638 525922
rect 159018 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 159638 508350
rect 159018 508226 159638 508294
rect 159018 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 159638 508226
rect 159018 508102 159638 508170
rect 159018 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 159638 508102
rect 159018 507978 159638 508046
rect 159018 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 159638 507978
rect 159018 490350 159638 507922
rect 159018 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 159638 490350
rect 159018 490226 159638 490294
rect 159018 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 159638 490226
rect 159018 490102 159638 490170
rect 159018 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 159638 490102
rect 159018 489978 159638 490046
rect 159018 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 159638 489978
rect 159018 472350 159638 489922
rect 159018 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 159638 472350
rect 159018 472226 159638 472294
rect 159018 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 159638 472226
rect 159018 472102 159638 472170
rect 159018 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 159638 472102
rect 159018 471978 159638 472046
rect 159018 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 159638 471978
rect 159018 454350 159638 471922
rect 159018 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 159638 454350
rect 159018 454226 159638 454294
rect 159018 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 159638 454226
rect 159018 454102 159638 454170
rect 159018 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 159638 454102
rect 159018 453978 159638 454046
rect 159018 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 159638 453978
rect 159018 436350 159638 453922
rect 159018 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 159638 436350
rect 159018 436226 159638 436294
rect 159018 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 159638 436226
rect 159018 436102 159638 436170
rect 159018 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 159638 436102
rect 159018 435978 159638 436046
rect 159018 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 159638 435978
rect 159018 418350 159638 435922
rect 159018 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 159638 418350
rect 159018 418226 159638 418294
rect 159018 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 159638 418226
rect 159018 418102 159638 418170
rect 159018 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 159638 418102
rect 159018 417978 159638 418046
rect 159018 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 159638 417978
rect 150332 407932 150388 407942
rect 132018 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 132638 406350
rect 132018 406226 132638 406294
rect 132018 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 132638 406226
rect 132018 406102 132638 406170
rect 132018 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 132638 406102
rect 132018 405978 132638 406046
rect 132018 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 132638 405978
rect 132018 388350 132638 405922
rect 132018 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 132638 388350
rect 132018 388226 132638 388294
rect 132018 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 132638 388226
rect 132018 388102 132638 388170
rect 132018 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 132638 388102
rect 132018 387978 132638 388046
rect 132018 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 132638 387978
rect 132018 370350 132638 387922
rect 132018 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 132638 370350
rect 132018 370226 132638 370294
rect 132018 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 132638 370226
rect 132018 370102 132638 370170
rect 132018 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 132638 370102
rect 132018 369978 132638 370046
rect 132018 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 132638 369978
rect 132018 352350 132638 369922
rect 159018 400350 159638 417922
rect 159018 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 159638 400350
rect 159018 400226 159638 400294
rect 159018 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 159638 400226
rect 159018 400102 159638 400170
rect 159018 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 159638 400102
rect 159018 399978 159638 400046
rect 159018 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 159638 399978
rect 159018 382350 159638 399922
rect 159018 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 159638 382350
rect 159018 382226 159638 382294
rect 159018 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 159638 382226
rect 159018 382102 159638 382170
rect 159018 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 159638 382102
rect 159018 381978 159638 382046
rect 159018 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 159638 381978
rect 159018 364350 159638 381922
rect 159018 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 159638 364350
rect 159018 364226 159638 364294
rect 159018 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 159638 364226
rect 159018 364102 159638 364170
rect 159018 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 159638 364102
rect 159018 363978 159638 364046
rect 159018 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 159638 363978
rect 132018 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 132638 352350
rect 132018 352226 132638 352294
rect 132018 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 132638 352226
rect 132018 352102 132638 352170
rect 132018 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 132638 352102
rect 132018 351978 132638 352046
rect 132018 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 132638 351978
rect 132018 334350 132638 351922
rect 139808 352350 140128 352384
rect 139808 352294 139878 352350
rect 139934 352294 140002 352350
rect 140058 352294 140128 352350
rect 139808 352226 140128 352294
rect 139808 352170 139878 352226
rect 139934 352170 140002 352226
rect 140058 352170 140128 352226
rect 139808 352102 140128 352170
rect 139808 352046 139878 352102
rect 139934 352046 140002 352102
rect 140058 352046 140128 352102
rect 139808 351978 140128 352046
rect 139808 351922 139878 351978
rect 139934 351922 140002 351978
rect 140058 351922 140128 351978
rect 139808 351888 140128 351922
rect 155168 346350 155488 346384
rect 155168 346294 155238 346350
rect 155294 346294 155362 346350
rect 155418 346294 155488 346350
rect 155168 346226 155488 346294
rect 155168 346170 155238 346226
rect 155294 346170 155362 346226
rect 155418 346170 155488 346226
rect 155168 346102 155488 346170
rect 155168 346046 155238 346102
rect 155294 346046 155362 346102
rect 155418 346046 155488 346102
rect 155168 345978 155488 346046
rect 155168 345922 155238 345978
rect 155294 345922 155362 345978
rect 155418 345922 155488 345978
rect 155168 345888 155488 345922
rect 159018 346350 159638 363922
rect 159018 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 159638 346350
rect 159018 346226 159638 346294
rect 159018 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 159638 346226
rect 159018 346102 159638 346170
rect 159018 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 159638 346102
rect 159018 345978 159638 346046
rect 159018 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 159638 345978
rect 132018 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 132638 334350
rect 132018 334226 132638 334294
rect 132018 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 132638 334226
rect 132018 334102 132638 334170
rect 132018 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 132638 334102
rect 132018 333978 132638 334046
rect 132018 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 132638 333978
rect 132018 316350 132638 333922
rect 139808 334350 140128 334384
rect 139808 334294 139878 334350
rect 139934 334294 140002 334350
rect 140058 334294 140128 334350
rect 139808 334226 140128 334294
rect 139808 334170 139878 334226
rect 139934 334170 140002 334226
rect 140058 334170 140128 334226
rect 139808 334102 140128 334170
rect 139808 334046 139878 334102
rect 139934 334046 140002 334102
rect 140058 334046 140128 334102
rect 139808 333978 140128 334046
rect 139808 333922 139878 333978
rect 139934 333922 140002 333978
rect 140058 333922 140128 333978
rect 139808 333888 140128 333922
rect 155168 328350 155488 328384
rect 155168 328294 155238 328350
rect 155294 328294 155362 328350
rect 155418 328294 155488 328350
rect 155168 328226 155488 328294
rect 155168 328170 155238 328226
rect 155294 328170 155362 328226
rect 155418 328170 155488 328226
rect 155168 328102 155488 328170
rect 155168 328046 155238 328102
rect 155294 328046 155362 328102
rect 155418 328046 155488 328102
rect 155168 327978 155488 328046
rect 155168 327922 155238 327978
rect 155294 327922 155362 327978
rect 155418 327922 155488 327978
rect 155168 327888 155488 327922
rect 159018 328350 159638 345922
rect 159018 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 159638 328350
rect 159018 328226 159638 328294
rect 159018 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 159638 328226
rect 159018 328102 159638 328170
rect 159018 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 159638 328102
rect 159018 327978 159638 328046
rect 159018 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 159638 327978
rect 132018 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 132638 316350
rect 132018 316226 132638 316294
rect 132018 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 132638 316226
rect 132018 316102 132638 316170
rect 132018 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 132638 316102
rect 132018 315978 132638 316046
rect 132018 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 132638 315978
rect 132018 298350 132638 315922
rect 132018 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 132638 298350
rect 132018 298226 132638 298294
rect 132018 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 132638 298226
rect 132018 298102 132638 298170
rect 132018 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 132638 298102
rect 132018 297978 132638 298046
rect 132018 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 132638 297978
rect 132018 280350 132638 297922
rect 159018 310350 159638 327922
rect 159018 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 159638 310350
rect 159018 310226 159638 310294
rect 159018 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 159638 310226
rect 159018 310102 159638 310170
rect 159018 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 159638 310102
rect 159018 309978 159638 310046
rect 159018 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 159638 309978
rect 159018 292350 159638 309922
rect 159018 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 159638 292350
rect 159018 292226 159638 292294
rect 159018 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 159638 292226
rect 159018 292102 159638 292170
rect 159018 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 159638 292102
rect 159018 291978 159638 292046
rect 159018 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 159638 291978
rect 159018 284908 159638 291922
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 568350 163358 585922
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 189738 580350 190358 596784
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 162738 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 163358 568350
rect 162738 568226 163358 568294
rect 162738 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 163358 568226
rect 162738 568102 163358 568170
rect 162738 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 163358 568102
rect 162738 567978 163358 568046
rect 162738 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 163358 567978
rect 162738 550350 163358 567922
rect 162738 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 163358 550350
rect 162738 550226 163358 550294
rect 162738 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 163358 550226
rect 162738 550102 163358 550170
rect 162738 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 163358 550102
rect 162738 549978 163358 550046
rect 162738 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 163358 549978
rect 162738 532350 163358 549922
rect 162738 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 163358 532350
rect 162738 532226 163358 532294
rect 162738 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 163358 532226
rect 162738 532102 163358 532170
rect 162738 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 163358 532102
rect 162738 531978 163358 532046
rect 162738 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 163358 531978
rect 162738 514350 163358 531922
rect 162738 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 163358 514350
rect 162738 514226 163358 514294
rect 162738 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 163358 514226
rect 162738 514102 163358 514170
rect 162738 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 163358 514102
rect 162738 513978 163358 514046
rect 162738 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 163358 513978
rect 162738 496350 163358 513922
rect 162738 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 163358 496350
rect 162738 496226 163358 496294
rect 162738 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 163358 496226
rect 162738 496102 163358 496170
rect 162738 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 163358 496102
rect 162738 495978 163358 496046
rect 162738 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 163358 495978
rect 162738 478350 163358 495922
rect 162738 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 163358 478350
rect 162738 478226 163358 478294
rect 162738 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 163358 478226
rect 162738 478102 163358 478170
rect 162738 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 163358 478102
rect 162738 477978 163358 478046
rect 162738 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 163358 477978
rect 162738 460350 163358 477922
rect 181356 573748 181412 573758
rect 178892 471268 178948 471278
rect 162738 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 163358 460350
rect 162738 460226 163358 460294
rect 162738 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 163358 460226
rect 162738 460102 163358 460170
rect 162738 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 163358 460102
rect 162738 459978 163358 460046
rect 162738 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 163358 459978
rect 162738 442350 163358 459922
rect 162738 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 163358 442350
rect 162738 442226 163358 442294
rect 162738 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 163358 442226
rect 162738 442102 163358 442170
rect 162738 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 163358 442102
rect 162738 441978 163358 442046
rect 162738 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 163358 441978
rect 162738 424350 163358 441922
rect 172172 467908 172228 467918
rect 162738 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 163358 424350
rect 162738 424226 163358 424294
rect 162738 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 163358 424226
rect 162738 424102 163358 424170
rect 162738 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 163358 424102
rect 162738 423978 163358 424046
rect 162738 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 163358 423978
rect 162738 406350 163358 423922
rect 162738 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 163358 406350
rect 162738 406226 163358 406294
rect 162738 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 163358 406226
rect 162738 406102 163358 406170
rect 162738 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 163358 406102
rect 162738 405978 163358 406046
rect 162738 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 163358 405978
rect 162738 388350 163358 405922
rect 162738 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 163358 388350
rect 162738 388226 163358 388294
rect 162738 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 163358 388226
rect 162738 388102 163358 388170
rect 162738 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 163358 388102
rect 162738 387978 163358 388046
rect 162738 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 163358 387978
rect 162738 370350 163358 387922
rect 162738 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 163358 370350
rect 162738 370226 163358 370294
rect 162738 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 163358 370226
rect 162738 370102 163358 370170
rect 162738 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 163358 370102
rect 162738 369978 163358 370046
rect 162738 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 163358 369978
rect 162738 352350 163358 369922
rect 162738 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 163358 352350
rect 162738 352226 163358 352294
rect 162738 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 163358 352226
rect 162738 352102 163358 352170
rect 162738 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 163358 352102
rect 162738 351978 163358 352046
rect 162738 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 163358 351978
rect 162738 334350 163358 351922
rect 162738 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 163358 334350
rect 162738 334226 163358 334294
rect 162738 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 163358 334226
rect 162738 334102 163358 334170
rect 162738 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 163358 334102
rect 162738 333978 163358 334046
rect 162738 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 163358 333978
rect 162738 316350 163358 333922
rect 167132 431956 167188 431966
rect 165900 322084 165956 322094
rect 165900 321748 165956 322028
rect 165900 321682 165956 321692
rect 162738 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 163358 316350
rect 162738 316226 163358 316294
rect 162738 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 163358 316226
rect 162738 316102 163358 316170
rect 162738 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 163358 316102
rect 162738 315978 163358 316046
rect 162738 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 163358 315978
rect 162738 298350 163358 315922
rect 162738 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 163358 298350
rect 162738 298226 163358 298294
rect 162738 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 163358 298226
rect 162738 298102 163358 298170
rect 162738 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 163358 298102
rect 162738 297978 163358 298046
rect 162738 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 163358 297978
rect 162738 282254 163358 297922
rect 165452 304948 165508 304958
rect 165452 284676 165508 304892
rect 165452 284610 165508 284620
rect 166348 286468 166404 286478
rect 132018 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 132638 280350
rect 132018 280226 132638 280294
rect 132018 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 132638 280226
rect 132018 280102 132638 280170
rect 132018 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 132638 280102
rect 132018 279978 132638 280046
rect 132018 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 132638 279978
rect 132018 262350 132638 279922
rect 147008 280350 147328 280384
rect 147008 280294 147078 280350
rect 147134 280294 147202 280350
rect 147258 280294 147328 280350
rect 147008 280226 147328 280294
rect 147008 280170 147078 280226
rect 147134 280170 147202 280226
rect 147258 280170 147328 280226
rect 147008 280102 147328 280170
rect 147008 280046 147078 280102
rect 147134 280046 147202 280102
rect 147258 280046 147328 280102
rect 147008 279978 147328 280046
rect 147008 279922 147078 279978
rect 147134 279922 147202 279978
rect 147258 279922 147328 279978
rect 147008 279888 147328 279922
rect 152832 280350 153152 280384
rect 152832 280294 152902 280350
rect 152958 280294 153026 280350
rect 153082 280294 153152 280350
rect 152832 280226 153152 280294
rect 152832 280170 152902 280226
rect 152958 280170 153026 280226
rect 153082 280170 153152 280226
rect 152832 280102 153152 280170
rect 152832 280046 152902 280102
rect 152958 280046 153026 280102
rect 153082 280046 153152 280102
rect 152832 279978 153152 280046
rect 152832 279922 152902 279978
rect 152958 279922 153026 279978
rect 153082 279922 153152 279978
rect 152832 279888 153152 279922
rect 158656 280350 158976 280384
rect 158656 280294 158726 280350
rect 158782 280294 158850 280350
rect 158906 280294 158976 280350
rect 158656 280226 158976 280294
rect 158656 280170 158726 280226
rect 158782 280170 158850 280226
rect 158906 280170 158976 280226
rect 158656 280102 158976 280170
rect 158656 280046 158726 280102
rect 158782 280046 158850 280102
rect 158906 280046 158976 280102
rect 158656 279978 158976 280046
rect 158656 279922 158726 279978
rect 158782 279922 158850 279978
rect 158906 279922 158976 279978
rect 158656 279888 158976 279922
rect 164480 280350 164800 280384
rect 164480 280294 164550 280350
rect 164606 280294 164674 280350
rect 164730 280294 164800 280350
rect 164480 280226 164800 280294
rect 164480 280170 164550 280226
rect 164606 280170 164674 280226
rect 164730 280170 164800 280226
rect 164480 280102 164800 280170
rect 164480 280046 164550 280102
rect 164606 280046 164674 280102
rect 164730 280046 164800 280102
rect 164480 279978 164800 280046
rect 164480 279922 164550 279978
rect 164606 279922 164674 279978
rect 164730 279922 164800 279978
rect 164480 279888 164800 279922
rect 153692 275698 153748 275708
rect 144096 274350 144416 274384
rect 144096 274294 144166 274350
rect 144222 274294 144290 274350
rect 144346 274294 144416 274350
rect 144096 274226 144416 274294
rect 144096 274170 144166 274226
rect 144222 274170 144290 274226
rect 144346 274170 144416 274226
rect 144096 274102 144416 274170
rect 144096 274046 144166 274102
rect 144222 274046 144290 274102
rect 144346 274046 144416 274102
rect 144096 273978 144416 274046
rect 144096 273922 144166 273978
rect 144222 273922 144290 273978
rect 144346 273922 144416 273978
rect 144096 273888 144416 273922
rect 149920 274350 150240 274384
rect 149920 274294 149990 274350
rect 150046 274294 150114 274350
rect 150170 274294 150240 274350
rect 149920 274226 150240 274294
rect 149920 274170 149990 274226
rect 150046 274170 150114 274226
rect 150170 274170 150240 274226
rect 149920 274102 150240 274170
rect 149920 274046 149990 274102
rect 150046 274046 150114 274102
rect 150170 274046 150240 274102
rect 149920 273978 150240 274046
rect 149920 273922 149990 273978
rect 150046 273922 150114 273978
rect 150170 273922 150240 273978
rect 149920 273888 150240 273922
rect 153692 267058 153748 275642
rect 155744 274350 156064 274384
rect 155744 274294 155814 274350
rect 155870 274294 155938 274350
rect 155994 274294 156064 274350
rect 155744 274226 156064 274294
rect 155744 274170 155814 274226
rect 155870 274170 155938 274226
rect 155994 274170 156064 274226
rect 155744 274102 156064 274170
rect 155744 274046 155814 274102
rect 155870 274046 155938 274102
rect 155994 274046 156064 274102
rect 155744 273978 156064 274046
rect 155744 273922 155814 273978
rect 155870 273922 155938 273978
rect 155994 273922 156064 273978
rect 155744 273888 156064 273922
rect 161568 274350 161888 274384
rect 161568 274294 161638 274350
rect 161694 274294 161762 274350
rect 161818 274294 161888 274350
rect 161568 274226 161888 274294
rect 161568 274170 161638 274226
rect 161694 274170 161762 274226
rect 161818 274170 161888 274226
rect 161568 274102 161888 274170
rect 161568 274046 161638 274102
rect 161694 274046 161762 274102
rect 161818 274046 161888 274102
rect 161568 273978 161888 274046
rect 161568 273922 161638 273978
rect 161694 273922 161762 273978
rect 161818 273922 161888 273978
rect 161568 273888 161888 273922
rect 153692 266992 153748 267002
rect 153804 270658 153860 270668
rect 153804 265438 153860 270602
rect 166348 268660 166404 286412
rect 167132 281316 167188 431900
rect 168812 428932 168868 428942
rect 168028 340138 168084 340148
rect 168028 339556 168084 340082
rect 168028 322498 168084 339500
rect 168028 322432 168084 322442
rect 168140 336868 168196 336878
rect 168140 320518 168196 336812
rect 168252 332836 168308 332846
rect 168252 320698 168308 332780
rect 168700 330932 168756 330942
rect 168364 329476 168420 329486
rect 168364 320878 168420 329420
rect 168700 329476 168756 330876
rect 168700 329410 168756 329420
rect 168364 320812 168420 320822
rect 168252 320632 168308 320642
rect 168140 320452 168196 320462
rect 168028 285460 168084 285470
rect 167132 281250 167188 281260
rect 167468 285348 167524 285358
rect 167468 280532 167524 285292
rect 167468 280466 167524 280476
rect 166348 267876 166404 268604
rect 166348 267810 166404 267820
rect 153804 265372 153860 265382
rect 132018 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 132638 262350
rect 132018 262226 132638 262294
rect 132018 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 132638 262226
rect 132018 262102 132638 262170
rect 132018 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 132638 262102
rect 132018 261978 132638 262046
rect 132018 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 132638 261978
rect 132018 244350 132638 261922
rect 162738 262350 163358 265522
rect 168028 265412 168084 285404
rect 168140 280532 168196 280542
rect 168140 278964 168196 280476
rect 168140 265860 168196 278908
rect 168140 265794 168196 265804
rect 168812 267058 168868 428876
rect 170492 380660 170548 380670
rect 168924 358596 168980 358606
rect 168924 326116 168980 358540
rect 168924 326050 168980 326060
rect 168924 313348 168980 313358
rect 168924 282436 168980 313292
rect 168924 282370 168980 282380
rect 168028 263844 168084 265356
rect 168028 263778 168084 263788
rect 162738 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 163358 262350
rect 162738 262226 163358 262294
rect 162738 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 163358 262226
rect 162738 262102 163358 262170
rect 162738 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 163358 262102
rect 162738 261978 163358 262046
rect 162738 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 163358 261978
rect 132018 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 132638 244350
rect 132018 244226 132638 244294
rect 132018 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 132638 244226
rect 132018 244102 132638 244170
rect 132018 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 132638 244102
rect 132018 243978 132638 244046
rect 132018 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 132638 243978
rect 132018 226350 132638 243922
rect 132018 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 132638 226350
rect 132018 226226 132638 226294
rect 132018 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 132638 226226
rect 132018 226102 132638 226170
rect 132018 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 132638 226102
rect 132018 225978 132638 226046
rect 132018 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 132638 225978
rect 132018 210574 132638 225922
rect 159018 256350 159638 260964
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 159018 210574 159638 219922
rect 162738 244350 163358 261922
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162738 226350 163358 243922
rect 168812 261828 168868 267002
rect 168812 236852 168868 261772
rect 170492 237718 170548 380604
rect 172172 277956 172228 467852
rect 175532 466228 175588 466238
rect 172172 277890 172228 277900
rect 173852 286916 173908 286926
rect 170492 237652 170548 237662
rect 168812 236786 168868 236796
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 162738 210574 163358 225922
rect 173852 222628 173908 286860
rect 175532 279076 175588 466172
rect 177996 313796 178052 313806
rect 177884 301476 177940 301486
rect 177212 296548 177268 296558
rect 177212 283556 177268 296492
rect 177212 283490 177268 283500
rect 175532 279010 175588 279020
rect 177884 278908 177940 301420
rect 177772 278852 177940 278908
rect 174636 272132 174692 272142
rect 174636 251218 174692 272076
rect 177772 267148 177828 278852
rect 177996 270838 178052 313740
rect 178892 280196 178948 471212
rect 179788 360836 179844 360846
rect 179788 352996 179844 360780
rect 179788 352930 179844 352940
rect 181244 316036 181300 316046
rect 179676 312676 179732 312686
rect 178892 280130 178948 280140
rect 179564 298116 179620 298126
rect 177884 270782 178052 270838
rect 177884 269758 177940 270782
rect 177996 270658 178052 270668
rect 177996 269892 178052 270602
rect 177996 269826 178052 269836
rect 177884 269702 178052 269758
rect 177772 267092 177940 267148
rect 174636 251152 174692 251162
rect 173852 222562 173908 222572
rect 177884 216132 177940 267092
rect 177884 216066 177940 216076
rect 177996 209412 178052 269702
rect 179564 239540 179620 298060
rect 179564 239474 179620 239484
rect 179676 210868 179732 312620
rect 181020 309316 181076 309326
rect 181020 214900 181076 309260
rect 181020 214834 181076 214844
rect 181132 307076 181188 307086
rect 179676 210802 179732 210812
rect 181132 209524 181188 307020
rect 181244 211092 181300 315980
rect 181356 266756 181412 573692
rect 183036 567924 183092 567934
rect 182924 402418 182980 402428
rect 182812 317156 182868 317166
rect 182700 305956 182756 305966
rect 181356 266690 181412 266700
rect 182252 285684 182308 285694
rect 182252 281988 182308 285628
rect 182252 236740 182308 281932
rect 182252 236674 182308 236684
rect 181244 211026 181300 211036
rect 182700 209636 182756 305900
rect 182812 210980 182868 317100
rect 182924 264516 182980 402362
rect 183036 265636 183092 567868
rect 187964 565124 188020 565134
rect 186396 550788 186452 550798
rect 183932 500612 183988 500622
rect 183932 285684 183988 500556
rect 184604 404038 184660 404048
rect 184492 320516 184548 320526
rect 183932 285618 183988 285628
rect 184380 311556 184436 311566
rect 183036 265570 183092 265580
rect 182924 264450 182980 264460
rect 184380 218148 184436 311500
rect 184380 218082 184436 218092
rect 182812 210914 182868 210924
rect 184492 210898 184548 320460
rect 184604 263396 184660 403982
rect 184604 263330 184660 263340
rect 184716 403318 184772 403328
rect 184716 261156 184772 403262
rect 186284 402598 186340 402608
rect 186172 304836 186228 304846
rect 186060 294756 186116 294766
rect 185724 282212 185780 282222
rect 184716 261090 184772 261100
rect 185612 280532 185668 280542
rect 185612 265412 185668 280476
rect 185612 236628 185668 265356
rect 185724 268772 185780 282156
rect 185724 239204 185780 268716
rect 185948 280420 186004 280430
rect 185948 279188 186004 280364
rect 185948 239988 186004 279132
rect 185948 239922 186004 239932
rect 185724 239138 185780 239148
rect 185612 236562 185668 236572
rect 186060 212996 186116 294700
rect 186060 212930 186116 212940
rect 186172 211316 186228 304780
rect 186284 262276 186340 402542
rect 186396 381358 186452 550732
rect 187852 536452 187908 536462
rect 187740 514948 187796 514958
rect 186396 381292 186452 381302
rect 187068 471940 187124 471950
rect 186508 363076 186564 363086
rect 186508 359828 186564 363020
rect 186508 359762 186564 359772
rect 186620 361956 186676 361966
rect 186396 359716 186452 359726
rect 186396 349636 186452 359660
rect 186620 356468 186676 361900
rect 186620 356402 186676 356412
rect 186396 349570 186452 349580
rect 186284 262210 186340 262220
rect 186396 314916 186452 314926
rect 186172 211250 186228 211260
rect 184492 210832 184548 210842
rect 186396 209748 186452 314860
rect 186956 296996 187012 297006
rect 186956 211204 187012 296940
rect 187068 296548 187124 471884
rect 187292 450436 187348 450446
rect 187068 296482 187124 296492
rect 187180 300356 187236 300366
rect 187068 288838 187124 288848
rect 187068 287364 187124 288782
rect 187068 287298 187124 287308
rect 187068 286468 187124 286478
rect 187068 285778 187124 286412
rect 187068 285712 187124 285722
rect 187068 282100 187124 282110
rect 187068 260036 187124 282044
rect 187068 259970 187124 259980
rect 187180 239652 187236 300300
rect 187292 282212 187348 450380
rect 187292 282146 187348 282156
rect 187404 443268 187460 443278
rect 187404 280420 187460 443212
rect 187628 436100 187684 436110
rect 187404 280354 187460 280364
rect 187516 299236 187572 299246
rect 187404 255556 187460 255566
rect 187180 239586 187236 239596
rect 187292 254436 187348 254446
rect 187292 223076 187348 254380
rect 187292 223010 187348 223020
rect 187404 219268 187460 255500
rect 187516 219716 187572 299180
rect 187628 280532 187684 436044
rect 187740 407638 187796 514892
rect 187852 407818 187908 536396
rect 187852 407752 187908 407762
rect 187740 407572 187796 407582
rect 187964 397378 188020 565068
rect 189738 562350 190358 579922
rect 189738 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 190358 562350
rect 189738 562226 190358 562294
rect 189738 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 190358 562226
rect 189738 562102 190358 562170
rect 189738 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 190358 562102
rect 189738 561978 190358 562046
rect 189738 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 190358 561978
rect 189738 544350 190358 561922
rect 189738 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 190358 544350
rect 189738 544226 190358 544294
rect 189738 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 190358 544226
rect 189738 544102 190358 544170
rect 189738 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 190358 544102
rect 189738 543978 190358 544046
rect 189738 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 190358 543978
rect 189738 526350 190358 543922
rect 189738 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 190358 526350
rect 189738 526226 190358 526294
rect 189738 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 190358 526226
rect 189738 526102 190358 526170
rect 189738 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 190358 526102
rect 189738 525978 190358 526046
rect 189738 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 190358 525978
rect 189532 522116 189588 522126
rect 187964 397312 188020 397322
rect 189420 421764 189476 421774
rect 189420 392532 189476 421708
rect 189420 392466 189476 392476
rect 189532 390718 189588 522060
rect 189532 390652 189588 390662
rect 189738 508350 190358 525922
rect 189738 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 190358 508350
rect 189738 508226 190358 508294
rect 189738 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 190358 508226
rect 189738 508102 190358 508170
rect 189738 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 190358 508102
rect 189738 507978 190358 508046
rect 189738 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 190358 507978
rect 189738 490350 190358 507922
rect 189738 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 190358 490350
rect 189738 490226 190358 490294
rect 189738 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 190358 490226
rect 189738 490102 190358 490170
rect 189738 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 190358 490102
rect 189738 489978 190358 490046
rect 189738 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 190358 489978
rect 189738 472350 190358 489922
rect 189738 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 190358 472350
rect 189738 472226 190358 472294
rect 189738 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 190358 472226
rect 189738 472102 190358 472170
rect 189738 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 190358 472102
rect 189738 471978 190358 472046
rect 189738 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 190358 471978
rect 189738 454350 190358 471922
rect 189738 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 190358 454350
rect 189738 454226 190358 454294
rect 189738 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 190358 454226
rect 189738 454102 190358 454170
rect 189738 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 190358 454102
rect 189738 453978 190358 454046
rect 189738 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 190358 453978
rect 189738 436350 190358 453922
rect 189738 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 190358 436350
rect 189738 436226 190358 436294
rect 189738 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 190358 436226
rect 189738 436102 190358 436170
rect 189738 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 190358 436102
rect 189738 435978 190358 436046
rect 189738 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 190358 435978
rect 189738 418350 190358 435922
rect 189738 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 190358 418350
rect 189738 418226 190358 418294
rect 189738 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 190358 418226
rect 189738 418102 190358 418170
rect 189738 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 190358 418102
rect 189738 417978 190358 418046
rect 189738 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 190358 417978
rect 189738 400350 190358 417922
rect 189738 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 190358 400350
rect 189738 400226 190358 400294
rect 189738 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 190358 400226
rect 189738 400102 190358 400170
rect 189738 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 190358 400102
rect 189738 399978 190358 400046
rect 189738 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 190358 399978
rect 189738 382350 190358 399922
rect 189738 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 190358 382350
rect 189738 382226 190358 382294
rect 189738 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 190358 382226
rect 189738 382102 190358 382170
rect 189738 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 190358 382102
rect 189738 381978 190358 382046
rect 189738 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 190358 381978
rect 189738 364350 190358 381922
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 193458 586350 194078 597744
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 568350 194078 585922
rect 193458 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 194078 568350
rect 193458 568226 194078 568294
rect 193458 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 194078 568226
rect 193458 568102 194078 568170
rect 193458 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 194078 568102
rect 193458 567978 194078 568046
rect 193458 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 194078 567978
rect 193458 550350 194078 567922
rect 201516 591332 201572 591342
rect 194448 562350 194768 562384
rect 194448 562294 194518 562350
rect 194574 562294 194642 562350
rect 194698 562294 194768 562350
rect 194448 562226 194768 562294
rect 194448 562170 194518 562226
rect 194574 562170 194642 562226
rect 194698 562170 194768 562226
rect 194448 562102 194768 562170
rect 194448 562046 194518 562102
rect 194574 562046 194642 562102
rect 194698 562046 194768 562102
rect 194448 561978 194768 562046
rect 194448 561922 194518 561978
rect 194574 561922 194642 561978
rect 194698 561922 194768 561978
rect 194448 561888 194768 561922
rect 193458 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 194078 550350
rect 193458 550226 194078 550294
rect 193458 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 194078 550226
rect 193458 550102 194078 550170
rect 193458 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 194078 550102
rect 193458 549978 194078 550046
rect 193458 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 194078 549978
rect 193458 532350 194078 549922
rect 194448 544350 194768 544384
rect 194448 544294 194518 544350
rect 194574 544294 194642 544350
rect 194698 544294 194768 544350
rect 194448 544226 194768 544294
rect 194448 544170 194518 544226
rect 194574 544170 194642 544226
rect 194698 544170 194768 544226
rect 194448 544102 194768 544170
rect 194448 544046 194518 544102
rect 194574 544046 194642 544102
rect 194698 544046 194768 544102
rect 194448 543978 194768 544046
rect 194448 543922 194518 543978
rect 194574 543922 194642 543978
rect 194698 543922 194768 543978
rect 194448 543888 194768 543922
rect 193458 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 194078 532350
rect 193458 532226 194078 532294
rect 193458 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 194078 532226
rect 193458 532102 194078 532170
rect 193458 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 194078 532102
rect 193458 531978 194078 532046
rect 193458 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 194078 531978
rect 193458 514350 194078 531922
rect 194448 526350 194768 526384
rect 194448 526294 194518 526350
rect 194574 526294 194642 526350
rect 194698 526294 194768 526350
rect 194448 526226 194768 526294
rect 194448 526170 194518 526226
rect 194574 526170 194642 526226
rect 194698 526170 194768 526226
rect 194448 526102 194768 526170
rect 194448 526046 194518 526102
rect 194574 526046 194642 526102
rect 194698 526046 194768 526102
rect 194448 525978 194768 526046
rect 194448 525922 194518 525978
rect 194574 525922 194642 525978
rect 194698 525922 194768 525978
rect 194448 525888 194768 525922
rect 193458 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 194078 514350
rect 193458 514226 194078 514294
rect 193458 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 194078 514226
rect 193458 514102 194078 514170
rect 193458 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 194078 514102
rect 193458 513978 194078 514046
rect 193458 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 194078 513978
rect 193458 496350 194078 513922
rect 194448 508350 194768 508384
rect 194448 508294 194518 508350
rect 194574 508294 194642 508350
rect 194698 508294 194768 508350
rect 194448 508226 194768 508294
rect 194448 508170 194518 508226
rect 194574 508170 194642 508226
rect 194698 508170 194768 508226
rect 194448 508102 194768 508170
rect 194448 508046 194518 508102
rect 194574 508046 194642 508102
rect 194698 508046 194768 508102
rect 194448 507978 194768 508046
rect 194448 507922 194518 507978
rect 194574 507922 194642 507978
rect 194698 507922 194768 507978
rect 194448 507888 194768 507922
rect 193458 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 194078 496350
rect 193458 496226 194078 496294
rect 193458 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 194078 496226
rect 193458 496102 194078 496170
rect 193458 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 194078 496102
rect 193458 495978 194078 496046
rect 193458 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 194078 495978
rect 193458 478350 194078 495922
rect 194448 490350 194768 490384
rect 194448 490294 194518 490350
rect 194574 490294 194642 490350
rect 194698 490294 194768 490350
rect 194448 490226 194768 490294
rect 194448 490170 194518 490226
rect 194574 490170 194642 490226
rect 194698 490170 194768 490226
rect 194448 490102 194768 490170
rect 194448 490046 194518 490102
rect 194574 490046 194642 490102
rect 194698 490046 194768 490102
rect 194448 489978 194768 490046
rect 194448 489922 194518 489978
rect 194574 489922 194642 489978
rect 194698 489922 194768 489978
rect 194448 489888 194768 489922
rect 193458 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 194078 478350
rect 193458 478226 194078 478294
rect 193458 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 194078 478226
rect 193458 478102 194078 478170
rect 193458 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 194078 478102
rect 193458 477978 194078 478046
rect 193458 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 194078 477978
rect 193458 460350 194078 477922
rect 194448 472350 194768 472384
rect 194448 472294 194518 472350
rect 194574 472294 194642 472350
rect 194698 472294 194768 472350
rect 194448 472226 194768 472294
rect 194448 472170 194518 472226
rect 194574 472170 194642 472226
rect 194698 472170 194768 472226
rect 194448 472102 194768 472170
rect 194448 472046 194518 472102
rect 194574 472046 194642 472102
rect 194698 472046 194768 472102
rect 194448 471978 194768 472046
rect 194448 471922 194518 471978
rect 194574 471922 194642 471978
rect 194698 471922 194768 471978
rect 194448 471888 194768 471922
rect 193458 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 194078 460350
rect 193458 460226 194078 460294
rect 193458 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 194078 460226
rect 193458 460102 194078 460170
rect 193458 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 194078 460102
rect 193458 459978 194078 460046
rect 193458 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 194078 459978
rect 193458 442350 194078 459922
rect 194448 454350 194768 454384
rect 194448 454294 194518 454350
rect 194574 454294 194642 454350
rect 194698 454294 194768 454350
rect 194448 454226 194768 454294
rect 194448 454170 194518 454226
rect 194574 454170 194642 454226
rect 194698 454170 194768 454226
rect 194448 454102 194768 454170
rect 194448 454046 194518 454102
rect 194574 454046 194642 454102
rect 194698 454046 194768 454102
rect 194448 453978 194768 454046
rect 194448 453922 194518 453978
rect 194574 453922 194642 453978
rect 194698 453922 194768 453978
rect 194448 453888 194768 453922
rect 193458 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 194078 442350
rect 193458 442226 194078 442294
rect 193458 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 194078 442226
rect 193458 442102 194078 442170
rect 193458 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 194078 442102
rect 193458 441978 194078 442046
rect 193458 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 194078 441978
rect 193458 424350 194078 441922
rect 194448 436350 194768 436384
rect 194448 436294 194518 436350
rect 194574 436294 194642 436350
rect 194698 436294 194768 436350
rect 194448 436226 194768 436294
rect 194448 436170 194518 436226
rect 194574 436170 194642 436226
rect 194698 436170 194768 436226
rect 194448 436102 194768 436170
rect 194448 436046 194518 436102
rect 194574 436046 194642 436102
rect 194698 436046 194768 436102
rect 194448 435978 194768 436046
rect 194448 435922 194518 435978
rect 194574 435922 194642 435978
rect 194698 435922 194768 435978
rect 194448 435888 194768 435922
rect 193458 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 194078 424350
rect 193458 424226 194078 424294
rect 193458 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 194078 424226
rect 193458 424102 194078 424170
rect 193458 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 194078 424102
rect 193458 423978 194078 424046
rect 193458 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 194078 423978
rect 193458 406350 194078 423922
rect 194448 418350 194768 418384
rect 194448 418294 194518 418350
rect 194574 418294 194642 418350
rect 194698 418294 194768 418350
rect 194448 418226 194768 418294
rect 194448 418170 194518 418226
rect 194574 418170 194642 418226
rect 194698 418170 194768 418226
rect 194448 418102 194768 418170
rect 194448 418046 194518 418102
rect 194574 418046 194642 418102
rect 194698 418046 194768 418102
rect 194448 417978 194768 418046
rect 194448 417922 194518 417978
rect 194574 417922 194642 417978
rect 194698 417922 194768 417978
rect 194448 417888 194768 417922
rect 193458 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 194078 406350
rect 193458 406226 194078 406294
rect 193458 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 194078 406226
rect 193458 406102 194078 406170
rect 193458 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 194078 406102
rect 193458 405978 194078 406046
rect 193458 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 194078 405978
rect 193458 388350 194078 405922
rect 193458 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 194078 388350
rect 193458 388226 194078 388294
rect 193458 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 194078 388226
rect 193458 388102 194078 388170
rect 193458 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 194078 388102
rect 193458 387978 194078 388046
rect 193458 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 194078 387978
rect 193458 370350 194078 387922
rect 201404 401698 201460 401708
rect 201404 382452 201460 401642
rect 201516 395780 201572 591276
rect 203196 591220 203252 591230
rect 203196 395892 203252 591164
rect 208124 591108 208180 591118
rect 203196 395826 203252 395836
rect 204652 590996 204708 591006
rect 201516 395714 201572 395724
rect 203196 393778 203252 393788
rect 201404 382386 201460 382396
rect 203084 393418 203140 393428
rect 203084 382452 203140 393362
rect 203196 382564 203252 393722
rect 204652 392756 204708 590940
rect 208012 590884 208068 590894
rect 206332 590772 206388 590782
rect 204652 392690 204708 392700
rect 204764 393958 204820 393968
rect 203196 382498 203252 382508
rect 204764 382564 204820 393902
rect 204764 382498 204820 382508
rect 204876 393238 204932 393248
rect 203084 382386 203140 382396
rect 204876 382452 204932 393182
rect 206332 392868 206388 590716
rect 208012 408100 208068 590828
rect 208012 408034 208068 408044
rect 208124 407764 208180 591052
rect 208124 407698 208180 407708
rect 208236 590660 208292 590670
rect 206668 406756 206724 406766
rect 206332 392802 206388 392812
rect 206444 398278 206500 398288
rect 204876 382386 204932 382396
rect 206444 382452 206500 398222
rect 206556 393598 206612 393608
rect 206556 382564 206612 393542
rect 206556 382498 206612 382508
rect 206444 382386 206500 382396
rect 201292 379862 201460 379918
rect 201292 379764 201348 379862
rect 201292 379698 201348 379708
rect 193458 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 194078 370350
rect 193458 370226 194078 370294
rect 193458 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 194078 370226
rect 193458 370102 194078 370170
rect 193458 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 194078 370102
rect 193458 369978 194078 370046
rect 193458 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 194078 369978
rect 190652 368116 190708 368126
rect 190652 368038 190708 368060
rect 190652 367972 190708 367982
rect 190652 366996 190708 367006
rect 190652 366598 190708 366940
rect 190652 366532 190708 366542
rect 190652 366436 190708 366456
rect 190652 366352 190708 366362
rect 190652 364644 190708 364656
rect 190652 364552 190708 364562
rect 189738 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 190358 364350
rect 189738 364226 190358 364294
rect 189738 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 190358 364226
rect 189738 364102 190358 364170
rect 189738 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 190358 364102
rect 189738 363978 190358 364046
rect 189738 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 190358 363978
rect 189738 346350 190358 363922
rect 189738 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 190358 346350
rect 189738 346226 190358 346294
rect 189738 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 190358 346226
rect 189738 346102 190358 346170
rect 189738 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 190358 346102
rect 189738 345978 190358 346046
rect 189738 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 190358 345978
rect 189738 328350 190358 345922
rect 189738 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 190358 328350
rect 189738 328226 190358 328294
rect 189738 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 190358 328226
rect 189738 328102 190358 328170
rect 189738 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 190358 328102
rect 189738 327978 190358 328046
rect 189738 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 190358 327978
rect 189738 310350 190358 327922
rect 193458 352350 194078 369922
rect 194448 364350 194768 364384
rect 194448 364294 194518 364350
rect 194574 364294 194642 364350
rect 194698 364294 194768 364350
rect 194448 364226 194768 364294
rect 194448 364170 194518 364226
rect 194574 364170 194642 364226
rect 194698 364170 194768 364226
rect 194448 364102 194768 364170
rect 194448 364046 194518 364102
rect 194574 364046 194642 364102
rect 194698 364046 194768 364102
rect 194448 363978 194768 364046
rect 194448 363922 194518 363978
rect 194574 363922 194642 363978
rect 194698 363922 194768 363978
rect 194448 363888 194768 363922
rect 193458 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 194078 352350
rect 193458 352226 194078 352294
rect 193458 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 194078 352226
rect 193458 352102 194078 352170
rect 193458 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 194078 352102
rect 193458 351978 194078 352046
rect 193458 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 194078 351978
rect 193458 334350 194078 351922
rect 194448 346350 194768 346384
rect 194448 346294 194518 346350
rect 194574 346294 194642 346350
rect 194698 346294 194768 346350
rect 194448 346226 194768 346294
rect 194448 346170 194518 346226
rect 194574 346170 194642 346226
rect 194698 346170 194768 346226
rect 194448 346102 194768 346170
rect 194448 346046 194518 346102
rect 194574 346046 194642 346102
rect 194698 346046 194768 346102
rect 194448 345978 194768 346046
rect 194448 345922 194518 345978
rect 194574 345922 194642 345978
rect 194698 345922 194768 345978
rect 194448 345888 194768 345922
rect 193458 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 194078 334350
rect 193458 334226 194078 334294
rect 193458 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 194078 334226
rect 193458 334102 194078 334170
rect 193458 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 194078 334102
rect 193458 333978 194078 334046
rect 193458 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 194078 333978
rect 190652 319396 190708 319406
rect 190652 319258 190708 319340
rect 190652 319192 190708 319202
rect 193458 316350 194078 333922
rect 194448 328350 194768 328384
rect 194448 328294 194518 328350
rect 194574 328294 194642 328350
rect 194698 328294 194768 328350
rect 194448 328226 194768 328294
rect 194448 328170 194518 328226
rect 194574 328170 194642 328226
rect 194698 328170 194768 328226
rect 194448 328102 194768 328170
rect 194448 328046 194518 328102
rect 194574 328046 194642 328102
rect 194698 328046 194768 328102
rect 194448 327978 194768 328046
rect 194448 327922 194518 327978
rect 194574 327922 194642 327978
rect 194698 327922 194768 327978
rect 194448 327888 194768 327922
rect 193458 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 194078 316350
rect 193458 316226 194078 316294
rect 193458 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 194078 316226
rect 193458 316102 194078 316170
rect 193458 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 194078 316102
rect 193458 315978 194078 316046
rect 193458 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 194078 315978
rect 189738 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 190358 310350
rect 189738 310226 190358 310294
rect 189738 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 190358 310226
rect 189738 310102 190358 310170
rect 189738 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 190358 310102
rect 189738 309978 190358 310046
rect 189738 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 190358 309978
rect 189532 308196 189588 308206
rect 187628 280466 187684 280476
rect 187740 303716 187796 303726
rect 187516 219650 187572 219660
rect 187628 257796 187684 257806
rect 187404 219202 187460 219212
rect 187628 214564 187684 257740
rect 187740 221396 187796 303660
rect 187964 302596 188020 302606
rect 187740 221330 187796 221340
rect 187852 295876 187908 295886
rect 187628 214498 187684 214508
rect 187852 212884 187908 295820
rect 187852 212818 187908 212828
rect 187964 211428 188020 302540
rect 188076 289940 188132 289950
rect 188076 289018 188132 289884
rect 188076 288952 188132 288962
rect 188076 288148 188132 288158
rect 188076 287398 188132 288092
rect 188076 287332 188132 287342
rect 188076 286580 188132 286590
rect 188076 285958 188132 286524
rect 188076 285892 188132 285902
rect 188076 284788 188132 284798
rect 188076 283978 188132 284732
rect 188076 283912 188132 283922
rect 188076 280644 188132 280654
rect 188076 270658 188132 280588
rect 188076 270592 188132 270602
rect 187964 211362 188020 211372
rect 186956 211138 187012 211148
rect 189532 209860 189588 308140
rect 189738 292350 190358 309922
rect 189738 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 190358 292350
rect 189738 292226 190358 292294
rect 189738 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 190358 292226
rect 189738 292102 190358 292170
rect 189738 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 190358 292102
rect 189738 291978 190358 292046
rect 189738 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 190358 291978
rect 189738 274350 190358 291922
rect 189738 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 190358 274350
rect 189738 274226 190358 274294
rect 189738 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 190358 274226
rect 189738 274102 190358 274170
rect 189738 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 190358 274102
rect 189738 273978 190358 274046
rect 189738 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 190358 273978
rect 189738 256350 190358 273922
rect 189738 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 190358 256350
rect 189738 256226 190358 256294
rect 189738 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 190358 256226
rect 189738 256102 190358 256170
rect 189738 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 190358 256102
rect 189738 255978 190358 256046
rect 189738 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 190358 255978
rect 189738 238350 190358 255922
rect 189738 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 190358 238350
rect 189738 238226 190358 238294
rect 189738 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 190358 238226
rect 189738 238102 190358 238170
rect 189738 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 190358 238102
rect 189738 237978 190358 238046
rect 189738 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 190358 237978
rect 189738 220350 190358 237922
rect 190428 310436 190484 310446
rect 190428 224980 190484 310380
rect 193458 298350 194078 315922
rect 194448 310350 194768 310384
rect 194448 310294 194518 310350
rect 194574 310294 194642 310350
rect 194698 310294 194768 310350
rect 194448 310226 194768 310294
rect 194448 310170 194518 310226
rect 194574 310170 194642 310226
rect 194698 310170 194768 310226
rect 194448 310102 194768 310170
rect 194448 310046 194518 310102
rect 194574 310046 194642 310102
rect 194698 310046 194768 310102
rect 194448 309978 194768 310046
rect 194448 309922 194518 309978
rect 194574 309922 194642 309978
rect 194698 309922 194768 309978
rect 194448 309888 194768 309922
rect 193458 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 194078 298350
rect 193458 298226 194078 298294
rect 193458 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 194078 298226
rect 193458 298102 194078 298170
rect 193458 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 194078 298102
rect 193458 297978 194078 298046
rect 193458 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 194078 297978
rect 190652 293076 190708 293086
rect 190652 292618 190708 293020
rect 190652 292552 190708 292562
rect 193458 280350 194078 297922
rect 194448 292350 194768 292384
rect 194448 292294 194518 292350
rect 194574 292294 194642 292350
rect 194698 292294 194768 292350
rect 194448 292226 194768 292294
rect 194448 292170 194518 292226
rect 194574 292170 194642 292226
rect 194698 292170 194768 292226
rect 194448 292102 194768 292170
rect 194448 292046 194518 292102
rect 194574 292046 194642 292102
rect 194698 292046 194768 292102
rect 194448 291978 194768 292046
rect 194448 291922 194518 291978
rect 194574 291922 194642 291978
rect 194698 291922 194768 291978
rect 194448 291888 194768 291922
rect 193458 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 194078 280350
rect 193458 280226 194078 280294
rect 193458 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 194078 280226
rect 193458 280102 194078 280170
rect 193458 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 194078 280102
rect 193458 279978 194078 280046
rect 193458 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 194078 279978
rect 193458 262350 194078 279922
rect 194448 274350 194768 274384
rect 194448 274294 194518 274350
rect 194574 274294 194642 274350
rect 194698 274294 194768 274350
rect 194448 274226 194768 274294
rect 194448 274170 194518 274226
rect 194574 274170 194642 274226
rect 194698 274170 194768 274226
rect 194448 274102 194768 274170
rect 194448 274046 194518 274102
rect 194574 274046 194642 274102
rect 194698 274046 194768 274102
rect 194448 273978 194768 274046
rect 194448 273922 194518 273978
rect 194574 273922 194642 273978
rect 194698 273922 194768 273978
rect 194448 273888 194768 273922
rect 193458 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 194078 262350
rect 193458 262226 194078 262294
rect 193458 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 194078 262226
rect 193458 262102 194078 262170
rect 193458 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 194078 262102
rect 193458 261978 194078 262046
rect 193458 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 194078 261978
rect 190652 260398 190708 260408
rect 190652 259812 190708 260342
rect 190652 259746 190708 259756
rect 190652 255780 190708 255790
rect 190652 255538 190708 255724
rect 190652 255472 190708 255482
rect 190652 252420 190708 252430
rect 190652 252118 190708 252364
rect 190652 252052 190708 252062
rect 190428 224914 190484 224924
rect 193458 244350 194078 261922
rect 194448 256350 194768 256384
rect 194448 256294 194518 256350
rect 194574 256294 194642 256350
rect 194698 256294 194768 256350
rect 194448 256226 194768 256294
rect 194448 256170 194518 256226
rect 194574 256170 194642 256226
rect 194698 256170 194768 256226
rect 194448 256102 194768 256170
rect 194448 256046 194518 256102
rect 194574 256046 194642 256102
rect 194698 256046 194768 256102
rect 194448 255978 194768 256046
rect 194448 255922 194518 255978
rect 194574 255922 194642 255978
rect 194698 255922 194768 255978
rect 194448 255888 194768 255922
rect 193458 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 194078 244350
rect 193458 244226 194078 244294
rect 193458 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 194078 244226
rect 193458 244102 194078 244170
rect 193458 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 194078 244102
rect 193458 243978 194078 244046
rect 193458 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 194078 243978
rect 193458 226350 194078 243922
rect 193458 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 194078 226350
rect 193458 226226 194078 226294
rect 193458 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 194078 226226
rect 193458 226102 194078 226170
rect 193458 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 194078 226102
rect 193458 225978 194078 226046
rect 193458 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 194078 225978
rect 189738 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 190358 220350
rect 189738 220226 190358 220294
rect 189738 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 190358 220226
rect 189738 220102 190358 220170
rect 189738 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 190358 220102
rect 189738 219978 190358 220046
rect 189738 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 190358 219978
rect 189738 210574 190358 219922
rect 193458 210574 194078 225922
rect 201404 213108 201460 379862
rect 202860 379764 202916 379774
rect 202860 372988 202916 379708
rect 202860 372932 203252 372988
rect 203196 214676 203252 372932
rect 206668 340138 206724 406700
rect 208124 404218 208180 404228
rect 208124 382452 208180 404162
rect 208236 399140 208292 590604
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 209468 568708 209524 568718
rect 209468 407876 209524 568652
rect 220458 567550 221078 579922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 568350 224798 585922
rect 224178 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 224798 568350
rect 224178 568226 224798 568294
rect 224178 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 224798 568226
rect 224178 568102 224798 568170
rect 224178 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 224798 568102
rect 224178 567978 224798 568046
rect 224178 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 224798 567978
rect 224178 567550 224798 567922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 251178 567550 251798 579922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 568350 255518 585922
rect 254898 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 255518 568350
rect 254898 568226 255518 568294
rect 254898 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 255518 568226
rect 254898 568102 255518 568170
rect 254898 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 255518 568102
rect 254898 567978 255518 568046
rect 254898 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 255518 567978
rect 254898 567550 255518 567922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 281898 567550 282518 579922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 568350 286238 585922
rect 285618 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 286238 568350
rect 285618 568226 286238 568294
rect 285618 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 286238 568226
rect 285618 568102 286238 568170
rect 285618 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 286238 568102
rect 285618 567978 286238 568046
rect 285618 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 286238 567978
rect 285618 567550 286238 567922
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 312618 567550 313238 579922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 568350 316958 585922
rect 316338 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 316958 568350
rect 316338 568226 316958 568294
rect 316338 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 316958 568226
rect 316338 568102 316958 568170
rect 316338 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 316958 568102
rect 316338 567978 316958 568046
rect 316338 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 316958 567978
rect 316338 567550 316958 567922
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 343338 567550 343958 579922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 568350 347678 585922
rect 347058 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 347678 568350
rect 347058 568226 347678 568294
rect 347058 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 347678 568226
rect 347058 568102 347678 568170
rect 347058 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 347678 568102
rect 347058 567978 347678 568046
rect 347058 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 347678 567978
rect 347058 567550 347678 567922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 374058 567550 374678 579922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 568350 378398 585922
rect 377778 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 378398 568350
rect 377778 568226 378398 568294
rect 377778 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 378398 568226
rect 377778 568102 378398 568170
rect 377778 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 378398 568102
rect 377778 567978 378398 568046
rect 377778 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 378398 567978
rect 377778 567550 378398 567922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 404778 567550 405398 579922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 568350 409118 585922
rect 408498 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 409118 568350
rect 408498 568226 409118 568294
rect 408498 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 409118 568226
rect 408498 568102 409118 568170
rect 408498 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 409118 568102
rect 408498 567978 409118 568046
rect 408498 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 409118 567978
rect 408498 567550 409118 567922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 435498 567550 436118 579922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 568350 439838 585922
rect 439218 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 439838 568350
rect 439218 568226 439838 568294
rect 439218 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 439838 568226
rect 439218 568102 439838 568170
rect 439218 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 439838 568102
rect 439218 567978 439838 568046
rect 439218 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 439838 567978
rect 439218 567550 439838 567922
rect 444332 590212 444388 590222
rect 225168 562350 225488 562384
rect 225168 562294 225238 562350
rect 225294 562294 225362 562350
rect 225418 562294 225488 562350
rect 225168 562226 225488 562294
rect 225168 562170 225238 562226
rect 225294 562170 225362 562226
rect 225418 562170 225488 562226
rect 225168 562102 225488 562170
rect 225168 562046 225238 562102
rect 225294 562046 225362 562102
rect 225418 562046 225488 562102
rect 225168 561978 225488 562046
rect 225168 561922 225238 561978
rect 225294 561922 225362 561978
rect 225418 561922 225488 561978
rect 225168 561888 225488 561922
rect 255888 562350 256208 562384
rect 255888 562294 255958 562350
rect 256014 562294 256082 562350
rect 256138 562294 256208 562350
rect 255888 562226 256208 562294
rect 255888 562170 255958 562226
rect 256014 562170 256082 562226
rect 256138 562170 256208 562226
rect 255888 562102 256208 562170
rect 255888 562046 255958 562102
rect 256014 562046 256082 562102
rect 256138 562046 256208 562102
rect 255888 561978 256208 562046
rect 255888 561922 255958 561978
rect 256014 561922 256082 561978
rect 256138 561922 256208 561978
rect 255888 561888 256208 561922
rect 286608 562350 286928 562384
rect 286608 562294 286678 562350
rect 286734 562294 286802 562350
rect 286858 562294 286928 562350
rect 286608 562226 286928 562294
rect 286608 562170 286678 562226
rect 286734 562170 286802 562226
rect 286858 562170 286928 562226
rect 286608 562102 286928 562170
rect 286608 562046 286678 562102
rect 286734 562046 286802 562102
rect 286858 562046 286928 562102
rect 286608 561978 286928 562046
rect 286608 561922 286678 561978
rect 286734 561922 286802 561978
rect 286858 561922 286928 561978
rect 286608 561888 286928 561922
rect 317328 562350 317648 562384
rect 317328 562294 317398 562350
rect 317454 562294 317522 562350
rect 317578 562294 317648 562350
rect 317328 562226 317648 562294
rect 317328 562170 317398 562226
rect 317454 562170 317522 562226
rect 317578 562170 317648 562226
rect 317328 562102 317648 562170
rect 317328 562046 317398 562102
rect 317454 562046 317522 562102
rect 317578 562046 317648 562102
rect 317328 561978 317648 562046
rect 317328 561922 317398 561978
rect 317454 561922 317522 561978
rect 317578 561922 317648 561978
rect 317328 561888 317648 561922
rect 348048 562350 348368 562384
rect 348048 562294 348118 562350
rect 348174 562294 348242 562350
rect 348298 562294 348368 562350
rect 348048 562226 348368 562294
rect 348048 562170 348118 562226
rect 348174 562170 348242 562226
rect 348298 562170 348368 562226
rect 348048 562102 348368 562170
rect 348048 562046 348118 562102
rect 348174 562046 348242 562102
rect 348298 562046 348368 562102
rect 348048 561978 348368 562046
rect 348048 561922 348118 561978
rect 348174 561922 348242 561978
rect 348298 561922 348368 561978
rect 348048 561888 348368 561922
rect 378768 562350 379088 562384
rect 378768 562294 378838 562350
rect 378894 562294 378962 562350
rect 379018 562294 379088 562350
rect 378768 562226 379088 562294
rect 378768 562170 378838 562226
rect 378894 562170 378962 562226
rect 379018 562170 379088 562226
rect 378768 562102 379088 562170
rect 378768 562046 378838 562102
rect 378894 562046 378962 562102
rect 379018 562046 379088 562102
rect 378768 561978 379088 562046
rect 378768 561922 378838 561978
rect 378894 561922 378962 561978
rect 379018 561922 379088 561978
rect 378768 561888 379088 561922
rect 409488 562350 409808 562384
rect 409488 562294 409558 562350
rect 409614 562294 409682 562350
rect 409738 562294 409808 562350
rect 409488 562226 409808 562294
rect 409488 562170 409558 562226
rect 409614 562170 409682 562226
rect 409738 562170 409808 562226
rect 409488 562102 409808 562170
rect 409488 562046 409558 562102
rect 409614 562046 409682 562102
rect 409738 562046 409808 562102
rect 409488 561978 409808 562046
rect 409488 561922 409558 561978
rect 409614 561922 409682 561978
rect 409738 561922 409808 561978
rect 409488 561888 409808 561922
rect 440208 562350 440528 562384
rect 440208 562294 440278 562350
rect 440334 562294 440402 562350
rect 440458 562294 440528 562350
rect 440208 562226 440528 562294
rect 440208 562170 440278 562226
rect 440334 562170 440402 562226
rect 440458 562170 440528 562226
rect 440208 562102 440528 562170
rect 440208 562046 440278 562102
rect 440334 562046 440402 562102
rect 440458 562046 440528 562102
rect 440208 561978 440528 562046
rect 440208 561922 440278 561978
rect 440334 561922 440402 561978
rect 440458 561922 440528 561978
rect 440208 561888 440528 561922
rect 209808 550350 210128 550384
rect 209808 550294 209878 550350
rect 209934 550294 210002 550350
rect 210058 550294 210128 550350
rect 209808 550226 210128 550294
rect 209808 550170 209878 550226
rect 209934 550170 210002 550226
rect 210058 550170 210128 550226
rect 209808 550102 210128 550170
rect 209808 550046 209878 550102
rect 209934 550046 210002 550102
rect 210058 550046 210128 550102
rect 209808 549978 210128 550046
rect 209808 549922 209878 549978
rect 209934 549922 210002 549978
rect 210058 549922 210128 549978
rect 209808 549888 210128 549922
rect 240528 550350 240848 550384
rect 240528 550294 240598 550350
rect 240654 550294 240722 550350
rect 240778 550294 240848 550350
rect 240528 550226 240848 550294
rect 240528 550170 240598 550226
rect 240654 550170 240722 550226
rect 240778 550170 240848 550226
rect 240528 550102 240848 550170
rect 240528 550046 240598 550102
rect 240654 550046 240722 550102
rect 240778 550046 240848 550102
rect 240528 549978 240848 550046
rect 240528 549922 240598 549978
rect 240654 549922 240722 549978
rect 240778 549922 240848 549978
rect 240528 549888 240848 549922
rect 271248 550350 271568 550384
rect 271248 550294 271318 550350
rect 271374 550294 271442 550350
rect 271498 550294 271568 550350
rect 271248 550226 271568 550294
rect 271248 550170 271318 550226
rect 271374 550170 271442 550226
rect 271498 550170 271568 550226
rect 271248 550102 271568 550170
rect 271248 550046 271318 550102
rect 271374 550046 271442 550102
rect 271498 550046 271568 550102
rect 271248 549978 271568 550046
rect 271248 549922 271318 549978
rect 271374 549922 271442 549978
rect 271498 549922 271568 549978
rect 271248 549888 271568 549922
rect 301968 550350 302288 550384
rect 301968 550294 302038 550350
rect 302094 550294 302162 550350
rect 302218 550294 302288 550350
rect 301968 550226 302288 550294
rect 301968 550170 302038 550226
rect 302094 550170 302162 550226
rect 302218 550170 302288 550226
rect 301968 550102 302288 550170
rect 301968 550046 302038 550102
rect 302094 550046 302162 550102
rect 302218 550046 302288 550102
rect 301968 549978 302288 550046
rect 301968 549922 302038 549978
rect 302094 549922 302162 549978
rect 302218 549922 302288 549978
rect 301968 549888 302288 549922
rect 332688 550350 333008 550384
rect 332688 550294 332758 550350
rect 332814 550294 332882 550350
rect 332938 550294 333008 550350
rect 332688 550226 333008 550294
rect 332688 550170 332758 550226
rect 332814 550170 332882 550226
rect 332938 550170 333008 550226
rect 332688 550102 333008 550170
rect 332688 550046 332758 550102
rect 332814 550046 332882 550102
rect 332938 550046 333008 550102
rect 332688 549978 333008 550046
rect 332688 549922 332758 549978
rect 332814 549922 332882 549978
rect 332938 549922 333008 549978
rect 332688 549888 333008 549922
rect 363408 550350 363728 550384
rect 363408 550294 363478 550350
rect 363534 550294 363602 550350
rect 363658 550294 363728 550350
rect 363408 550226 363728 550294
rect 363408 550170 363478 550226
rect 363534 550170 363602 550226
rect 363658 550170 363728 550226
rect 363408 550102 363728 550170
rect 363408 550046 363478 550102
rect 363534 550046 363602 550102
rect 363658 550046 363728 550102
rect 363408 549978 363728 550046
rect 363408 549922 363478 549978
rect 363534 549922 363602 549978
rect 363658 549922 363728 549978
rect 363408 549888 363728 549922
rect 394128 550350 394448 550384
rect 394128 550294 394198 550350
rect 394254 550294 394322 550350
rect 394378 550294 394448 550350
rect 394128 550226 394448 550294
rect 394128 550170 394198 550226
rect 394254 550170 394322 550226
rect 394378 550170 394448 550226
rect 394128 550102 394448 550170
rect 394128 550046 394198 550102
rect 394254 550046 394322 550102
rect 394378 550046 394448 550102
rect 394128 549978 394448 550046
rect 394128 549922 394198 549978
rect 394254 549922 394322 549978
rect 394378 549922 394448 549978
rect 394128 549888 394448 549922
rect 424848 550350 425168 550384
rect 424848 550294 424918 550350
rect 424974 550294 425042 550350
rect 425098 550294 425168 550350
rect 424848 550226 425168 550294
rect 424848 550170 424918 550226
rect 424974 550170 425042 550226
rect 425098 550170 425168 550226
rect 424848 550102 425168 550170
rect 424848 550046 424918 550102
rect 424974 550046 425042 550102
rect 425098 550046 425168 550102
rect 424848 549978 425168 550046
rect 424848 549922 424918 549978
rect 424974 549922 425042 549978
rect 425098 549922 425168 549978
rect 424848 549888 425168 549922
rect 225168 544350 225488 544384
rect 225168 544294 225238 544350
rect 225294 544294 225362 544350
rect 225418 544294 225488 544350
rect 225168 544226 225488 544294
rect 225168 544170 225238 544226
rect 225294 544170 225362 544226
rect 225418 544170 225488 544226
rect 225168 544102 225488 544170
rect 225168 544046 225238 544102
rect 225294 544046 225362 544102
rect 225418 544046 225488 544102
rect 225168 543978 225488 544046
rect 225168 543922 225238 543978
rect 225294 543922 225362 543978
rect 225418 543922 225488 543978
rect 225168 543888 225488 543922
rect 255888 544350 256208 544384
rect 255888 544294 255958 544350
rect 256014 544294 256082 544350
rect 256138 544294 256208 544350
rect 255888 544226 256208 544294
rect 255888 544170 255958 544226
rect 256014 544170 256082 544226
rect 256138 544170 256208 544226
rect 255888 544102 256208 544170
rect 255888 544046 255958 544102
rect 256014 544046 256082 544102
rect 256138 544046 256208 544102
rect 255888 543978 256208 544046
rect 255888 543922 255958 543978
rect 256014 543922 256082 543978
rect 256138 543922 256208 543978
rect 255888 543888 256208 543922
rect 286608 544350 286928 544384
rect 286608 544294 286678 544350
rect 286734 544294 286802 544350
rect 286858 544294 286928 544350
rect 286608 544226 286928 544294
rect 286608 544170 286678 544226
rect 286734 544170 286802 544226
rect 286858 544170 286928 544226
rect 286608 544102 286928 544170
rect 286608 544046 286678 544102
rect 286734 544046 286802 544102
rect 286858 544046 286928 544102
rect 286608 543978 286928 544046
rect 286608 543922 286678 543978
rect 286734 543922 286802 543978
rect 286858 543922 286928 543978
rect 286608 543888 286928 543922
rect 317328 544350 317648 544384
rect 317328 544294 317398 544350
rect 317454 544294 317522 544350
rect 317578 544294 317648 544350
rect 317328 544226 317648 544294
rect 317328 544170 317398 544226
rect 317454 544170 317522 544226
rect 317578 544170 317648 544226
rect 317328 544102 317648 544170
rect 317328 544046 317398 544102
rect 317454 544046 317522 544102
rect 317578 544046 317648 544102
rect 317328 543978 317648 544046
rect 317328 543922 317398 543978
rect 317454 543922 317522 543978
rect 317578 543922 317648 543978
rect 317328 543888 317648 543922
rect 348048 544350 348368 544384
rect 348048 544294 348118 544350
rect 348174 544294 348242 544350
rect 348298 544294 348368 544350
rect 348048 544226 348368 544294
rect 348048 544170 348118 544226
rect 348174 544170 348242 544226
rect 348298 544170 348368 544226
rect 348048 544102 348368 544170
rect 348048 544046 348118 544102
rect 348174 544046 348242 544102
rect 348298 544046 348368 544102
rect 348048 543978 348368 544046
rect 348048 543922 348118 543978
rect 348174 543922 348242 543978
rect 348298 543922 348368 543978
rect 348048 543888 348368 543922
rect 378768 544350 379088 544384
rect 378768 544294 378838 544350
rect 378894 544294 378962 544350
rect 379018 544294 379088 544350
rect 378768 544226 379088 544294
rect 378768 544170 378838 544226
rect 378894 544170 378962 544226
rect 379018 544170 379088 544226
rect 378768 544102 379088 544170
rect 378768 544046 378838 544102
rect 378894 544046 378962 544102
rect 379018 544046 379088 544102
rect 378768 543978 379088 544046
rect 378768 543922 378838 543978
rect 378894 543922 378962 543978
rect 379018 543922 379088 543978
rect 378768 543888 379088 543922
rect 409488 544350 409808 544384
rect 409488 544294 409558 544350
rect 409614 544294 409682 544350
rect 409738 544294 409808 544350
rect 409488 544226 409808 544294
rect 409488 544170 409558 544226
rect 409614 544170 409682 544226
rect 409738 544170 409808 544226
rect 409488 544102 409808 544170
rect 409488 544046 409558 544102
rect 409614 544046 409682 544102
rect 409738 544046 409808 544102
rect 409488 543978 409808 544046
rect 409488 543922 409558 543978
rect 409614 543922 409682 543978
rect 409738 543922 409808 543978
rect 409488 543888 409808 543922
rect 440208 544350 440528 544384
rect 440208 544294 440278 544350
rect 440334 544294 440402 544350
rect 440458 544294 440528 544350
rect 440208 544226 440528 544294
rect 440208 544170 440278 544226
rect 440334 544170 440402 544226
rect 440458 544170 440528 544226
rect 440208 544102 440528 544170
rect 440208 544046 440278 544102
rect 440334 544046 440402 544102
rect 440458 544046 440528 544102
rect 440208 543978 440528 544046
rect 440208 543922 440278 543978
rect 440334 543922 440402 543978
rect 440458 543922 440528 543978
rect 440208 543888 440528 543922
rect 209808 532350 210128 532384
rect 209808 532294 209878 532350
rect 209934 532294 210002 532350
rect 210058 532294 210128 532350
rect 209808 532226 210128 532294
rect 209808 532170 209878 532226
rect 209934 532170 210002 532226
rect 210058 532170 210128 532226
rect 209808 532102 210128 532170
rect 209808 532046 209878 532102
rect 209934 532046 210002 532102
rect 210058 532046 210128 532102
rect 209808 531978 210128 532046
rect 209808 531922 209878 531978
rect 209934 531922 210002 531978
rect 210058 531922 210128 531978
rect 209808 531888 210128 531922
rect 240528 532350 240848 532384
rect 240528 532294 240598 532350
rect 240654 532294 240722 532350
rect 240778 532294 240848 532350
rect 240528 532226 240848 532294
rect 240528 532170 240598 532226
rect 240654 532170 240722 532226
rect 240778 532170 240848 532226
rect 240528 532102 240848 532170
rect 240528 532046 240598 532102
rect 240654 532046 240722 532102
rect 240778 532046 240848 532102
rect 240528 531978 240848 532046
rect 240528 531922 240598 531978
rect 240654 531922 240722 531978
rect 240778 531922 240848 531978
rect 240528 531888 240848 531922
rect 271248 532350 271568 532384
rect 271248 532294 271318 532350
rect 271374 532294 271442 532350
rect 271498 532294 271568 532350
rect 271248 532226 271568 532294
rect 271248 532170 271318 532226
rect 271374 532170 271442 532226
rect 271498 532170 271568 532226
rect 271248 532102 271568 532170
rect 271248 532046 271318 532102
rect 271374 532046 271442 532102
rect 271498 532046 271568 532102
rect 271248 531978 271568 532046
rect 271248 531922 271318 531978
rect 271374 531922 271442 531978
rect 271498 531922 271568 531978
rect 271248 531888 271568 531922
rect 301968 532350 302288 532384
rect 301968 532294 302038 532350
rect 302094 532294 302162 532350
rect 302218 532294 302288 532350
rect 301968 532226 302288 532294
rect 301968 532170 302038 532226
rect 302094 532170 302162 532226
rect 302218 532170 302288 532226
rect 301968 532102 302288 532170
rect 301968 532046 302038 532102
rect 302094 532046 302162 532102
rect 302218 532046 302288 532102
rect 301968 531978 302288 532046
rect 301968 531922 302038 531978
rect 302094 531922 302162 531978
rect 302218 531922 302288 531978
rect 301968 531888 302288 531922
rect 332688 532350 333008 532384
rect 332688 532294 332758 532350
rect 332814 532294 332882 532350
rect 332938 532294 333008 532350
rect 332688 532226 333008 532294
rect 332688 532170 332758 532226
rect 332814 532170 332882 532226
rect 332938 532170 333008 532226
rect 332688 532102 333008 532170
rect 332688 532046 332758 532102
rect 332814 532046 332882 532102
rect 332938 532046 333008 532102
rect 332688 531978 333008 532046
rect 332688 531922 332758 531978
rect 332814 531922 332882 531978
rect 332938 531922 333008 531978
rect 332688 531888 333008 531922
rect 363408 532350 363728 532384
rect 363408 532294 363478 532350
rect 363534 532294 363602 532350
rect 363658 532294 363728 532350
rect 363408 532226 363728 532294
rect 363408 532170 363478 532226
rect 363534 532170 363602 532226
rect 363658 532170 363728 532226
rect 363408 532102 363728 532170
rect 363408 532046 363478 532102
rect 363534 532046 363602 532102
rect 363658 532046 363728 532102
rect 363408 531978 363728 532046
rect 363408 531922 363478 531978
rect 363534 531922 363602 531978
rect 363658 531922 363728 531978
rect 363408 531888 363728 531922
rect 394128 532350 394448 532384
rect 394128 532294 394198 532350
rect 394254 532294 394322 532350
rect 394378 532294 394448 532350
rect 394128 532226 394448 532294
rect 394128 532170 394198 532226
rect 394254 532170 394322 532226
rect 394378 532170 394448 532226
rect 394128 532102 394448 532170
rect 394128 532046 394198 532102
rect 394254 532046 394322 532102
rect 394378 532046 394448 532102
rect 394128 531978 394448 532046
rect 394128 531922 394198 531978
rect 394254 531922 394322 531978
rect 394378 531922 394448 531978
rect 394128 531888 394448 531922
rect 424848 532350 425168 532384
rect 424848 532294 424918 532350
rect 424974 532294 425042 532350
rect 425098 532294 425168 532350
rect 424848 532226 425168 532294
rect 424848 532170 424918 532226
rect 424974 532170 425042 532226
rect 425098 532170 425168 532226
rect 424848 532102 425168 532170
rect 424848 532046 424918 532102
rect 424974 532046 425042 532102
rect 425098 532046 425168 532102
rect 424848 531978 425168 532046
rect 424848 531922 424918 531978
rect 424974 531922 425042 531978
rect 425098 531922 425168 531978
rect 424848 531888 425168 531922
rect 225168 526350 225488 526384
rect 225168 526294 225238 526350
rect 225294 526294 225362 526350
rect 225418 526294 225488 526350
rect 225168 526226 225488 526294
rect 225168 526170 225238 526226
rect 225294 526170 225362 526226
rect 225418 526170 225488 526226
rect 225168 526102 225488 526170
rect 225168 526046 225238 526102
rect 225294 526046 225362 526102
rect 225418 526046 225488 526102
rect 225168 525978 225488 526046
rect 225168 525922 225238 525978
rect 225294 525922 225362 525978
rect 225418 525922 225488 525978
rect 225168 525888 225488 525922
rect 255888 526350 256208 526384
rect 255888 526294 255958 526350
rect 256014 526294 256082 526350
rect 256138 526294 256208 526350
rect 255888 526226 256208 526294
rect 255888 526170 255958 526226
rect 256014 526170 256082 526226
rect 256138 526170 256208 526226
rect 255888 526102 256208 526170
rect 255888 526046 255958 526102
rect 256014 526046 256082 526102
rect 256138 526046 256208 526102
rect 255888 525978 256208 526046
rect 255888 525922 255958 525978
rect 256014 525922 256082 525978
rect 256138 525922 256208 525978
rect 255888 525888 256208 525922
rect 286608 526350 286928 526384
rect 286608 526294 286678 526350
rect 286734 526294 286802 526350
rect 286858 526294 286928 526350
rect 286608 526226 286928 526294
rect 286608 526170 286678 526226
rect 286734 526170 286802 526226
rect 286858 526170 286928 526226
rect 286608 526102 286928 526170
rect 286608 526046 286678 526102
rect 286734 526046 286802 526102
rect 286858 526046 286928 526102
rect 286608 525978 286928 526046
rect 286608 525922 286678 525978
rect 286734 525922 286802 525978
rect 286858 525922 286928 525978
rect 286608 525888 286928 525922
rect 317328 526350 317648 526384
rect 317328 526294 317398 526350
rect 317454 526294 317522 526350
rect 317578 526294 317648 526350
rect 317328 526226 317648 526294
rect 317328 526170 317398 526226
rect 317454 526170 317522 526226
rect 317578 526170 317648 526226
rect 317328 526102 317648 526170
rect 317328 526046 317398 526102
rect 317454 526046 317522 526102
rect 317578 526046 317648 526102
rect 317328 525978 317648 526046
rect 317328 525922 317398 525978
rect 317454 525922 317522 525978
rect 317578 525922 317648 525978
rect 317328 525888 317648 525922
rect 348048 526350 348368 526384
rect 348048 526294 348118 526350
rect 348174 526294 348242 526350
rect 348298 526294 348368 526350
rect 348048 526226 348368 526294
rect 348048 526170 348118 526226
rect 348174 526170 348242 526226
rect 348298 526170 348368 526226
rect 348048 526102 348368 526170
rect 348048 526046 348118 526102
rect 348174 526046 348242 526102
rect 348298 526046 348368 526102
rect 348048 525978 348368 526046
rect 348048 525922 348118 525978
rect 348174 525922 348242 525978
rect 348298 525922 348368 525978
rect 348048 525888 348368 525922
rect 378768 526350 379088 526384
rect 378768 526294 378838 526350
rect 378894 526294 378962 526350
rect 379018 526294 379088 526350
rect 378768 526226 379088 526294
rect 378768 526170 378838 526226
rect 378894 526170 378962 526226
rect 379018 526170 379088 526226
rect 378768 526102 379088 526170
rect 378768 526046 378838 526102
rect 378894 526046 378962 526102
rect 379018 526046 379088 526102
rect 378768 525978 379088 526046
rect 378768 525922 378838 525978
rect 378894 525922 378962 525978
rect 379018 525922 379088 525978
rect 378768 525888 379088 525922
rect 409488 526350 409808 526384
rect 409488 526294 409558 526350
rect 409614 526294 409682 526350
rect 409738 526294 409808 526350
rect 409488 526226 409808 526294
rect 409488 526170 409558 526226
rect 409614 526170 409682 526226
rect 409738 526170 409808 526226
rect 409488 526102 409808 526170
rect 409488 526046 409558 526102
rect 409614 526046 409682 526102
rect 409738 526046 409808 526102
rect 409488 525978 409808 526046
rect 409488 525922 409558 525978
rect 409614 525922 409682 525978
rect 409738 525922 409808 525978
rect 409488 525888 409808 525922
rect 440208 526350 440528 526384
rect 440208 526294 440278 526350
rect 440334 526294 440402 526350
rect 440458 526294 440528 526350
rect 440208 526226 440528 526294
rect 440208 526170 440278 526226
rect 440334 526170 440402 526226
rect 440458 526170 440528 526226
rect 440208 526102 440528 526170
rect 440208 526046 440278 526102
rect 440334 526046 440402 526102
rect 440458 526046 440528 526102
rect 440208 525978 440528 526046
rect 440208 525922 440278 525978
rect 440334 525922 440402 525978
rect 440458 525922 440528 525978
rect 440208 525888 440528 525922
rect 209808 514350 210128 514384
rect 209808 514294 209878 514350
rect 209934 514294 210002 514350
rect 210058 514294 210128 514350
rect 209808 514226 210128 514294
rect 209808 514170 209878 514226
rect 209934 514170 210002 514226
rect 210058 514170 210128 514226
rect 209808 514102 210128 514170
rect 209808 514046 209878 514102
rect 209934 514046 210002 514102
rect 210058 514046 210128 514102
rect 209808 513978 210128 514046
rect 209808 513922 209878 513978
rect 209934 513922 210002 513978
rect 210058 513922 210128 513978
rect 209808 513888 210128 513922
rect 240528 514350 240848 514384
rect 240528 514294 240598 514350
rect 240654 514294 240722 514350
rect 240778 514294 240848 514350
rect 240528 514226 240848 514294
rect 240528 514170 240598 514226
rect 240654 514170 240722 514226
rect 240778 514170 240848 514226
rect 240528 514102 240848 514170
rect 240528 514046 240598 514102
rect 240654 514046 240722 514102
rect 240778 514046 240848 514102
rect 240528 513978 240848 514046
rect 240528 513922 240598 513978
rect 240654 513922 240722 513978
rect 240778 513922 240848 513978
rect 240528 513888 240848 513922
rect 271248 514350 271568 514384
rect 271248 514294 271318 514350
rect 271374 514294 271442 514350
rect 271498 514294 271568 514350
rect 271248 514226 271568 514294
rect 271248 514170 271318 514226
rect 271374 514170 271442 514226
rect 271498 514170 271568 514226
rect 271248 514102 271568 514170
rect 271248 514046 271318 514102
rect 271374 514046 271442 514102
rect 271498 514046 271568 514102
rect 271248 513978 271568 514046
rect 271248 513922 271318 513978
rect 271374 513922 271442 513978
rect 271498 513922 271568 513978
rect 271248 513888 271568 513922
rect 301968 514350 302288 514384
rect 301968 514294 302038 514350
rect 302094 514294 302162 514350
rect 302218 514294 302288 514350
rect 301968 514226 302288 514294
rect 301968 514170 302038 514226
rect 302094 514170 302162 514226
rect 302218 514170 302288 514226
rect 301968 514102 302288 514170
rect 301968 514046 302038 514102
rect 302094 514046 302162 514102
rect 302218 514046 302288 514102
rect 301968 513978 302288 514046
rect 301968 513922 302038 513978
rect 302094 513922 302162 513978
rect 302218 513922 302288 513978
rect 301968 513888 302288 513922
rect 332688 514350 333008 514384
rect 332688 514294 332758 514350
rect 332814 514294 332882 514350
rect 332938 514294 333008 514350
rect 332688 514226 333008 514294
rect 332688 514170 332758 514226
rect 332814 514170 332882 514226
rect 332938 514170 333008 514226
rect 332688 514102 333008 514170
rect 332688 514046 332758 514102
rect 332814 514046 332882 514102
rect 332938 514046 333008 514102
rect 332688 513978 333008 514046
rect 332688 513922 332758 513978
rect 332814 513922 332882 513978
rect 332938 513922 333008 513978
rect 332688 513888 333008 513922
rect 363408 514350 363728 514384
rect 363408 514294 363478 514350
rect 363534 514294 363602 514350
rect 363658 514294 363728 514350
rect 363408 514226 363728 514294
rect 363408 514170 363478 514226
rect 363534 514170 363602 514226
rect 363658 514170 363728 514226
rect 363408 514102 363728 514170
rect 363408 514046 363478 514102
rect 363534 514046 363602 514102
rect 363658 514046 363728 514102
rect 363408 513978 363728 514046
rect 363408 513922 363478 513978
rect 363534 513922 363602 513978
rect 363658 513922 363728 513978
rect 363408 513888 363728 513922
rect 394128 514350 394448 514384
rect 394128 514294 394198 514350
rect 394254 514294 394322 514350
rect 394378 514294 394448 514350
rect 394128 514226 394448 514294
rect 394128 514170 394198 514226
rect 394254 514170 394322 514226
rect 394378 514170 394448 514226
rect 394128 514102 394448 514170
rect 394128 514046 394198 514102
rect 394254 514046 394322 514102
rect 394378 514046 394448 514102
rect 394128 513978 394448 514046
rect 394128 513922 394198 513978
rect 394254 513922 394322 513978
rect 394378 513922 394448 513978
rect 394128 513888 394448 513922
rect 424848 514350 425168 514384
rect 424848 514294 424918 514350
rect 424974 514294 425042 514350
rect 425098 514294 425168 514350
rect 424848 514226 425168 514294
rect 424848 514170 424918 514226
rect 424974 514170 425042 514226
rect 425098 514170 425168 514226
rect 424848 514102 425168 514170
rect 424848 514046 424918 514102
rect 424974 514046 425042 514102
rect 425098 514046 425168 514102
rect 424848 513978 425168 514046
rect 424848 513922 424918 513978
rect 424974 513922 425042 513978
rect 425098 513922 425168 513978
rect 424848 513888 425168 513922
rect 225168 508350 225488 508384
rect 225168 508294 225238 508350
rect 225294 508294 225362 508350
rect 225418 508294 225488 508350
rect 225168 508226 225488 508294
rect 225168 508170 225238 508226
rect 225294 508170 225362 508226
rect 225418 508170 225488 508226
rect 225168 508102 225488 508170
rect 225168 508046 225238 508102
rect 225294 508046 225362 508102
rect 225418 508046 225488 508102
rect 225168 507978 225488 508046
rect 225168 507922 225238 507978
rect 225294 507922 225362 507978
rect 225418 507922 225488 507978
rect 225168 507888 225488 507922
rect 255888 508350 256208 508384
rect 255888 508294 255958 508350
rect 256014 508294 256082 508350
rect 256138 508294 256208 508350
rect 255888 508226 256208 508294
rect 255888 508170 255958 508226
rect 256014 508170 256082 508226
rect 256138 508170 256208 508226
rect 255888 508102 256208 508170
rect 255888 508046 255958 508102
rect 256014 508046 256082 508102
rect 256138 508046 256208 508102
rect 255888 507978 256208 508046
rect 255888 507922 255958 507978
rect 256014 507922 256082 507978
rect 256138 507922 256208 507978
rect 255888 507888 256208 507922
rect 286608 508350 286928 508384
rect 286608 508294 286678 508350
rect 286734 508294 286802 508350
rect 286858 508294 286928 508350
rect 286608 508226 286928 508294
rect 286608 508170 286678 508226
rect 286734 508170 286802 508226
rect 286858 508170 286928 508226
rect 286608 508102 286928 508170
rect 286608 508046 286678 508102
rect 286734 508046 286802 508102
rect 286858 508046 286928 508102
rect 286608 507978 286928 508046
rect 286608 507922 286678 507978
rect 286734 507922 286802 507978
rect 286858 507922 286928 507978
rect 286608 507888 286928 507922
rect 317328 508350 317648 508384
rect 317328 508294 317398 508350
rect 317454 508294 317522 508350
rect 317578 508294 317648 508350
rect 317328 508226 317648 508294
rect 317328 508170 317398 508226
rect 317454 508170 317522 508226
rect 317578 508170 317648 508226
rect 317328 508102 317648 508170
rect 317328 508046 317398 508102
rect 317454 508046 317522 508102
rect 317578 508046 317648 508102
rect 317328 507978 317648 508046
rect 317328 507922 317398 507978
rect 317454 507922 317522 507978
rect 317578 507922 317648 507978
rect 317328 507888 317648 507922
rect 348048 508350 348368 508384
rect 348048 508294 348118 508350
rect 348174 508294 348242 508350
rect 348298 508294 348368 508350
rect 348048 508226 348368 508294
rect 348048 508170 348118 508226
rect 348174 508170 348242 508226
rect 348298 508170 348368 508226
rect 348048 508102 348368 508170
rect 348048 508046 348118 508102
rect 348174 508046 348242 508102
rect 348298 508046 348368 508102
rect 348048 507978 348368 508046
rect 348048 507922 348118 507978
rect 348174 507922 348242 507978
rect 348298 507922 348368 507978
rect 348048 507888 348368 507922
rect 378768 508350 379088 508384
rect 378768 508294 378838 508350
rect 378894 508294 378962 508350
rect 379018 508294 379088 508350
rect 378768 508226 379088 508294
rect 378768 508170 378838 508226
rect 378894 508170 378962 508226
rect 379018 508170 379088 508226
rect 378768 508102 379088 508170
rect 378768 508046 378838 508102
rect 378894 508046 378962 508102
rect 379018 508046 379088 508102
rect 378768 507978 379088 508046
rect 378768 507922 378838 507978
rect 378894 507922 378962 507978
rect 379018 507922 379088 507978
rect 378768 507888 379088 507922
rect 409488 508350 409808 508384
rect 409488 508294 409558 508350
rect 409614 508294 409682 508350
rect 409738 508294 409808 508350
rect 409488 508226 409808 508294
rect 409488 508170 409558 508226
rect 409614 508170 409682 508226
rect 409738 508170 409808 508226
rect 409488 508102 409808 508170
rect 409488 508046 409558 508102
rect 409614 508046 409682 508102
rect 409738 508046 409808 508102
rect 409488 507978 409808 508046
rect 409488 507922 409558 507978
rect 409614 507922 409682 507978
rect 409738 507922 409808 507978
rect 409488 507888 409808 507922
rect 440208 508350 440528 508384
rect 440208 508294 440278 508350
rect 440334 508294 440402 508350
rect 440458 508294 440528 508350
rect 440208 508226 440528 508294
rect 440208 508170 440278 508226
rect 440334 508170 440402 508226
rect 440458 508170 440528 508226
rect 440208 508102 440528 508170
rect 440208 508046 440278 508102
rect 440334 508046 440402 508102
rect 440458 508046 440528 508102
rect 440208 507978 440528 508046
rect 440208 507922 440278 507978
rect 440334 507922 440402 507978
rect 440458 507922 440528 507978
rect 440208 507888 440528 507922
rect 209808 496350 210128 496384
rect 209808 496294 209878 496350
rect 209934 496294 210002 496350
rect 210058 496294 210128 496350
rect 209808 496226 210128 496294
rect 209808 496170 209878 496226
rect 209934 496170 210002 496226
rect 210058 496170 210128 496226
rect 209808 496102 210128 496170
rect 209808 496046 209878 496102
rect 209934 496046 210002 496102
rect 210058 496046 210128 496102
rect 209808 495978 210128 496046
rect 209808 495922 209878 495978
rect 209934 495922 210002 495978
rect 210058 495922 210128 495978
rect 209808 495888 210128 495922
rect 240528 496350 240848 496384
rect 240528 496294 240598 496350
rect 240654 496294 240722 496350
rect 240778 496294 240848 496350
rect 240528 496226 240848 496294
rect 240528 496170 240598 496226
rect 240654 496170 240722 496226
rect 240778 496170 240848 496226
rect 240528 496102 240848 496170
rect 240528 496046 240598 496102
rect 240654 496046 240722 496102
rect 240778 496046 240848 496102
rect 240528 495978 240848 496046
rect 240528 495922 240598 495978
rect 240654 495922 240722 495978
rect 240778 495922 240848 495978
rect 240528 495888 240848 495922
rect 271248 496350 271568 496384
rect 271248 496294 271318 496350
rect 271374 496294 271442 496350
rect 271498 496294 271568 496350
rect 271248 496226 271568 496294
rect 271248 496170 271318 496226
rect 271374 496170 271442 496226
rect 271498 496170 271568 496226
rect 271248 496102 271568 496170
rect 271248 496046 271318 496102
rect 271374 496046 271442 496102
rect 271498 496046 271568 496102
rect 271248 495978 271568 496046
rect 271248 495922 271318 495978
rect 271374 495922 271442 495978
rect 271498 495922 271568 495978
rect 271248 495888 271568 495922
rect 301968 496350 302288 496384
rect 301968 496294 302038 496350
rect 302094 496294 302162 496350
rect 302218 496294 302288 496350
rect 301968 496226 302288 496294
rect 301968 496170 302038 496226
rect 302094 496170 302162 496226
rect 302218 496170 302288 496226
rect 301968 496102 302288 496170
rect 301968 496046 302038 496102
rect 302094 496046 302162 496102
rect 302218 496046 302288 496102
rect 301968 495978 302288 496046
rect 301968 495922 302038 495978
rect 302094 495922 302162 495978
rect 302218 495922 302288 495978
rect 301968 495888 302288 495922
rect 332688 496350 333008 496384
rect 332688 496294 332758 496350
rect 332814 496294 332882 496350
rect 332938 496294 333008 496350
rect 332688 496226 333008 496294
rect 332688 496170 332758 496226
rect 332814 496170 332882 496226
rect 332938 496170 333008 496226
rect 332688 496102 333008 496170
rect 332688 496046 332758 496102
rect 332814 496046 332882 496102
rect 332938 496046 333008 496102
rect 332688 495978 333008 496046
rect 332688 495922 332758 495978
rect 332814 495922 332882 495978
rect 332938 495922 333008 495978
rect 332688 495888 333008 495922
rect 363408 496350 363728 496384
rect 363408 496294 363478 496350
rect 363534 496294 363602 496350
rect 363658 496294 363728 496350
rect 363408 496226 363728 496294
rect 363408 496170 363478 496226
rect 363534 496170 363602 496226
rect 363658 496170 363728 496226
rect 363408 496102 363728 496170
rect 363408 496046 363478 496102
rect 363534 496046 363602 496102
rect 363658 496046 363728 496102
rect 363408 495978 363728 496046
rect 363408 495922 363478 495978
rect 363534 495922 363602 495978
rect 363658 495922 363728 495978
rect 363408 495888 363728 495922
rect 394128 496350 394448 496384
rect 394128 496294 394198 496350
rect 394254 496294 394322 496350
rect 394378 496294 394448 496350
rect 394128 496226 394448 496294
rect 394128 496170 394198 496226
rect 394254 496170 394322 496226
rect 394378 496170 394448 496226
rect 394128 496102 394448 496170
rect 394128 496046 394198 496102
rect 394254 496046 394322 496102
rect 394378 496046 394448 496102
rect 394128 495978 394448 496046
rect 394128 495922 394198 495978
rect 394254 495922 394322 495978
rect 394378 495922 394448 495978
rect 394128 495888 394448 495922
rect 424848 496350 425168 496384
rect 424848 496294 424918 496350
rect 424974 496294 425042 496350
rect 425098 496294 425168 496350
rect 424848 496226 425168 496294
rect 424848 496170 424918 496226
rect 424974 496170 425042 496226
rect 425098 496170 425168 496226
rect 424848 496102 425168 496170
rect 424848 496046 424918 496102
rect 424974 496046 425042 496102
rect 425098 496046 425168 496102
rect 424848 495978 425168 496046
rect 424848 495922 424918 495978
rect 424974 495922 425042 495978
rect 425098 495922 425168 495978
rect 424848 495888 425168 495922
rect 225168 490350 225488 490384
rect 225168 490294 225238 490350
rect 225294 490294 225362 490350
rect 225418 490294 225488 490350
rect 225168 490226 225488 490294
rect 225168 490170 225238 490226
rect 225294 490170 225362 490226
rect 225418 490170 225488 490226
rect 225168 490102 225488 490170
rect 225168 490046 225238 490102
rect 225294 490046 225362 490102
rect 225418 490046 225488 490102
rect 225168 489978 225488 490046
rect 225168 489922 225238 489978
rect 225294 489922 225362 489978
rect 225418 489922 225488 489978
rect 225168 489888 225488 489922
rect 255888 490350 256208 490384
rect 255888 490294 255958 490350
rect 256014 490294 256082 490350
rect 256138 490294 256208 490350
rect 255888 490226 256208 490294
rect 255888 490170 255958 490226
rect 256014 490170 256082 490226
rect 256138 490170 256208 490226
rect 255888 490102 256208 490170
rect 255888 490046 255958 490102
rect 256014 490046 256082 490102
rect 256138 490046 256208 490102
rect 255888 489978 256208 490046
rect 255888 489922 255958 489978
rect 256014 489922 256082 489978
rect 256138 489922 256208 489978
rect 255888 489888 256208 489922
rect 286608 490350 286928 490384
rect 286608 490294 286678 490350
rect 286734 490294 286802 490350
rect 286858 490294 286928 490350
rect 286608 490226 286928 490294
rect 286608 490170 286678 490226
rect 286734 490170 286802 490226
rect 286858 490170 286928 490226
rect 286608 490102 286928 490170
rect 286608 490046 286678 490102
rect 286734 490046 286802 490102
rect 286858 490046 286928 490102
rect 286608 489978 286928 490046
rect 286608 489922 286678 489978
rect 286734 489922 286802 489978
rect 286858 489922 286928 489978
rect 286608 489888 286928 489922
rect 317328 490350 317648 490384
rect 317328 490294 317398 490350
rect 317454 490294 317522 490350
rect 317578 490294 317648 490350
rect 317328 490226 317648 490294
rect 317328 490170 317398 490226
rect 317454 490170 317522 490226
rect 317578 490170 317648 490226
rect 317328 490102 317648 490170
rect 317328 490046 317398 490102
rect 317454 490046 317522 490102
rect 317578 490046 317648 490102
rect 317328 489978 317648 490046
rect 317328 489922 317398 489978
rect 317454 489922 317522 489978
rect 317578 489922 317648 489978
rect 317328 489888 317648 489922
rect 348048 490350 348368 490384
rect 348048 490294 348118 490350
rect 348174 490294 348242 490350
rect 348298 490294 348368 490350
rect 348048 490226 348368 490294
rect 348048 490170 348118 490226
rect 348174 490170 348242 490226
rect 348298 490170 348368 490226
rect 348048 490102 348368 490170
rect 348048 490046 348118 490102
rect 348174 490046 348242 490102
rect 348298 490046 348368 490102
rect 348048 489978 348368 490046
rect 348048 489922 348118 489978
rect 348174 489922 348242 489978
rect 348298 489922 348368 489978
rect 348048 489888 348368 489922
rect 378768 490350 379088 490384
rect 378768 490294 378838 490350
rect 378894 490294 378962 490350
rect 379018 490294 379088 490350
rect 378768 490226 379088 490294
rect 378768 490170 378838 490226
rect 378894 490170 378962 490226
rect 379018 490170 379088 490226
rect 378768 490102 379088 490170
rect 378768 490046 378838 490102
rect 378894 490046 378962 490102
rect 379018 490046 379088 490102
rect 378768 489978 379088 490046
rect 378768 489922 378838 489978
rect 378894 489922 378962 489978
rect 379018 489922 379088 489978
rect 378768 489888 379088 489922
rect 409488 490350 409808 490384
rect 409488 490294 409558 490350
rect 409614 490294 409682 490350
rect 409738 490294 409808 490350
rect 409488 490226 409808 490294
rect 409488 490170 409558 490226
rect 409614 490170 409682 490226
rect 409738 490170 409808 490226
rect 409488 490102 409808 490170
rect 409488 490046 409558 490102
rect 409614 490046 409682 490102
rect 409738 490046 409808 490102
rect 409488 489978 409808 490046
rect 409488 489922 409558 489978
rect 409614 489922 409682 489978
rect 409738 489922 409808 489978
rect 409488 489888 409808 489922
rect 440208 490350 440528 490384
rect 440208 490294 440278 490350
rect 440334 490294 440402 490350
rect 440458 490294 440528 490350
rect 440208 490226 440528 490294
rect 440208 490170 440278 490226
rect 440334 490170 440402 490226
rect 440458 490170 440528 490226
rect 440208 490102 440528 490170
rect 440208 490046 440278 490102
rect 440334 490046 440402 490102
rect 440458 490046 440528 490102
rect 440208 489978 440528 490046
rect 440208 489922 440278 489978
rect 440334 489922 440402 489978
rect 440458 489922 440528 489978
rect 440208 489888 440528 489922
rect 209808 478350 210128 478384
rect 209808 478294 209878 478350
rect 209934 478294 210002 478350
rect 210058 478294 210128 478350
rect 209808 478226 210128 478294
rect 209808 478170 209878 478226
rect 209934 478170 210002 478226
rect 210058 478170 210128 478226
rect 209808 478102 210128 478170
rect 209808 478046 209878 478102
rect 209934 478046 210002 478102
rect 210058 478046 210128 478102
rect 209808 477978 210128 478046
rect 209808 477922 209878 477978
rect 209934 477922 210002 477978
rect 210058 477922 210128 477978
rect 209808 477888 210128 477922
rect 240528 478350 240848 478384
rect 240528 478294 240598 478350
rect 240654 478294 240722 478350
rect 240778 478294 240848 478350
rect 240528 478226 240848 478294
rect 240528 478170 240598 478226
rect 240654 478170 240722 478226
rect 240778 478170 240848 478226
rect 240528 478102 240848 478170
rect 240528 478046 240598 478102
rect 240654 478046 240722 478102
rect 240778 478046 240848 478102
rect 240528 477978 240848 478046
rect 240528 477922 240598 477978
rect 240654 477922 240722 477978
rect 240778 477922 240848 477978
rect 240528 477888 240848 477922
rect 271248 478350 271568 478384
rect 271248 478294 271318 478350
rect 271374 478294 271442 478350
rect 271498 478294 271568 478350
rect 271248 478226 271568 478294
rect 271248 478170 271318 478226
rect 271374 478170 271442 478226
rect 271498 478170 271568 478226
rect 271248 478102 271568 478170
rect 271248 478046 271318 478102
rect 271374 478046 271442 478102
rect 271498 478046 271568 478102
rect 271248 477978 271568 478046
rect 271248 477922 271318 477978
rect 271374 477922 271442 477978
rect 271498 477922 271568 477978
rect 271248 477888 271568 477922
rect 301968 478350 302288 478384
rect 301968 478294 302038 478350
rect 302094 478294 302162 478350
rect 302218 478294 302288 478350
rect 301968 478226 302288 478294
rect 301968 478170 302038 478226
rect 302094 478170 302162 478226
rect 302218 478170 302288 478226
rect 301968 478102 302288 478170
rect 301968 478046 302038 478102
rect 302094 478046 302162 478102
rect 302218 478046 302288 478102
rect 301968 477978 302288 478046
rect 301968 477922 302038 477978
rect 302094 477922 302162 477978
rect 302218 477922 302288 477978
rect 301968 477888 302288 477922
rect 332688 478350 333008 478384
rect 332688 478294 332758 478350
rect 332814 478294 332882 478350
rect 332938 478294 333008 478350
rect 332688 478226 333008 478294
rect 332688 478170 332758 478226
rect 332814 478170 332882 478226
rect 332938 478170 333008 478226
rect 332688 478102 333008 478170
rect 332688 478046 332758 478102
rect 332814 478046 332882 478102
rect 332938 478046 333008 478102
rect 332688 477978 333008 478046
rect 332688 477922 332758 477978
rect 332814 477922 332882 477978
rect 332938 477922 333008 477978
rect 332688 477888 333008 477922
rect 363408 478350 363728 478384
rect 363408 478294 363478 478350
rect 363534 478294 363602 478350
rect 363658 478294 363728 478350
rect 363408 478226 363728 478294
rect 363408 478170 363478 478226
rect 363534 478170 363602 478226
rect 363658 478170 363728 478226
rect 363408 478102 363728 478170
rect 363408 478046 363478 478102
rect 363534 478046 363602 478102
rect 363658 478046 363728 478102
rect 363408 477978 363728 478046
rect 363408 477922 363478 477978
rect 363534 477922 363602 477978
rect 363658 477922 363728 477978
rect 363408 477888 363728 477922
rect 394128 478350 394448 478384
rect 394128 478294 394198 478350
rect 394254 478294 394322 478350
rect 394378 478294 394448 478350
rect 394128 478226 394448 478294
rect 394128 478170 394198 478226
rect 394254 478170 394322 478226
rect 394378 478170 394448 478226
rect 394128 478102 394448 478170
rect 394128 478046 394198 478102
rect 394254 478046 394322 478102
rect 394378 478046 394448 478102
rect 394128 477978 394448 478046
rect 394128 477922 394198 477978
rect 394254 477922 394322 477978
rect 394378 477922 394448 477978
rect 394128 477888 394448 477922
rect 424848 478350 425168 478384
rect 424848 478294 424918 478350
rect 424974 478294 425042 478350
rect 425098 478294 425168 478350
rect 424848 478226 425168 478294
rect 424848 478170 424918 478226
rect 424974 478170 425042 478226
rect 425098 478170 425168 478226
rect 424848 478102 425168 478170
rect 424848 478046 424918 478102
rect 424974 478046 425042 478102
rect 425098 478046 425168 478102
rect 424848 477978 425168 478046
rect 424848 477922 424918 477978
rect 424974 477922 425042 477978
rect 425098 477922 425168 477978
rect 424848 477888 425168 477922
rect 225168 472350 225488 472384
rect 225168 472294 225238 472350
rect 225294 472294 225362 472350
rect 225418 472294 225488 472350
rect 225168 472226 225488 472294
rect 225168 472170 225238 472226
rect 225294 472170 225362 472226
rect 225418 472170 225488 472226
rect 225168 472102 225488 472170
rect 225168 472046 225238 472102
rect 225294 472046 225362 472102
rect 225418 472046 225488 472102
rect 225168 471978 225488 472046
rect 225168 471922 225238 471978
rect 225294 471922 225362 471978
rect 225418 471922 225488 471978
rect 225168 471888 225488 471922
rect 255888 472350 256208 472384
rect 255888 472294 255958 472350
rect 256014 472294 256082 472350
rect 256138 472294 256208 472350
rect 255888 472226 256208 472294
rect 255888 472170 255958 472226
rect 256014 472170 256082 472226
rect 256138 472170 256208 472226
rect 255888 472102 256208 472170
rect 255888 472046 255958 472102
rect 256014 472046 256082 472102
rect 256138 472046 256208 472102
rect 255888 471978 256208 472046
rect 255888 471922 255958 471978
rect 256014 471922 256082 471978
rect 256138 471922 256208 471978
rect 255888 471888 256208 471922
rect 286608 472350 286928 472384
rect 286608 472294 286678 472350
rect 286734 472294 286802 472350
rect 286858 472294 286928 472350
rect 286608 472226 286928 472294
rect 286608 472170 286678 472226
rect 286734 472170 286802 472226
rect 286858 472170 286928 472226
rect 286608 472102 286928 472170
rect 286608 472046 286678 472102
rect 286734 472046 286802 472102
rect 286858 472046 286928 472102
rect 286608 471978 286928 472046
rect 286608 471922 286678 471978
rect 286734 471922 286802 471978
rect 286858 471922 286928 471978
rect 286608 471888 286928 471922
rect 317328 472350 317648 472384
rect 317328 472294 317398 472350
rect 317454 472294 317522 472350
rect 317578 472294 317648 472350
rect 317328 472226 317648 472294
rect 317328 472170 317398 472226
rect 317454 472170 317522 472226
rect 317578 472170 317648 472226
rect 317328 472102 317648 472170
rect 317328 472046 317398 472102
rect 317454 472046 317522 472102
rect 317578 472046 317648 472102
rect 317328 471978 317648 472046
rect 317328 471922 317398 471978
rect 317454 471922 317522 471978
rect 317578 471922 317648 471978
rect 317328 471888 317648 471922
rect 348048 472350 348368 472384
rect 348048 472294 348118 472350
rect 348174 472294 348242 472350
rect 348298 472294 348368 472350
rect 348048 472226 348368 472294
rect 348048 472170 348118 472226
rect 348174 472170 348242 472226
rect 348298 472170 348368 472226
rect 348048 472102 348368 472170
rect 348048 472046 348118 472102
rect 348174 472046 348242 472102
rect 348298 472046 348368 472102
rect 348048 471978 348368 472046
rect 348048 471922 348118 471978
rect 348174 471922 348242 471978
rect 348298 471922 348368 471978
rect 348048 471888 348368 471922
rect 378768 472350 379088 472384
rect 378768 472294 378838 472350
rect 378894 472294 378962 472350
rect 379018 472294 379088 472350
rect 378768 472226 379088 472294
rect 378768 472170 378838 472226
rect 378894 472170 378962 472226
rect 379018 472170 379088 472226
rect 378768 472102 379088 472170
rect 378768 472046 378838 472102
rect 378894 472046 378962 472102
rect 379018 472046 379088 472102
rect 378768 471978 379088 472046
rect 378768 471922 378838 471978
rect 378894 471922 378962 471978
rect 379018 471922 379088 471978
rect 378768 471888 379088 471922
rect 409488 472350 409808 472384
rect 409488 472294 409558 472350
rect 409614 472294 409682 472350
rect 409738 472294 409808 472350
rect 409488 472226 409808 472294
rect 409488 472170 409558 472226
rect 409614 472170 409682 472226
rect 409738 472170 409808 472226
rect 409488 472102 409808 472170
rect 409488 472046 409558 472102
rect 409614 472046 409682 472102
rect 409738 472046 409808 472102
rect 409488 471978 409808 472046
rect 409488 471922 409558 471978
rect 409614 471922 409682 471978
rect 409738 471922 409808 471978
rect 409488 471888 409808 471922
rect 440208 472350 440528 472384
rect 440208 472294 440278 472350
rect 440334 472294 440402 472350
rect 440458 472294 440528 472350
rect 440208 472226 440528 472294
rect 440208 472170 440278 472226
rect 440334 472170 440402 472226
rect 440458 472170 440528 472226
rect 440208 472102 440528 472170
rect 440208 472046 440278 472102
rect 440334 472046 440402 472102
rect 440458 472046 440528 472102
rect 440208 471978 440528 472046
rect 440208 471922 440278 471978
rect 440334 471922 440402 471978
rect 440458 471922 440528 471978
rect 440208 471888 440528 471922
rect 209808 460350 210128 460384
rect 209808 460294 209878 460350
rect 209934 460294 210002 460350
rect 210058 460294 210128 460350
rect 209808 460226 210128 460294
rect 209808 460170 209878 460226
rect 209934 460170 210002 460226
rect 210058 460170 210128 460226
rect 209808 460102 210128 460170
rect 209808 460046 209878 460102
rect 209934 460046 210002 460102
rect 210058 460046 210128 460102
rect 209808 459978 210128 460046
rect 209808 459922 209878 459978
rect 209934 459922 210002 459978
rect 210058 459922 210128 459978
rect 209808 459888 210128 459922
rect 240528 460350 240848 460384
rect 240528 460294 240598 460350
rect 240654 460294 240722 460350
rect 240778 460294 240848 460350
rect 240528 460226 240848 460294
rect 240528 460170 240598 460226
rect 240654 460170 240722 460226
rect 240778 460170 240848 460226
rect 240528 460102 240848 460170
rect 240528 460046 240598 460102
rect 240654 460046 240722 460102
rect 240778 460046 240848 460102
rect 240528 459978 240848 460046
rect 240528 459922 240598 459978
rect 240654 459922 240722 459978
rect 240778 459922 240848 459978
rect 240528 459888 240848 459922
rect 271248 460350 271568 460384
rect 271248 460294 271318 460350
rect 271374 460294 271442 460350
rect 271498 460294 271568 460350
rect 271248 460226 271568 460294
rect 271248 460170 271318 460226
rect 271374 460170 271442 460226
rect 271498 460170 271568 460226
rect 271248 460102 271568 460170
rect 271248 460046 271318 460102
rect 271374 460046 271442 460102
rect 271498 460046 271568 460102
rect 271248 459978 271568 460046
rect 271248 459922 271318 459978
rect 271374 459922 271442 459978
rect 271498 459922 271568 459978
rect 271248 459888 271568 459922
rect 301968 460350 302288 460384
rect 301968 460294 302038 460350
rect 302094 460294 302162 460350
rect 302218 460294 302288 460350
rect 301968 460226 302288 460294
rect 301968 460170 302038 460226
rect 302094 460170 302162 460226
rect 302218 460170 302288 460226
rect 301968 460102 302288 460170
rect 301968 460046 302038 460102
rect 302094 460046 302162 460102
rect 302218 460046 302288 460102
rect 301968 459978 302288 460046
rect 301968 459922 302038 459978
rect 302094 459922 302162 459978
rect 302218 459922 302288 459978
rect 301968 459888 302288 459922
rect 332688 460350 333008 460384
rect 332688 460294 332758 460350
rect 332814 460294 332882 460350
rect 332938 460294 333008 460350
rect 332688 460226 333008 460294
rect 332688 460170 332758 460226
rect 332814 460170 332882 460226
rect 332938 460170 333008 460226
rect 332688 460102 333008 460170
rect 332688 460046 332758 460102
rect 332814 460046 332882 460102
rect 332938 460046 333008 460102
rect 332688 459978 333008 460046
rect 332688 459922 332758 459978
rect 332814 459922 332882 459978
rect 332938 459922 333008 459978
rect 332688 459888 333008 459922
rect 363408 460350 363728 460384
rect 363408 460294 363478 460350
rect 363534 460294 363602 460350
rect 363658 460294 363728 460350
rect 363408 460226 363728 460294
rect 363408 460170 363478 460226
rect 363534 460170 363602 460226
rect 363658 460170 363728 460226
rect 363408 460102 363728 460170
rect 363408 460046 363478 460102
rect 363534 460046 363602 460102
rect 363658 460046 363728 460102
rect 363408 459978 363728 460046
rect 363408 459922 363478 459978
rect 363534 459922 363602 459978
rect 363658 459922 363728 459978
rect 363408 459888 363728 459922
rect 394128 460350 394448 460384
rect 394128 460294 394198 460350
rect 394254 460294 394322 460350
rect 394378 460294 394448 460350
rect 394128 460226 394448 460294
rect 394128 460170 394198 460226
rect 394254 460170 394322 460226
rect 394378 460170 394448 460226
rect 394128 460102 394448 460170
rect 394128 460046 394198 460102
rect 394254 460046 394322 460102
rect 394378 460046 394448 460102
rect 394128 459978 394448 460046
rect 394128 459922 394198 459978
rect 394254 459922 394322 459978
rect 394378 459922 394448 459978
rect 394128 459888 394448 459922
rect 424848 460350 425168 460384
rect 424848 460294 424918 460350
rect 424974 460294 425042 460350
rect 425098 460294 425168 460350
rect 424848 460226 425168 460294
rect 424848 460170 424918 460226
rect 424974 460170 425042 460226
rect 425098 460170 425168 460226
rect 424848 460102 425168 460170
rect 424848 460046 424918 460102
rect 424974 460046 425042 460102
rect 425098 460046 425168 460102
rect 424848 459978 425168 460046
rect 424848 459922 424918 459978
rect 424974 459922 425042 459978
rect 425098 459922 425168 459978
rect 424848 459888 425168 459922
rect 225168 454350 225488 454384
rect 225168 454294 225238 454350
rect 225294 454294 225362 454350
rect 225418 454294 225488 454350
rect 225168 454226 225488 454294
rect 225168 454170 225238 454226
rect 225294 454170 225362 454226
rect 225418 454170 225488 454226
rect 225168 454102 225488 454170
rect 225168 454046 225238 454102
rect 225294 454046 225362 454102
rect 225418 454046 225488 454102
rect 225168 453978 225488 454046
rect 225168 453922 225238 453978
rect 225294 453922 225362 453978
rect 225418 453922 225488 453978
rect 225168 453888 225488 453922
rect 255888 454350 256208 454384
rect 255888 454294 255958 454350
rect 256014 454294 256082 454350
rect 256138 454294 256208 454350
rect 255888 454226 256208 454294
rect 255888 454170 255958 454226
rect 256014 454170 256082 454226
rect 256138 454170 256208 454226
rect 255888 454102 256208 454170
rect 255888 454046 255958 454102
rect 256014 454046 256082 454102
rect 256138 454046 256208 454102
rect 255888 453978 256208 454046
rect 255888 453922 255958 453978
rect 256014 453922 256082 453978
rect 256138 453922 256208 453978
rect 255888 453888 256208 453922
rect 286608 454350 286928 454384
rect 286608 454294 286678 454350
rect 286734 454294 286802 454350
rect 286858 454294 286928 454350
rect 286608 454226 286928 454294
rect 286608 454170 286678 454226
rect 286734 454170 286802 454226
rect 286858 454170 286928 454226
rect 286608 454102 286928 454170
rect 286608 454046 286678 454102
rect 286734 454046 286802 454102
rect 286858 454046 286928 454102
rect 286608 453978 286928 454046
rect 286608 453922 286678 453978
rect 286734 453922 286802 453978
rect 286858 453922 286928 453978
rect 286608 453888 286928 453922
rect 317328 454350 317648 454384
rect 317328 454294 317398 454350
rect 317454 454294 317522 454350
rect 317578 454294 317648 454350
rect 317328 454226 317648 454294
rect 317328 454170 317398 454226
rect 317454 454170 317522 454226
rect 317578 454170 317648 454226
rect 317328 454102 317648 454170
rect 317328 454046 317398 454102
rect 317454 454046 317522 454102
rect 317578 454046 317648 454102
rect 317328 453978 317648 454046
rect 317328 453922 317398 453978
rect 317454 453922 317522 453978
rect 317578 453922 317648 453978
rect 317328 453888 317648 453922
rect 348048 454350 348368 454384
rect 348048 454294 348118 454350
rect 348174 454294 348242 454350
rect 348298 454294 348368 454350
rect 348048 454226 348368 454294
rect 348048 454170 348118 454226
rect 348174 454170 348242 454226
rect 348298 454170 348368 454226
rect 348048 454102 348368 454170
rect 348048 454046 348118 454102
rect 348174 454046 348242 454102
rect 348298 454046 348368 454102
rect 348048 453978 348368 454046
rect 348048 453922 348118 453978
rect 348174 453922 348242 453978
rect 348298 453922 348368 453978
rect 348048 453888 348368 453922
rect 378768 454350 379088 454384
rect 378768 454294 378838 454350
rect 378894 454294 378962 454350
rect 379018 454294 379088 454350
rect 378768 454226 379088 454294
rect 378768 454170 378838 454226
rect 378894 454170 378962 454226
rect 379018 454170 379088 454226
rect 378768 454102 379088 454170
rect 378768 454046 378838 454102
rect 378894 454046 378962 454102
rect 379018 454046 379088 454102
rect 378768 453978 379088 454046
rect 378768 453922 378838 453978
rect 378894 453922 378962 453978
rect 379018 453922 379088 453978
rect 378768 453888 379088 453922
rect 409488 454350 409808 454384
rect 409488 454294 409558 454350
rect 409614 454294 409682 454350
rect 409738 454294 409808 454350
rect 409488 454226 409808 454294
rect 409488 454170 409558 454226
rect 409614 454170 409682 454226
rect 409738 454170 409808 454226
rect 409488 454102 409808 454170
rect 409488 454046 409558 454102
rect 409614 454046 409682 454102
rect 409738 454046 409808 454102
rect 409488 453978 409808 454046
rect 409488 453922 409558 453978
rect 409614 453922 409682 453978
rect 409738 453922 409808 453978
rect 409488 453888 409808 453922
rect 440208 454350 440528 454384
rect 440208 454294 440278 454350
rect 440334 454294 440402 454350
rect 440458 454294 440528 454350
rect 440208 454226 440528 454294
rect 440208 454170 440278 454226
rect 440334 454170 440402 454226
rect 440458 454170 440528 454226
rect 440208 454102 440528 454170
rect 440208 454046 440278 454102
rect 440334 454046 440402 454102
rect 440458 454046 440528 454102
rect 440208 453978 440528 454046
rect 440208 453922 440278 453978
rect 440334 453922 440402 453978
rect 440458 453922 440528 453978
rect 440208 453888 440528 453922
rect 209808 442350 210128 442384
rect 209808 442294 209878 442350
rect 209934 442294 210002 442350
rect 210058 442294 210128 442350
rect 209808 442226 210128 442294
rect 209808 442170 209878 442226
rect 209934 442170 210002 442226
rect 210058 442170 210128 442226
rect 209808 442102 210128 442170
rect 209808 442046 209878 442102
rect 209934 442046 210002 442102
rect 210058 442046 210128 442102
rect 209808 441978 210128 442046
rect 209808 441922 209878 441978
rect 209934 441922 210002 441978
rect 210058 441922 210128 441978
rect 209808 441888 210128 441922
rect 240528 442350 240848 442384
rect 240528 442294 240598 442350
rect 240654 442294 240722 442350
rect 240778 442294 240848 442350
rect 240528 442226 240848 442294
rect 240528 442170 240598 442226
rect 240654 442170 240722 442226
rect 240778 442170 240848 442226
rect 240528 442102 240848 442170
rect 240528 442046 240598 442102
rect 240654 442046 240722 442102
rect 240778 442046 240848 442102
rect 240528 441978 240848 442046
rect 240528 441922 240598 441978
rect 240654 441922 240722 441978
rect 240778 441922 240848 441978
rect 240528 441888 240848 441922
rect 271248 442350 271568 442384
rect 271248 442294 271318 442350
rect 271374 442294 271442 442350
rect 271498 442294 271568 442350
rect 271248 442226 271568 442294
rect 271248 442170 271318 442226
rect 271374 442170 271442 442226
rect 271498 442170 271568 442226
rect 271248 442102 271568 442170
rect 271248 442046 271318 442102
rect 271374 442046 271442 442102
rect 271498 442046 271568 442102
rect 271248 441978 271568 442046
rect 271248 441922 271318 441978
rect 271374 441922 271442 441978
rect 271498 441922 271568 441978
rect 271248 441888 271568 441922
rect 301968 442350 302288 442384
rect 301968 442294 302038 442350
rect 302094 442294 302162 442350
rect 302218 442294 302288 442350
rect 301968 442226 302288 442294
rect 301968 442170 302038 442226
rect 302094 442170 302162 442226
rect 302218 442170 302288 442226
rect 301968 442102 302288 442170
rect 301968 442046 302038 442102
rect 302094 442046 302162 442102
rect 302218 442046 302288 442102
rect 301968 441978 302288 442046
rect 301968 441922 302038 441978
rect 302094 441922 302162 441978
rect 302218 441922 302288 441978
rect 301968 441888 302288 441922
rect 332688 442350 333008 442384
rect 332688 442294 332758 442350
rect 332814 442294 332882 442350
rect 332938 442294 333008 442350
rect 332688 442226 333008 442294
rect 332688 442170 332758 442226
rect 332814 442170 332882 442226
rect 332938 442170 333008 442226
rect 332688 442102 333008 442170
rect 332688 442046 332758 442102
rect 332814 442046 332882 442102
rect 332938 442046 333008 442102
rect 332688 441978 333008 442046
rect 332688 441922 332758 441978
rect 332814 441922 332882 441978
rect 332938 441922 333008 441978
rect 332688 441888 333008 441922
rect 363408 442350 363728 442384
rect 363408 442294 363478 442350
rect 363534 442294 363602 442350
rect 363658 442294 363728 442350
rect 363408 442226 363728 442294
rect 363408 442170 363478 442226
rect 363534 442170 363602 442226
rect 363658 442170 363728 442226
rect 363408 442102 363728 442170
rect 363408 442046 363478 442102
rect 363534 442046 363602 442102
rect 363658 442046 363728 442102
rect 363408 441978 363728 442046
rect 363408 441922 363478 441978
rect 363534 441922 363602 441978
rect 363658 441922 363728 441978
rect 363408 441888 363728 441922
rect 394128 442350 394448 442384
rect 394128 442294 394198 442350
rect 394254 442294 394322 442350
rect 394378 442294 394448 442350
rect 394128 442226 394448 442294
rect 394128 442170 394198 442226
rect 394254 442170 394322 442226
rect 394378 442170 394448 442226
rect 394128 442102 394448 442170
rect 394128 442046 394198 442102
rect 394254 442046 394322 442102
rect 394378 442046 394448 442102
rect 394128 441978 394448 442046
rect 394128 441922 394198 441978
rect 394254 441922 394322 441978
rect 394378 441922 394448 441978
rect 394128 441888 394448 441922
rect 424848 442350 425168 442384
rect 424848 442294 424918 442350
rect 424974 442294 425042 442350
rect 425098 442294 425168 442350
rect 424848 442226 425168 442294
rect 424848 442170 424918 442226
rect 424974 442170 425042 442226
rect 425098 442170 425168 442226
rect 424848 442102 425168 442170
rect 424848 442046 424918 442102
rect 424974 442046 425042 442102
rect 425098 442046 425168 442102
rect 424848 441978 425168 442046
rect 424848 441922 424918 441978
rect 424974 441922 425042 441978
rect 425098 441922 425168 441978
rect 424848 441888 425168 441922
rect 225168 436350 225488 436384
rect 225168 436294 225238 436350
rect 225294 436294 225362 436350
rect 225418 436294 225488 436350
rect 225168 436226 225488 436294
rect 225168 436170 225238 436226
rect 225294 436170 225362 436226
rect 225418 436170 225488 436226
rect 225168 436102 225488 436170
rect 225168 436046 225238 436102
rect 225294 436046 225362 436102
rect 225418 436046 225488 436102
rect 225168 435978 225488 436046
rect 225168 435922 225238 435978
rect 225294 435922 225362 435978
rect 225418 435922 225488 435978
rect 225168 435888 225488 435922
rect 255888 436350 256208 436384
rect 255888 436294 255958 436350
rect 256014 436294 256082 436350
rect 256138 436294 256208 436350
rect 255888 436226 256208 436294
rect 255888 436170 255958 436226
rect 256014 436170 256082 436226
rect 256138 436170 256208 436226
rect 255888 436102 256208 436170
rect 255888 436046 255958 436102
rect 256014 436046 256082 436102
rect 256138 436046 256208 436102
rect 255888 435978 256208 436046
rect 255888 435922 255958 435978
rect 256014 435922 256082 435978
rect 256138 435922 256208 435978
rect 255888 435888 256208 435922
rect 286608 436350 286928 436384
rect 286608 436294 286678 436350
rect 286734 436294 286802 436350
rect 286858 436294 286928 436350
rect 286608 436226 286928 436294
rect 286608 436170 286678 436226
rect 286734 436170 286802 436226
rect 286858 436170 286928 436226
rect 286608 436102 286928 436170
rect 286608 436046 286678 436102
rect 286734 436046 286802 436102
rect 286858 436046 286928 436102
rect 286608 435978 286928 436046
rect 286608 435922 286678 435978
rect 286734 435922 286802 435978
rect 286858 435922 286928 435978
rect 286608 435888 286928 435922
rect 317328 436350 317648 436384
rect 317328 436294 317398 436350
rect 317454 436294 317522 436350
rect 317578 436294 317648 436350
rect 317328 436226 317648 436294
rect 317328 436170 317398 436226
rect 317454 436170 317522 436226
rect 317578 436170 317648 436226
rect 317328 436102 317648 436170
rect 317328 436046 317398 436102
rect 317454 436046 317522 436102
rect 317578 436046 317648 436102
rect 317328 435978 317648 436046
rect 317328 435922 317398 435978
rect 317454 435922 317522 435978
rect 317578 435922 317648 435978
rect 317328 435888 317648 435922
rect 348048 436350 348368 436384
rect 348048 436294 348118 436350
rect 348174 436294 348242 436350
rect 348298 436294 348368 436350
rect 348048 436226 348368 436294
rect 348048 436170 348118 436226
rect 348174 436170 348242 436226
rect 348298 436170 348368 436226
rect 348048 436102 348368 436170
rect 348048 436046 348118 436102
rect 348174 436046 348242 436102
rect 348298 436046 348368 436102
rect 348048 435978 348368 436046
rect 348048 435922 348118 435978
rect 348174 435922 348242 435978
rect 348298 435922 348368 435978
rect 348048 435888 348368 435922
rect 378768 436350 379088 436384
rect 378768 436294 378838 436350
rect 378894 436294 378962 436350
rect 379018 436294 379088 436350
rect 378768 436226 379088 436294
rect 378768 436170 378838 436226
rect 378894 436170 378962 436226
rect 379018 436170 379088 436226
rect 378768 436102 379088 436170
rect 378768 436046 378838 436102
rect 378894 436046 378962 436102
rect 379018 436046 379088 436102
rect 378768 435978 379088 436046
rect 378768 435922 378838 435978
rect 378894 435922 378962 435978
rect 379018 435922 379088 435978
rect 378768 435888 379088 435922
rect 409488 436350 409808 436384
rect 409488 436294 409558 436350
rect 409614 436294 409682 436350
rect 409738 436294 409808 436350
rect 409488 436226 409808 436294
rect 409488 436170 409558 436226
rect 409614 436170 409682 436226
rect 409738 436170 409808 436226
rect 409488 436102 409808 436170
rect 409488 436046 409558 436102
rect 409614 436046 409682 436102
rect 409738 436046 409808 436102
rect 409488 435978 409808 436046
rect 409488 435922 409558 435978
rect 409614 435922 409682 435978
rect 409738 435922 409808 435978
rect 409488 435888 409808 435922
rect 440208 436350 440528 436384
rect 440208 436294 440278 436350
rect 440334 436294 440402 436350
rect 440458 436294 440528 436350
rect 440208 436226 440528 436294
rect 440208 436170 440278 436226
rect 440334 436170 440402 436226
rect 440458 436170 440528 436226
rect 440208 436102 440528 436170
rect 440208 436046 440278 436102
rect 440334 436046 440402 436102
rect 440458 436046 440528 436102
rect 440208 435978 440528 436046
rect 440208 435922 440278 435978
rect 440334 435922 440402 435978
rect 440458 435922 440528 435978
rect 440208 435888 440528 435922
rect 209808 424350 210128 424384
rect 209808 424294 209878 424350
rect 209934 424294 210002 424350
rect 210058 424294 210128 424350
rect 209808 424226 210128 424294
rect 209808 424170 209878 424226
rect 209934 424170 210002 424226
rect 210058 424170 210128 424226
rect 209808 424102 210128 424170
rect 209808 424046 209878 424102
rect 209934 424046 210002 424102
rect 210058 424046 210128 424102
rect 209808 423978 210128 424046
rect 209808 423922 209878 423978
rect 209934 423922 210002 423978
rect 210058 423922 210128 423978
rect 209808 423888 210128 423922
rect 240528 424350 240848 424384
rect 240528 424294 240598 424350
rect 240654 424294 240722 424350
rect 240778 424294 240848 424350
rect 240528 424226 240848 424294
rect 240528 424170 240598 424226
rect 240654 424170 240722 424226
rect 240778 424170 240848 424226
rect 240528 424102 240848 424170
rect 240528 424046 240598 424102
rect 240654 424046 240722 424102
rect 240778 424046 240848 424102
rect 240528 423978 240848 424046
rect 240528 423922 240598 423978
rect 240654 423922 240722 423978
rect 240778 423922 240848 423978
rect 240528 423888 240848 423922
rect 271248 424350 271568 424384
rect 271248 424294 271318 424350
rect 271374 424294 271442 424350
rect 271498 424294 271568 424350
rect 271248 424226 271568 424294
rect 271248 424170 271318 424226
rect 271374 424170 271442 424226
rect 271498 424170 271568 424226
rect 271248 424102 271568 424170
rect 271248 424046 271318 424102
rect 271374 424046 271442 424102
rect 271498 424046 271568 424102
rect 271248 423978 271568 424046
rect 271248 423922 271318 423978
rect 271374 423922 271442 423978
rect 271498 423922 271568 423978
rect 271248 423888 271568 423922
rect 301968 424350 302288 424384
rect 301968 424294 302038 424350
rect 302094 424294 302162 424350
rect 302218 424294 302288 424350
rect 301968 424226 302288 424294
rect 301968 424170 302038 424226
rect 302094 424170 302162 424226
rect 302218 424170 302288 424226
rect 301968 424102 302288 424170
rect 301968 424046 302038 424102
rect 302094 424046 302162 424102
rect 302218 424046 302288 424102
rect 301968 423978 302288 424046
rect 301968 423922 302038 423978
rect 302094 423922 302162 423978
rect 302218 423922 302288 423978
rect 301968 423888 302288 423922
rect 332688 424350 333008 424384
rect 332688 424294 332758 424350
rect 332814 424294 332882 424350
rect 332938 424294 333008 424350
rect 332688 424226 333008 424294
rect 332688 424170 332758 424226
rect 332814 424170 332882 424226
rect 332938 424170 333008 424226
rect 332688 424102 333008 424170
rect 332688 424046 332758 424102
rect 332814 424046 332882 424102
rect 332938 424046 333008 424102
rect 332688 423978 333008 424046
rect 332688 423922 332758 423978
rect 332814 423922 332882 423978
rect 332938 423922 333008 423978
rect 332688 423888 333008 423922
rect 363408 424350 363728 424384
rect 363408 424294 363478 424350
rect 363534 424294 363602 424350
rect 363658 424294 363728 424350
rect 363408 424226 363728 424294
rect 363408 424170 363478 424226
rect 363534 424170 363602 424226
rect 363658 424170 363728 424226
rect 363408 424102 363728 424170
rect 363408 424046 363478 424102
rect 363534 424046 363602 424102
rect 363658 424046 363728 424102
rect 363408 423978 363728 424046
rect 363408 423922 363478 423978
rect 363534 423922 363602 423978
rect 363658 423922 363728 423978
rect 363408 423888 363728 423922
rect 394128 424350 394448 424384
rect 394128 424294 394198 424350
rect 394254 424294 394322 424350
rect 394378 424294 394448 424350
rect 394128 424226 394448 424294
rect 394128 424170 394198 424226
rect 394254 424170 394322 424226
rect 394378 424170 394448 424226
rect 394128 424102 394448 424170
rect 394128 424046 394198 424102
rect 394254 424046 394322 424102
rect 394378 424046 394448 424102
rect 394128 423978 394448 424046
rect 394128 423922 394198 423978
rect 394254 423922 394322 423978
rect 394378 423922 394448 423978
rect 394128 423888 394448 423922
rect 424848 424350 425168 424384
rect 424848 424294 424918 424350
rect 424974 424294 425042 424350
rect 425098 424294 425168 424350
rect 424848 424226 425168 424294
rect 424848 424170 424918 424226
rect 424974 424170 425042 424226
rect 425098 424170 425168 424226
rect 424848 424102 425168 424170
rect 424848 424046 424918 424102
rect 424974 424046 425042 424102
rect 425098 424046 425168 424102
rect 424848 423978 425168 424046
rect 424848 423922 424918 423978
rect 424974 423922 425042 423978
rect 425098 423922 425168 423978
rect 424848 423888 425168 423922
rect 225168 418350 225488 418384
rect 225168 418294 225238 418350
rect 225294 418294 225362 418350
rect 225418 418294 225488 418350
rect 225168 418226 225488 418294
rect 225168 418170 225238 418226
rect 225294 418170 225362 418226
rect 225418 418170 225488 418226
rect 225168 418102 225488 418170
rect 225168 418046 225238 418102
rect 225294 418046 225362 418102
rect 225418 418046 225488 418102
rect 225168 417978 225488 418046
rect 225168 417922 225238 417978
rect 225294 417922 225362 417978
rect 225418 417922 225488 417978
rect 225168 417888 225488 417922
rect 255888 418350 256208 418384
rect 255888 418294 255958 418350
rect 256014 418294 256082 418350
rect 256138 418294 256208 418350
rect 255888 418226 256208 418294
rect 255888 418170 255958 418226
rect 256014 418170 256082 418226
rect 256138 418170 256208 418226
rect 255888 418102 256208 418170
rect 255888 418046 255958 418102
rect 256014 418046 256082 418102
rect 256138 418046 256208 418102
rect 255888 417978 256208 418046
rect 255888 417922 255958 417978
rect 256014 417922 256082 417978
rect 256138 417922 256208 417978
rect 255888 417888 256208 417922
rect 286608 418350 286928 418384
rect 286608 418294 286678 418350
rect 286734 418294 286802 418350
rect 286858 418294 286928 418350
rect 286608 418226 286928 418294
rect 286608 418170 286678 418226
rect 286734 418170 286802 418226
rect 286858 418170 286928 418226
rect 286608 418102 286928 418170
rect 286608 418046 286678 418102
rect 286734 418046 286802 418102
rect 286858 418046 286928 418102
rect 286608 417978 286928 418046
rect 286608 417922 286678 417978
rect 286734 417922 286802 417978
rect 286858 417922 286928 417978
rect 286608 417888 286928 417922
rect 317328 418350 317648 418384
rect 317328 418294 317398 418350
rect 317454 418294 317522 418350
rect 317578 418294 317648 418350
rect 317328 418226 317648 418294
rect 317328 418170 317398 418226
rect 317454 418170 317522 418226
rect 317578 418170 317648 418226
rect 317328 418102 317648 418170
rect 317328 418046 317398 418102
rect 317454 418046 317522 418102
rect 317578 418046 317648 418102
rect 317328 417978 317648 418046
rect 317328 417922 317398 417978
rect 317454 417922 317522 417978
rect 317578 417922 317648 417978
rect 317328 417888 317648 417922
rect 348048 418350 348368 418384
rect 348048 418294 348118 418350
rect 348174 418294 348242 418350
rect 348298 418294 348368 418350
rect 348048 418226 348368 418294
rect 348048 418170 348118 418226
rect 348174 418170 348242 418226
rect 348298 418170 348368 418226
rect 348048 418102 348368 418170
rect 348048 418046 348118 418102
rect 348174 418046 348242 418102
rect 348298 418046 348368 418102
rect 348048 417978 348368 418046
rect 348048 417922 348118 417978
rect 348174 417922 348242 417978
rect 348298 417922 348368 417978
rect 348048 417888 348368 417922
rect 378768 418350 379088 418384
rect 378768 418294 378838 418350
rect 378894 418294 378962 418350
rect 379018 418294 379088 418350
rect 378768 418226 379088 418294
rect 378768 418170 378838 418226
rect 378894 418170 378962 418226
rect 379018 418170 379088 418226
rect 378768 418102 379088 418170
rect 378768 418046 378838 418102
rect 378894 418046 378962 418102
rect 379018 418046 379088 418102
rect 378768 417978 379088 418046
rect 378768 417922 378838 417978
rect 378894 417922 378962 417978
rect 379018 417922 379088 417978
rect 378768 417888 379088 417922
rect 409488 418350 409808 418384
rect 409488 418294 409558 418350
rect 409614 418294 409682 418350
rect 409738 418294 409808 418350
rect 409488 418226 409808 418294
rect 409488 418170 409558 418226
rect 409614 418170 409682 418226
rect 409738 418170 409808 418226
rect 409488 418102 409808 418170
rect 409488 418046 409558 418102
rect 409614 418046 409682 418102
rect 409738 418046 409808 418102
rect 409488 417978 409808 418046
rect 409488 417922 409558 417978
rect 409614 417922 409682 417978
rect 409738 417922 409808 417978
rect 409488 417888 409808 417922
rect 440208 418350 440528 418384
rect 440208 418294 440278 418350
rect 440334 418294 440402 418350
rect 440458 418294 440528 418350
rect 440208 418226 440528 418294
rect 440208 418170 440278 418226
rect 440334 418170 440402 418226
rect 440458 418170 440528 418226
rect 440208 418102 440528 418170
rect 440208 418046 440278 418102
rect 440334 418046 440402 418102
rect 440458 418046 440528 418102
rect 440208 417978 440528 418046
rect 440208 417922 440278 417978
rect 440334 417922 440402 417978
rect 440458 417922 440528 417978
rect 440208 417888 440528 417922
rect 355404 410116 355460 410126
rect 354396 409798 354452 409808
rect 289772 409438 289828 409448
rect 288876 409258 288932 409268
rect 209468 407810 209524 407820
rect 209916 404398 209972 404408
rect 208236 399074 208292 399084
rect 209804 402778 209860 402788
rect 208124 382386 208180 382396
rect 209804 382452 209860 402722
rect 209916 382564 209972 404342
rect 209916 382498 209972 382508
rect 220458 400350 221078 408466
rect 220458 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 221078 400350
rect 220458 400226 221078 400294
rect 220458 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 221078 400226
rect 220458 400102 221078 400170
rect 220458 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 221078 400102
rect 220458 399978 221078 400046
rect 220458 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 221078 399978
rect 209804 382386 209860 382396
rect 220458 382350 221078 399922
rect 220458 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 221078 382350
rect 220458 382226 221078 382294
rect 220458 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 221078 382226
rect 220458 382102 221078 382170
rect 220458 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 221078 382102
rect 220458 381978 221078 382046
rect 220458 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 221078 381978
rect 214172 379652 214228 379662
rect 214172 379204 214228 379596
rect 214172 379138 214228 379148
rect 214396 379652 214452 379662
rect 214396 379092 214452 379596
rect 214396 379026 214452 379036
rect 209808 370350 210128 370384
rect 209808 370294 209878 370350
rect 209934 370294 210002 370350
rect 210058 370294 210128 370350
rect 209808 370226 210128 370294
rect 209808 370170 209878 370226
rect 209934 370170 210002 370226
rect 210058 370170 210128 370226
rect 209808 370102 210128 370170
rect 209808 370046 209878 370102
rect 209934 370046 210002 370102
rect 210058 370046 210128 370102
rect 209808 369978 210128 370046
rect 209808 369922 209878 369978
rect 209934 369922 210002 369978
rect 210058 369922 210128 369978
rect 209808 369888 210128 369922
rect 210812 368038 210868 368048
rect 209808 352350 210128 352384
rect 209808 352294 209878 352350
rect 209934 352294 210002 352350
rect 210058 352294 210128 352350
rect 209808 352226 210128 352294
rect 209808 352170 209878 352226
rect 209934 352170 210002 352226
rect 210058 352170 210128 352226
rect 209808 352102 210128 352170
rect 209808 352046 209878 352102
rect 209934 352046 210002 352102
rect 210058 352046 210128 352102
rect 209808 351978 210128 352046
rect 209808 351922 209878 351978
rect 209934 351922 210002 351978
rect 210058 351922 210128 351978
rect 209808 351888 210128 351922
rect 206668 340072 206724 340082
rect 209808 334350 210128 334384
rect 209808 334294 209878 334350
rect 209934 334294 210002 334350
rect 210058 334294 210128 334350
rect 209808 334226 210128 334294
rect 209808 334170 209878 334226
rect 209934 334170 210002 334226
rect 210058 334170 210128 334226
rect 209808 334102 210128 334170
rect 209808 334046 209878 334102
rect 209934 334046 210002 334102
rect 210058 334046 210128 334102
rect 209808 333978 210128 334046
rect 209808 333922 209878 333978
rect 209934 333922 210002 333978
rect 210058 333922 210128 333978
rect 209808 333888 210128 333922
rect 209808 316350 210128 316384
rect 209808 316294 209878 316350
rect 209934 316294 210002 316350
rect 210058 316294 210128 316350
rect 209808 316226 210128 316294
rect 209808 316170 209878 316226
rect 209934 316170 210002 316226
rect 210058 316170 210128 316226
rect 209808 316102 210128 316170
rect 209808 316046 209878 316102
rect 209934 316046 210002 316102
rect 210058 316046 210128 316102
rect 209808 315978 210128 316046
rect 209808 315922 209878 315978
rect 209934 315922 210002 315978
rect 210058 315922 210128 315978
rect 209808 315888 210128 315922
rect 209808 298350 210128 298384
rect 209808 298294 209878 298350
rect 209934 298294 210002 298350
rect 210058 298294 210128 298350
rect 209808 298226 210128 298294
rect 209808 298170 209878 298226
rect 209934 298170 210002 298226
rect 210058 298170 210128 298226
rect 209808 298102 210128 298170
rect 209808 298046 209878 298102
rect 209934 298046 210002 298102
rect 210058 298046 210128 298102
rect 209808 297978 210128 298046
rect 209808 297922 209878 297978
rect 209934 297922 210002 297978
rect 210058 297922 210128 297978
rect 209808 297888 210128 297922
rect 209808 280350 210128 280384
rect 209808 280294 209878 280350
rect 209934 280294 210002 280350
rect 210058 280294 210128 280350
rect 209808 280226 210128 280294
rect 209808 280170 209878 280226
rect 209934 280170 210002 280226
rect 210058 280170 210128 280226
rect 209808 280102 210128 280170
rect 209808 280046 209878 280102
rect 209934 280046 210002 280102
rect 210058 280046 210128 280102
rect 209808 279978 210128 280046
rect 209808 279922 209878 279978
rect 209934 279922 210002 279978
rect 210058 279922 210128 279978
rect 209808 279888 210128 279922
rect 209808 262350 210128 262384
rect 209808 262294 209878 262350
rect 209934 262294 210002 262350
rect 210058 262294 210128 262350
rect 209808 262226 210128 262294
rect 209808 262170 209878 262226
rect 209934 262170 210002 262226
rect 210058 262170 210128 262226
rect 209808 262102 210128 262170
rect 209808 262046 209878 262102
rect 209934 262046 210002 262102
rect 210058 262046 210128 262102
rect 209808 261978 210128 262046
rect 209808 261922 209878 261978
rect 209934 261922 210002 261978
rect 210058 261922 210128 261978
rect 209808 261888 210128 261922
rect 209808 244350 210128 244384
rect 209808 244294 209878 244350
rect 209934 244294 210002 244350
rect 210058 244294 210128 244350
rect 209808 244226 210128 244294
rect 209808 244170 209878 244226
rect 209934 244170 210002 244226
rect 210058 244170 210128 244226
rect 209808 244102 210128 244170
rect 209808 244046 209878 244102
rect 209934 244046 210002 244102
rect 210058 244046 210128 244102
rect 209808 243978 210128 244046
rect 209808 243922 209878 243978
rect 209934 243922 210002 243978
rect 210058 243922 210128 243978
rect 209808 243888 210128 243922
rect 209916 236964 209972 236974
rect 209916 231058 209972 236908
rect 209916 230992 209972 231002
rect 210812 216244 210868 367982
rect 214172 366598 214228 366608
rect 214172 216356 214228 366542
rect 217532 366418 217588 366428
rect 214284 364618 214340 364628
rect 214284 219828 214340 364562
rect 214284 219762 214340 219772
rect 214172 216290 214228 216300
rect 210812 216178 210868 216188
rect 203196 214610 203252 214620
rect 217532 213220 217588 366362
rect 220458 364350 221078 381922
rect 224178 406350 224798 408466
rect 224178 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 224798 406350
rect 224178 406226 224798 406294
rect 224178 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 224798 406226
rect 224178 406102 224798 406170
rect 224178 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 224798 406102
rect 224178 405978 224798 406046
rect 224178 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 224798 405978
rect 224178 388350 224798 405922
rect 229964 406644 230020 406654
rect 224178 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 224798 388350
rect 224178 388226 224798 388294
rect 224178 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 224798 388226
rect 224178 388102 224798 388170
rect 224178 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 224798 388102
rect 224178 387978 224798 388046
rect 224178 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 224798 387978
rect 222012 379540 222068 379550
rect 222012 372178 222068 379484
rect 224028 379540 224084 379550
rect 224028 378838 224084 379484
rect 224028 378772 224084 378782
rect 222012 372112 222068 372122
rect 220458 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 221078 364350
rect 220458 364226 221078 364294
rect 220458 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 221078 364226
rect 220458 364102 221078 364170
rect 220458 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 221078 364102
rect 220458 363978 221078 364046
rect 220458 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 221078 363978
rect 220458 346350 221078 363922
rect 220458 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 221078 346350
rect 220458 346226 221078 346294
rect 220458 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 221078 346226
rect 220458 346102 221078 346170
rect 220458 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 221078 346102
rect 220458 345978 221078 346046
rect 220458 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 221078 345978
rect 220458 328350 221078 345922
rect 220458 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 221078 328350
rect 220458 328226 221078 328294
rect 220458 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 221078 328226
rect 220458 328102 221078 328170
rect 220458 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 221078 328102
rect 220458 327978 221078 328046
rect 220458 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 221078 327978
rect 217644 319258 217700 319268
rect 217644 222740 217700 319202
rect 217644 222674 217700 222684
rect 220458 310350 221078 327922
rect 220458 310294 220554 310350
rect 220610 310294 220678 310350
rect 220734 310294 220802 310350
rect 220858 310294 220926 310350
rect 220982 310294 221078 310350
rect 220458 310226 221078 310294
rect 220458 310170 220554 310226
rect 220610 310170 220678 310226
rect 220734 310170 220802 310226
rect 220858 310170 220926 310226
rect 220982 310170 221078 310226
rect 220458 310102 221078 310170
rect 220458 310046 220554 310102
rect 220610 310046 220678 310102
rect 220734 310046 220802 310102
rect 220858 310046 220926 310102
rect 220982 310046 221078 310102
rect 220458 309978 221078 310046
rect 220458 309922 220554 309978
rect 220610 309922 220678 309978
rect 220734 309922 220802 309978
rect 220858 309922 220926 309978
rect 220982 309922 221078 309978
rect 220458 292350 221078 309922
rect 220458 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 221078 292350
rect 220458 292226 221078 292294
rect 220458 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 221078 292226
rect 220458 292102 221078 292170
rect 220458 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 221078 292102
rect 220458 291978 221078 292046
rect 220458 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 221078 291978
rect 220458 274350 221078 291922
rect 220458 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 221078 274350
rect 220458 274226 221078 274294
rect 220458 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 221078 274226
rect 220458 274102 221078 274170
rect 220458 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 221078 274102
rect 220458 273978 221078 274046
rect 220458 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 221078 273978
rect 220458 256350 221078 273922
rect 220458 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 221078 256350
rect 220458 256226 221078 256294
rect 220458 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 221078 256226
rect 220458 256102 221078 256170
rect 220458 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 221078 256102
rect 220458 255978 221078 256046
rect 220458 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 221078 255978
rect 220458 238350 221078 255922
rect 220458 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 221078 238350
rect 220458 238226 221078 238294
rect 220458 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 221078 238226
rect 220458 238102 221078 238170
rect 220458 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 221078 238102
rect 220458 237978 221078 238046
rect 220458 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 221078 237978
rect 217532 213154 217588 213164
rect 220458 220350 221078 237922
rect 220458 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 221078 220350
rect 220458 220226 221078 220294
rect 220458 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 221078 220226
rect 220458 220102 221078 220170
rect 220458 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 221078 220102
rect 220458 219978 221078 220046
rect 220458 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 221078 219978
rect 201404 213042 201460 213052
rect 220458 210574 221078 219922
rect 224178 370350 224798 387922
rect 226716 394858 226772 394868
rect 226716 382116 226772 394802
rect 226716 382050 226772 382060
rect 227612 379540 227668 379550
rect 225148 379316 225204 379326
rect 225148 377398 225204 379260
rect 225148 377332 225204 377342
rect 225820 379316 225876 379326
rect 225820 377218 225876 379260
rect 225820 377152 225876 377162
rect 224178 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 224798 370350
rect 224178 370226 224798 370294
rect 224178 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 224798 370226
rect 224178 370102 224798 370170
rect 224178 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 224798 370102
rect 224178 369978 224798 370046
rect 224178 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 224798 369978
rect 224178 352350 224798 369922
rect 225168 364350 225488 364384
rect 225168 364294 225238 364350
rect 225294 364294 225362 364350
rect 225418 364294 225488 364350
rect 225168 364226 225488 364294
rect 225168 364170 225238 364226
rect 225294 364170 225362 364226
rect 225418 364170 225488 364226
rect 225168 364102 225488 364170
rect 225168 364046 225238 364102
rect 225294 364046 225362 364102
rect 225418 364046 225488 364102
rect 225168 363978 225488 364046
rect 225168 363922 225238 363978
rect 225294 363922 225362 363978
rect 225418 363922 225488 363978
rect 225168 363888 225488 363922
rect 224178 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 224798 352350
rect 224178 352226 224798 352294
rect 224178 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 224798 352226
rect 224178 352102 224798 352170
rect 224178 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 224798 352102
rect 224178 351978 224798 352046
rect 224178 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 224798 351978
rect 224178 334350 224798 351922
rect 225168 346350 225488 346384
rect 225168 346294 225238 346350
rect 225294 346294 225362 346350
rect 225418 346294 225488 346350
rect 225168 346226 225488 346294
rect 225168 346170 225238 346226
rect 225294 346170 225362 346226
rect 225418 346170 225488 346226
rect 225168 346102 225488 346170
rect 225168 346046 225238 346102
rect 225294 346046 225362 346102
rect 225418 346046 225488 346102
rect 225168 345978 225488 346046
rect 225168 345922 225238 345978
rect 225294 345922 225362 345978
rect 225418 345922 225488 345978
rect 225168 345888 225488 345922
rect 224178 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 224798 334350
rect 224178 334226 224798 334294
rect 224178 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 224798 334226
rect 224178 334102 224798 334170
rect 224178 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 224798 334102
rect 224178 333978 224798 334046
rect 224178 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 224798 333978
rect 224178 316350 224798 333922
rect 225168 328350 225488 328384
rect 225168 328294 225238 328350
rect 225294 328294 225362 328350
rect 225418 328294 225488 328350
rect 225168 328226 225488 328294
rect 225168 328170 225238 328226
rect 225294 328170 225362 328226
rect 225418 328170 225488 328226
rect 225168 328102 225488 328170
rect 225168 328046 225238 328102
rect 225294 328046 225362 328102
rect 225418 328046 225488 328102
rect 225168 327978 225488 328046
rect 225168 327922 225238 327978
rect 225294 327922 225362 327978
rect 225418 327922 225488 327978
rect 225168 327888 225488 327922
rect 224178 316294 224274 316350
rect 224330 316294 224398 316350
rect 224454 316294 224522 316350
rect 224578 316294 224646 316350
rect 224702 316294 224798 316350
rect 224178 316226 224798 316294
rect 224178 316170 224274 316226
rect 224330 316170 224398 316226
rect 224454 316170 224522 316226
rect 224578 316170 224646 316226
rect 224702 316170 224798 316226
rect 224178 316102 224798 316170
rect 224178 316046 224274 316102
rect 224330 316046 224398 316102
rect 224454 316046 224522 316102
rect 224578 316046 224646 316102
rect 224702 316046 224798 316102
rect 224178 315978 224798 316046
rect 224178 315922 224274 315978
rect 224330 315922 224398 315978
rect 224454 315922 224522 315978
rect 224578 315922 224646 315978
rect 224702 315922 224798 315978
rect 224178 298350 224798 315922
rect 225168 310350 225488 310384
rect 225168 310294 225238 310350
rect 225294 310294 225362 310350
rect 225418 310294 225488 310350
rect 225168 310226 225488 310294
rect 225168 310170 225238 310226
rect 225294 310170 225362 310226
rect 225418 310170 225488 310226
rect 225168 310102 225488 310170
rect 225168 310046 225238 310102
rect 225294 310046 225362 310102
rect 225418 310046 225488 310102
rect 225168 309978 225488 310046
rect 225168 309922 225238 309978
rect 225294 309922 225362 309978
rect 225418 309922 225488 309978
rect 225168 309888 225488 309922
rect 224178 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 224798 298350
rect 224178 298226 224798 298294
rect 224178 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 224798 298226
rect 224178 298102 224798 298170
rect 224178 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 224798 298102
rect 224178 297978 224798 298046
rect 224178 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 224798 297978
rect 224178 280350 224798 297922
rect 225168 292350 225488 292384
rect 225168 292294 225238 292350
rect 225294 292294 225362 292350
rect 225418 292294 225488 292350
rect 225168 292226 225488 292294
rect 225168 292170 225238 292226
rect 225294 292170 225362 292226
rect 225418 292170 225488 292226
rect 225168 292102 225488 292170
rect 225168 292046 225238 292102
rect 225294 292046 225362 292102
rect 225418 292046 225488 292102
rect 225168 291978 225488 292046
rect 225168 291922 225238 291978
rect 225294 291922 225362 291978
rect 225418 291922 225488 291978
rect 225168 291888 225488 291922
rect 224178 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 224798 280350
rect 224178 280226 224798 280294
rect 224178 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 224798 280226
rect 224178 280102 224798 280170
rect 224178 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 224798 280102
rect 224178 279978 224798 280046
rect 224178 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 224798 279978
rect 224178 262350 224798 279922
rect 225168 274350 225488 274384
rect 225168 274294 225238 274350
rect 225294 274294 225362 274350
rect 225418 274294 225488 274350
rect 225168 274226 225488 274294
rect 225168 274170 225238 274226
rect 225294 274170 225362 274226
rect 225418 274170 225488 274226
rect 225168 274102 225488 274170
rect 225168 274046 225238 274102
rect 225294 274046 225362 274102
rect 225418 274046 225488 274102
rect 225168 273978 225488 274046
rect 225168 273922 225238 273978
rect 225294 273922 225362 273978
rect 225418 273922 225488 273978
rect 225168 273888 225488 273922
rect 224178 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 224798 262350
rect 224178 262226 224798 262294
rect 224178 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 224798 262226
rect 224178 262102 224798 262170
rect 224178 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 224798 262102
rect 224178 261978 224798 262046
rect 224178 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 224798 261978
rect 224178 244350 224798 261922
rect 225168 256350 225488 256384
rect 225168 256294 225238 256350
rect 225294 256294 225362 256350
rect 225418 256294 225488 256350
rect 225168 256226 225488 256294
rect 225168 256170 225238 256226
rect 225294 256170 225362 256226
rect 225418 256170 225488 256226
rect 225168 256102 225488 256170
rect 225168 256046 225238 256102
rect 225294 256046 225362 256102
rect 225418 256046 225488 256102
rect 225168 255978 225488 256046
rect 225168 255922 225238 255978
rect 225294 255922 225362 255978
rect 225418 255922 225488 255978
rect 225168 255888 225488 255922
rect 224178 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 224798 244350
rect 224178 244226 224798 244294
rect 224178 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 224798 244226
rect 224178 244102 224798 244170
rect 224178 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 224798 244102
rect 224178 243978 224798 244046
rect 224178 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 224798 243978
rect 224178 226350 224798 243922
rect 224178 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 224798 226350
rect 224178 226226 224798 226294
rect 224178 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 224798 226226
rect 224178 226102 224798 226170
rect 224178 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 224798 226102
rect 224178 225978 224798 226046
rect 224178 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 224798 225978
rect 224178 210574 224798 225922
rect 225148 236964 225204 236974
rect 225148 224218 225204 236908
rect 225148 224152 225204 224162
rect 227612 212660 227668 379484
rect 227836 379316 227892 379326
rect 227836 372988 227892 379260
rect 227836 372932 228228 372988
rect 228172 214228 228228 372932
rect 229964 272098 230020 406588
rect 251178 400350 251798 408466
rect 251178 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 251798 400350
rect 251178 400226 251798 400294
rect 251178 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 251798 400226
rect 251178 400102 251798 400170
rect 251178 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 251798 400102
rect 251178 399978 251798 400046
rect 251178 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 251798 399978
rect 239484 398458 239540 398468
rect 239372 392698 239428 392708
rect 235116 386036 235172 386046
rect 232764 381444 232820 381454
rect 229964 272032 230020 272042
rect 230076 379540 230132 379550
rect 228172 214162 228228 214172
rect 230076 212772 230132 379484
rect 232540 379316 232596 379326
rect 232540 373798 232596 379260
rect 232540 373732 232596 373742
rect 230972 272098 231028 272108
rect 230972 265438 231028 272042
rect 230972 239428 231028 265382
rect 232764 240548 232820 381388
rect 235116 293878 235172 385980
rect 238364 384916 238420 384926
rect 237804 383124 237860 383134
rect 237692 380772 237748 380782
rect 235452 379540 235508 379550
rect 235452 361228 235508 379484
rect 235116 293812 235172 293822
rect 235228 361172 235508 361228
rect 232764 240482 232820 240492
rect 230972 239362 231028 239372
rect 233436 236964 233492 236974
rect 233436 224218 233492 236908
rect 235228 233492 235284 361172
rect 237692 302428 237748 380716
rect 237804 311698 237860 383068
rect 237804 311632 237860 311642
rect 236908 302372 237748 302428
rect 236908 295678 236964 302372
rect 236796 295622 236964 295678
rect 236796 294058 236852 295622
rect 238364 294778 238420 384860
rect 238364 294712 238420 294722
rect 238476 384468 238532 384478
rect 236012 287398 236068 287408
rect 236012 236404 236068 287342
rect 236236 285958 236292 285968
rect 236124 283978 236180 283988
rect 236124 240548 236180 283922
rect 236124 240482 236180 240492
rect 236012 236338 236068 236348
rect 236236 236292 236292 285902
rect 236348 270658 236404 270668
rect 236348 241678 236404 270602
rect 236348 241612 236404 241622
rect 236796 239316 236852 294002
rect 238476 239876 238532 384412
rect 238588 384356 238644 384366
rect 238588 376318 238644 384300
rect 238588 376252 238644 376262
rect 239372 260398 239428 392642
rect 239484 288838 239540 398402
rect 250236 392338 250292 392348
rect 241836 384580 241892 384590
rect 241500 381444 241556 381454
rect 240156 380884 240212 380894
rect 239708 294778 239764 294788
rect 239484 288772 239540 288782
rect 239596 292618 239652 292628
rect 239372 260332 239428 260342
rect 239484 285778 239540 285788
rect 238476 239810 238532 239820
rect 239372 252118 239428 252128
rect 236796 239250 236852 239260
rect 236796 237076 236852 237086
rect 236236 236226 236292 236236
rect 236684 236964 236740 236974
rect 235228 233426 235284 233436
rect 236684 231418 236740 236908
rect 236684 231352 236740 231362
rect 236796 231238 236852 237020
rect 236796 231172 236852 231182
rect 238476 236964 238532 236974
rect 238476 227638 238532 236908
rect 238476 227572 238532 227582
rect 233436 224152 233492 224162
rect 239372 219940 239428 252062
rect 239484 236516 239540 285722
rect 239484 236450 239540 236460
rect 239372 219874 239428 219884
rect 230076 212706 230132 212716
rect 227612 212594 227668 212604
rect 239596 211438 239652 292562
rect 239708 216468 239764 294722
rect 239820 293878 239876 293888
rect 239820 234658 239876 293822
rect 239820 220108 239876 234602
rect 239932 289018 239988 289028
rect 239932 234388 239988 288962
rect 239932 234322 239988 234332
rect 240044 236964 240100 236974
rect 240044 227818 240100 236908
rect 240156 235060 240212 380828
rect 240528 370350 240848 370384
rect 240528 370294 240598 370350
rect 240654 370294 240722 370350
rect 240778 370294 240848 370350
rect 240528 370226 240848 370294
rect 240528 370170 240598 370226
rect 240654 370170 240722 370226
rect 240778 370170 240848 370226
rect 240528 370102 240848 370170
rect 240528 370046 240598 370102
rect 240654 370046 240722 370102
rect 240778 370046 240848 370102
rect 240528 369978 240848 370046
rect 240528 369922 240598 369978
rect 240654 369922 240722 369978
rect 240778 369922 240848 369978
rect 240528 369888 240848 369922
rect 240528 352350 240848 352384
rect 240528 352294 240598 352350
rect 240654 352294 240722 352350
rect 240778 352294 240848 352350
rect 240528 352226 240848 352294
rect 240528 352170 240598 352226
rect 240654 352170 240722 352226
rect 240778 352170 240848 352226
rect 240528 352102 240848 352170
rect 240528 352046 240598 352102
rect 240654 352046 240722 352102
rect 240778 352046 240848 352102
rect 240528 351978 240848 352046
rect 240528 351922 240598 351978
rect 240654 351922 240722 351978
rect 240778 351922 240848 351978
rect 240528 351888 240848 351922
rect 240528 334350 240848 334384
rect 240528 334294 240598 334350
rect 240654 334294 240722 334350
rect 240778 334294 240848 334350
rect 240528 334226 240848 334294
rect 240528 334170 240598 334226
rect 240654 334170 240722 334226
rect 240778 334170 240848 334226
rect 240528 334102 240848 334170
rect 240528 334046 240598 334102
rect 240654 334046 240722 334102
rect 240778 334046 240848 334102
rect 240528 333978 240848 334046
rect 240528 333922 240598 333978
rect 240654 333922 240722 333978
rect 240778 333922 240848 333978
rect 240528 333888 240848 333922
rect 240528 316350 240848 316384
rect 240528 316294 240598 316350
rect 240654 316294 240722 316350
rect 240778 316294 240848 316350
rect 240528 316226 240848 316294
rect 240528 316170 240598 316226
rect 240654 316170 240722 316226
rect 240778 316170 240848 316226
rect 240528 316102 240848 316170
rect 240528 316046 240598 316102
rect 240654 316046 240722 316102
rect 240778 316046 240848 316102
rect 240528 315978 240848 316046
rect 240528 315922 240598 315978
rect 240654 315922 240722 315978
rect 240778 315922 240848 315978
rect 240528 315888 240848 315922
rect 240528 298350 240848 298384
rect 240528 298294 240598 298350
rect 240654 298294 240722 298350
rect 240778 298294 240848 298350
rect 240528 298226 240848 298294
rect 240528 298170 240598 298226
rect 240654 298170 240722 298226
rect 240778 298170 240848 298226
rect 240528 298102 240848 298170
rect 240528 298046 240598 298102
rect 240654 298046 240722 298102
rect 240778 298046 240848 298102
rect 240528 297978 240848 298046
rect 240528 297922 240598 297978
rect 240654 297922 240722 297978
rect 240778 297922 240848 297978
rect 240528 297888 240848 297922
rect 240528 280350 240848 280384
rect 240528 280294 240598 280350
rect 240654 280294 240722 280350
rect 240778 280294 240848 280350
rect 240528 280226 240848 280294
rect 240528 280170 240598 280226
rect 240654 280170 240722 280226
rect 240778 280170 240848 280226
rect 240528 280102 240848 280170
rect 240528 280046 240598 280102
rect 240654 280046 240722 280102
rect 240778 280046 240848 280102
rect 240528 279978 240848 280046
rect 240528 279922 240598 279978
rect 240654 279922 240722 279978
rect 240778 279922 240848 279978
rect 240528 279888 240848 279922
rect 240528 262350 240848 262384
rect 240528 262294 240598 262350
rect 240654 262294 240722 262350
rect 240778 262294 240848 262350
rect 240528 262226 240848 262294
rect 240528 262170 240598 262226
rect 240654 262170 240722 262226
rect 240778 262170 240848 262226
rect 240528 262102 240848 262170
rect 240528 262046 240598 262102
rect 240654 262046 240722 262102
rect 240778 262046 240848 262102
rect 240528 261978 240848 262046
rect 240528 261922 240598 261978
rect 240654 261922 240722 261978
rect 240778 261922 240848 261978
rect 240528 261888 240848 261922
rect 241052 255538 241108 255548
rect 240528 244350 240848 244384
rect 240528 244294 240598 244350
rect 240654 244294 240722 244350
rect 240778 244294 240848 244350
rect 240528 244226 240848 244294
rect 240528 244170 240598 244226
rect 240654 244170 240722 244226
rect 240778 244170 240848 244226
rect 240528 244102 240848 244170
rect 240528 244046 240598 244102
rect 240654 244046 240722 244102
rect 240778 244046 240848 244102
rect 240528 243978 240848 244046
rect 240528 243922 240598 243978
rect 240654 243922 240722 243978
rect 240778 243922 240848 243978
rect 240528 243888 240848 243922
rect 240156 234994 240212 235004
rect 240044 227752 240100 227762
rect 239820 220052 240212 220108
rect 239708 216402 239764 216412
rect 239596 211372 239652 211382
rect 240156 211258 240212 220052
rect 240156 211192 240212 211202
rect 241052 211078 241108 255482
rect 241164 251218 241220 251228
rect 241164 241858 241220 251162
rect 241164 241792 241220 241802
rect 241500 235172 241556 381388
rect 241500 235106 241556 235116
rect 241724 380660 241780 380670
rect 241724 234612 241780 380604
rect 241836 239764 241892 384524
rect 250236 382004 250292 392282
rect 250236 381938 250292 381948
rect 251178 382350 251798 399922
rect 251178 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 251798 382350
rect 251178 382226 251798 382294
rect 251178 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 251798 382226
rect 251178 382102 251798 382170
rect 251178 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 251798 382102
rect 251178 381978 251798 382046
rect 251178 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 251798 381978
rect 251178 380638 251798 381922
rect 254898 406350 255518 408466
rect 254898 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 255518 406350
rect 254898 406226 255518 406294
rect 254898 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 255518 406226
rect 254898 406102 255518 406170
rect 254898 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 255518 406102
rect 254898 405978 255518 406046
rect 254898 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 255518 405978
rect 254898 388350 255518 405922
rect 280476 406644 280532 406654
rect 267036 398998 267092 399008
rect 254898 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 255518 388350
rect 254898 388226 255518 388294
rect 254898 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 255518 388226
rect 254898 388102 255518 388170
rect 254898 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 255518 388102
rect 254898 387978 255518 388046
rect 254898 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 255518 387978
rect 254898 380638 255518 387922
rect 260316 392518 260372 392528
rect 260316 382004 260372 392462
rect 260316 381938 260372 381948
rect 267036 382004 267092 398942
rect 267036 381938 267092 381948
rect 280476 380458 280532 406588
rect 281898 400350 282518 408466
rect 281898 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 282518 400350
rect 281898 400226 282518 400294
rect 281898 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 282518 400226
rect 281898 400102 282518 400170
rect 281898 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 282518 400102
rect 281898 399978 282518 400046
rect 281898 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 282518 399978
rect 281708 395578 281764 395588
rect 281708 382004 281764 395522
rect 281708 381938 281764 381948
rect 281898 382350 282518 399922
rect 281898 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 282518 382350
rect 281898 382226 282518 382294
rect 281898 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 282518 382226
rect 281898 382102 282518 382170
rect 281898 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 282518 382102
rect 281898 381978 282518 382046
rect 281898 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 282518 381978
rect 281898 380638 282518 381922
rect 285618 406350 286238 408466
rect 285618 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 286238 406350
rect 285618 406226 286238 406294
rect 285618 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 286238 406226
rect 285618 406102 286238 406170
rect 285618 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 286238 406102
rect 285618 405978 286238 406046
rect 285618 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 286238 405978
rect 285618 388350 286238 405922
rect 285618 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 286238 388350
rect 285618 388226 286238 388294
rect 285618 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 286238 388226
rect 285618 388102 286238 388170
rect 285618 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 286238 388102
rect 285618 387978 286238 388046
rect 285618 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 286238 387978
rect 285618 380638 286238 387922
rect 288092 407458 288148 407468
rect 288092 382788 288148 407402
rect 288092 382722 288148 382732
rect 288876 382004 288932 409202
rect 289772 409220 289828 409382
rect 289772 409154 289828 409164
rect 291452 409438 291508 409448
rect 288876 381938 288932 381948
rect 290556 405658 290612 405668
rect 290556 382004 290612 405602
rect 291452 382788 291508 409382
rect 295596 409078 295652 409088
rect 295596 408996 295652 409022
rect 295596 408930 295652 408940
rect 300636 408100 300692 408110
rect 299852 407998 299908 408008
rect 295596 406644 295652 406654
rect 291452 382722 291508 382732
rect 293916 390898 293972 390908
rect 290556 381938 290612 381948
rect 293916 382004 293972 390842
rect 293916 381938 293972 381948
rect 295596 380638 295652 406588
rect 299852 380818 299908 407942
rect 300636 407998 300692 408044
rect 300636 407932 300692 407942
rect 301532 405478 301588 405488
rect 301532 382116 301588 405422
rect 312618 400350 313238 408466
rect 312618 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 313238 400350
rect 312618 400226 313238 400294
rect 312618 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 313238 400226
rect 312618 400102 313238 400170
rect 312618 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 313238 400102
rect 312618 399978 313238 400046
rect 312618 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 313238 399978
rect 301532 382050 301588 382060
rect 312396 396838 312452 396848
rect 312396 382004 312452 396782
rect 312396 381938 312452 381948
rect 312618 382350 313238 399922
rect 316338 406350 316958 408466
rect 316338 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 316958 406350
rect 316338 406226 316958 406294
rect 316338 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 316958 406226
rect 316338 406102 316958 406170
rect 316338 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 316958 406102
rect 316338 405978 316958 406046
rect 316338 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 316958 405978
rect 312618 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 313238 382350
rect 312618 382226 313238 382294
rect 312618 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 313238 382226
rect 312618 382102 313238 382170
rect 312618 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 313238 382102
rect 312618 381978 313238 382046
rect 299852 380752 299908 380762
rect 312618 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 313238 381978
rect 314076 396658 314132 396668
rect 314076 382004 314132 396602
rect 314076 381938 314132 381948
rect 315756 391078 315812 391088
rect 315756 382004 315812 391022
rect 315756 381938 315812 381948
rect 316338 388350 316958 405922
rect 339612 407818 339668 407828
rect 316338 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 316958 388350
rect 316338 388226 316958 388294
rect 316338 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 316958 388226
rect 316338 388102 316958 388170
rect 316338 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 316958 388102
rect 316338 387978 316958 388046
rect 316338 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 316958 387978
rect 312618 380638 313238 381922
rect 315756 381358 315812 381368
rect 295596 380572 295652 380582
rect 280476 380392 280532 380402
rect 315756 379764 315812 381302
rect 316338 380638 316958 387922
rect 322588 390538 322644 390548
rect 322588 382004 322644 390482
rect 322588 381938 322644 381948
rect 338604 380638 338660 380648
rect 315756 379698 315812 379708
rect 338492 380458 338548 380468
rect 271248 370350 271568 370384
rect 271248 370294 271318 370350
rect 271374 370294 271442 370350
rect 271498 370294 271568 370350
rect 271248 370226 271568 370294
rect 271248 370170 271318 370226
rect 271374 370170 271442 370226
rect 271498 370170 271568 370226
rect 271248 370102 271568 370170
rect 271248 370046 271318 370102
rect 271374 370046 271442 370102
rect 271498 370046 271568 370102
rect 271248 369978 271568 370046
rect 271248 369922 271318 369978
rect 271374 369922 271442 369978
rect 271498 369922 271568 369978
rect 271248 369888 271568 369922
rect 301968 370350 302288 370384
rect 301968 370294 302038 370350
rect 302094 370294 302162 370350
rect 302218 370294 302288 370350
rect 301968 370226 302288 370294
rect 301968 370170 302038 370226
rect 302094 370170 302162 370226
rect 302218 370170 302288 370226
rect 301968 370102 302288 370170
rect 301968 370046 302038 370102
rect 302094 370046 302162 370102
rect 302218 370046 302288 370102
rect 301968 369978 302288 370046
rect 301968 369922 302038 369978
rect 302094 369922 302162 369978
rect 302218 369922 302288 369978
rect 301968 369888 302288 369922
rect 332688 370350 333008 370384
rect 332688 370294 332758 370350
rect 332814 370294 332882 370350
rect 332938 370294 333008 370350
rect 332688 370226 333008 370294
rect 332688 370170 332758 370226
rect 332814 370170 332882 370226
rect 332938 370170 333008 370226
rect 332688 370102 333008 370170
rect 332688 370046 332758 370102
rect 332814 370046 332882 370102
rect 332938 370046 333008 370102
rect 332688 369978 333008 370046
rect 332688 369922 332758 369978
rect 332814 369922 332882 369978
rect 332938 369922 333008 369978
rect 332688 369888 333008 369922
rect 255888 364350 256208 364384
rect 255888 364294 255958 364350
rect 256014 364294 256082 364350
rect 256138 364294 256208 364350
rect 255888 364226 256208 364294
rect 255888 364170 255958 364226
rect 256014 364170 256082 364226
rect 256138 364170 256208 364226
rect 255888 364102 256208 364170
rect 255888 364046 255958 364102
rect 256014 364046 256082 364102
rect 256138 364046 256208 364102
rect 255888 363978 256208 364046
rect 255888 363922 255958 363978
rect 256014 363922 256082 363978
rect 256138 363922 256208 363978
rect 255888 363888 256208 363922
rect 286608 364350 286928 364384
rect 286608 364294 286678 364350
rect 286734 364294 286802 364350
rect 286858 364294 286928 364350
rect 286608 364226 286928 364294
rect 286608 364170 286678 364226
rect 286734 364170 286802 364226
rect 286858 364170 286928 364226
rect 286608 364102 286928 364170
rect 286608 364046 286678 364102
rect 286734 364046 286802 364102
rect 286858 364046 286928 364102
rect 286608 363978 286928 364046
rect 286608 363922 286678 363978
rect 286734 363922 286802 363978
rect 286858 363922 286928 363978
rect 286608 363888 286928 363922
rect 317328 364350 317648 364384
rect 317328 364294 317398 364350
rect 317454 364294 317522 364350
rect 317578 364294 317648 364350
rect 317328 364226 317648 364294
rect 317328 364170 317398 364226
rect 317454 364170 317522 364226
rect 317578 364170 317648 364226
rect 317328 364102 317648 364170
rect 317328 364046 317398 364102
rect 317454 364046 317522 364102
rect 317578 364046 317648 364102
rect 317328 363978 317648 364046
rect 317328 363922 317398 363978
rect 317454 363922 317522 363978
rect 317578 363922 317648 363978
rect 317328 363888 317648 363922
rect 271248 352350 271568 352384
rect 271248 352294 271318 352350
rect 271374 352294 271442 352350
rect 271498 352294 271568 352350
rect 271248 352226 271568 352294
rect 271248 352170 271318 352226
rect 271374 352170 271442 352226
rect 271498 352170 271568 352226
rect 271248 352102 271568 352170
rect 271248 352046 271318 352102
rect 271374 352046 271442 352102
rect 271498 352046 271568 352102
rect 271248 351978 271568 352046
rect 271248 351922 271318 351978
rect 271374 351922 271442 351978
rect 271498 351922 271568 351978
rect 271248 351888 271568 351922
rect 301968 352350 302288 352384
rect 301968 352294 302038 352350
rect 302094 352294 302162 352350
rect 302218 352294 302288 352350
rect 301968 352226 302288 352294
rect 301968 352170 302038 352226
rect 302094 352170 302162 352226
rect 302218 352170 302288 352226
rect 301968 352102 302288 352170
rect 301968 352046 302038 352102
rect 302094 352046 302162 352102
rect 302218 352046 302288 352102
rect 301968 351978 302288 352046
rect 301968 351922 302038 351978
rect 302094 351922 302162 351978
rect 302218 351922 302288 351978
rect 301968 351888 302288 351922
rect 332688 352350 333008 352384
rect 332688 352294 332758 352350
rect 332814 352294 332882 352350
rect 332938 352294 333008 352350
rect 332688 352226 333008 352294
rect 332688 352170 332758 352226
rect 332814 352170 332882 352226
rect 332938 352170 333008 352226
rect 332688 352102 333008 352170
rect 332688 352046 332758 352102
rect 332814 352046 332882 352102
rect 332938 352046 333008 352102
rect 332688 351978 333008 352046
rect 332688 351922 332758 351978
rect 332814 351922 332882 351978
rect 332938 351922 333008 351978
rect 332688 351888 333008 351922
rect 255888 346350 256208 346384
rect 255888 346294 255958 346350
rect 256014 346294 256082 346350
rect 256138 346294 256208 346350
rect 255888 346226 256208 346294
rect 255888 346170 255958 346226
rect 256014 346170 256082 346226
rect 256138 346170 256208 346226
rect 255888 346102 256208 346170
rect 255888 346046 255958 346102
rect 256014 346046 256082 346102
rect 256138 346046 256208 346102
rect 255888 345978 256208 346046
rect 255888 345922 255958 345978
rect 256014 345922 256082 345978
rect 256138 345922 256208 345978
rect 255888 345888 256208 345922
rect 286608 346350 286928 346384
rect 286608 346294 286678 346350
rect 286734 346294 286802 346350
rect 286858 346294 286928 346350
rect 286608 346226 286928 346294
rect 286608 346170 286678 346226
rect 286734 346170 286802 346226
rect 286858 346170 286928 346226
rect 286608 346102 286928 346170
rect 286608 346046 286678 346102
rect 286734 346046 286802 346102
rect 286858 346046 286928 346102
rect 286608 345978 286928 346046
rect 286608 345922 286678 345978
rect 286734 345922 286802 345978
rect 286858 345922 286928 345978
rect 286608 345888 286928 345922
rect 317328 346350 317648 346384
rect 317328 346294 317398 346350
rect 317454 346294 317522 346350
rect 317578 346294 317648 346350
rect 317328 346226 317648 346294
rect 317328 346170 317398 346226
rect 317454 346170 317522 346226
rect 317578 346170 317648 346226
rect 317328 346102 317648 346170
rect 317328 346046 317398 346102
rect 317454 346046 317522 346102
rect 317578 346046 317648 346102
rect 317328 345978 317648 346046
rect 317328 345922 317398 345978
rect 317454 345922 317522 345978
rect 317578 345922 317648 345978
rect 317328 345888 317648 345922
rect 338156 342478 338212 342488
rect 271248 334350 271568 334384
rect 271248 334294 271318 334350
rect 271374 334294 271442 334350
rect 271498 334294 271568 334350
rect 271248 334226 271568 334294
rect 271248 334170 271318 334226
rect 271374 334170 271442 334226
rect 271498 334170 271568 334226
rect 271248 334102 271568 334170
rect 271248 334046 271318 334102
rect 271374 334046 271442 334102
rect 271498 334046 271568 334102
rect 271248 333978 271568 334046
rect 271248 333922 271318 333978
rect 271374 333922 271442 333978
rect 271498 333922 271568 333978
rect 271248 333888 271568 333922
rect 301968 334350 302288 334384
rect 301968 334294 302038 334350
rect 302094 334294 302162 334350
rect 302218 334294 302288 334350
rect 301968 334226 302288 334294
rect 301968 334170 302038 334226
rect 302094 334170 302162 334226
rect 302218 334170 302288 334226
rect 301968 334102 302288 334170
rect 301968 334046 302038 334102
rect 302094 334046 302162 334102
rect 302218 334046 302288 334102
rect 301968 333978 302288 334046
rect 301968 333922 302038 333978
rect 302094 333922 302162 333978
rect 302218 333922 302288 333978
rect 301968 333888 302288 333922
rect 332688 334350 333008 334384
rect 332688 334294 332758 334350
rect 332814 334294 332882 334350
rect 332938 334294 333008 334350
rect 332688 334226 333008 334294
rect 332688 334170 332758 334226
rect 332814 334170 332882 334226
rect 332938 334170 333008 334226
rect 332688 334102 333008 334170
rect 332688 334046 332758 334102
rect 332814 334046 332882 334102
rect 332938 334046 333008 334102
rect 332688 333978 333008 334046
rect 332688 333922 332758 333978
rect 332814 333922 332882 333978
rect 332938 333922 333008 333978
rect 332688 333888 333008 333922
rect 255888 328350 256208 328384
rect 255888 328294 255958 328350
rect 256014 328294 256082 328350
rect 256138 328294 256208 328350
rect 255888 328226 256208 328294
rect 255888 328170 255958 328226
rect 256014 328170 256082 328226
rect 256138 328170 256208 328226
rect 255888 328102 256208 328170
rect 255888 328046 255958 328102
rect 256014 328046 256082 328102
rect 256138 328046 256208 328102
rect 255888 327978 256208 328046
rect 255888 327922 255958 327978
rect 256014 327922 256082 327978
rect 256138 327922 256208 327978
rect 255888 327888 256208 327922
rect 286608 328350 286928 328384
rect 286608 328294 286678 328350
rect 286734 328294 286802 328350
rect 286858 328294 286928 328350
rect 286608 328226 286928 328294
rect 286608 328170 286678 328226
rect 286734 328170 286802 328226
rect 286858 328170 286928 328226
rect 286608 328102 286928 328170
rect 286608 328046 286678 328102
rect 286734 328046 286802 328102
rect 286858 328046 286928 328102
rect 286608 327978 286928 328046
rect 286608 327922 286678 327978
rect 286734 327922 286802 327978
rect 286858 327922 286928 327978
rect 286608 327888 286928 327922
rect 317328 328350 317648 328384
rect 317328 328294 317398 328350
rect 317454 328294 317522 328350
rect 317578 328294 317648 328350
rect 317328 328226 317648 328294
rect 317328 328170 317398 328226
rect 317454 328170 317522 328226
rect 317578 328170 317648 328226
rect 317328 328102 317648 328170
rect 317328 328046 317398 328102
rect 317454 328046 317522 328102
rect 317578 328046 317648 328102
rect 317328 327978 317648 328046
rect 317328 327922 317398 327978
rect 317454 327922 317522 327978
rect 317578 327922 317648 327978
rect 317328 327888 317648 327922
rect 271248 316350 271568 316384
rect 271248 316294 271318 316350
rect 271374 316294 271442 316350
rect 271498 316294 271568 316350
rect 271248 316226 271568 316294
rect 271248 316170 271318 316226
rect 271374 316170 271442 316226
rect 271498 316170 271568 316226
rect 271248 316102 271568 316170
rect 271248 316046 271318 316102
rect 271374 316046 271442 316102
rect 271498 316046 271568 316102
rect 271248 315978 271568 316046
rect 271248 315922 271318 315978
rect 271374 315922 271442 315978
rect 271498 315922 271568 315978
rect 271248 315888 271568 315922
rect 301968 316350 302288 316384
rect 301968 316294 302038 316350
rect 302094 316294 302162 316350
rect 302218 316294 302288 316350
rect 301968 316226 302288 316294
rect 301968 316170 302038 316226
rect 302094 316170 302162 316226
rect 302218 316170 302288 316226
rect 301968 316102 302288 316170
rect 301968 316046 302038 316102
rect 302094 316046 302162 316102
rect 302218 316046 302288 316102
rect 301968 315978 302288 316046
rect 301968 315922 302038 315978
rect 302094 315922 302162 315978
rect 302218 315922 302288 315978
rect 301968 315888 302288 315922
rect 332688 316350 333008 316384
rect 332688 316294 332758 316350
rect 332814 316294 332882 316350
rect 332938 316294 333008 316350
rect 332688 316226 333008 316294
rect 332688 316170 332758 316226
rect 332814 316170 332882 316226
rect 332938 316170 333008 316226
rect 332688 316102 333008 316170
rect 332688 316046 332758 316102
rect 332814 316046 332882 316102
rect 332938 316046 333008 316102
rect 332688 315978 333008 316046
rect 332688 315922 332758 315978
rect 332814 315922 332882 315978
rect 332938 315922 333008 315978
rect 332688 315888 333008 315922
rect 255888 310350 256208 310384
rect 255888 310294 255958 310350
rect 256014 310294 256082 310350
rect 256138 310294 256208 310350
rect 255888 310226 256208 310294
rect 255888 310170 255958 310226
rect 256014 310170 256082 310226
rect 256138 310170 256208 310226
rect 255888 310102 256208 310170
rect 255888 310046 255958 310102
rect 256014 310046 256082 310102
rect 256138 310046 256208 310102
rect 255888 309978 256208 310046
rect 255888 309922 255958 309978
rect 256014 309922 256082 309978
rect 256138 309922 256208 309978
rect 255888 309888 256208 309922
rect 286608 310350 286928 310384
rect 286608 310294 286678 310350
rect 286734 310294 286802 310350
rect 286858 310294 286928 310350
rect 286608 310226 286928 310294
rect 286608 310170 286678 310226
rect 286734 310170 286802 310226
rect 286858 310170 286928 310226
rect 286608 310102 286928 310170
rect 286608 310046 286678 310102
rect 286734 310046 286802 310102
rect 286858 310046 286928 310102
rect 286608 309978 286928 310046
rect 286608 309922 286678 309978
rect 286734 309922 286802 309978
rect 286858 309922 286928 309978
rect 286608 309888 286928 309922
rect 317328 310350 317648 310384
rect 317328 310294 317398 310350
rect 317454 310294 317522 310350
rect 317578 310294 317648 310350
rect 317328 310226 317648 310294
rect 317328 310170 317398 310226
rect 317454 310170 317522 310226
rect 317578 310170 317648 310226
rect 317328 310102 317648 310170
rect 317328 310046 317398 310102
rect 317454 310046 317522 310102
rect 317578 310046 317648 310102
rect 317328 309978 317648 310046
rect 317328 309922 317398 309978
rect 317454 309922 317522 309978
rect 317578 309922 317648 309978
rect 317328 309888 317648 309922
rect 271248 298350 271568 298384
rect 271248 298294 271318 298350
rect 271374 298294 271442 298350
rect 271498 298294 271568 298350
rect 271248 298226 271568 298294
rect 271248 298170 271318 298226
rect 271374 298170 271442 298226
rect 271498 298170 271568 298226
rect 271248 298102 271568 298170
rect 271248 298046 271318 298102
rect 271374 298046 271442 298102
rect 271498 298046 271568 298102
rect 271248 297978 271568 298046
rect 271248 297922 271318 297978
rect 271374 297922 271442 297978
rect 271498 297922 271568 297978
rect 271248 297888 271568 297922
rect 301968 298350 302288 298384
rect 301968 298294 302038 298350
rect 302094 298294 302162 298350
rect 302218 298294 302288 298350
rect 301968 298226 302288 298294
rect 301968 298170 302038 298226
rect 302094 298170 302162 298226
rect 302218 298170 302288 298226
rect 301968 298102 302288 298170
rect 301968 298046 302038 298102
rect 302094 298046 302162 298102
rect 302218 298046 302288 298102
rect 301968 297978 302288 298046
rect 301968 297922 302038 297978
rect 302094 297922 302162 297978
rect 302218 297922 302288 297978
rect 301968 297888 302288 297922
rect 332688 298350 333008 298384
rect 332688 298294 332758 298350
rect 332814 298294 332882 298350
rect 332938 298294 333008 298350
rect 332688 298226 333008 298294
rect 332688 298170 332758 298226
rect 332814 298170 332882 298226
rect 332938 298170 333008 298226
rect 332688 298102 333008 298170
rect 332688 298046 332758 298102
rect 332814 298046 332882 298102
rect 332938 298046 333008 298102
rect 332688 297978 333008 298046
rect 332688 297922 332758 297978
rect 332814 297922 332882 297978
rect 332938 297922 333008 297978
rect 332688 297888 333008 297922
rect 255888 292350 256208 292384
rect 255888 292294 255958 292350
rect 256014 292294 256082 292350
rect 256138 292294 256208 292350
rect 255888 292226 256208 292294
rect 255888 292170 255958 292226
rect 256014 292170 256082 292226
rect 256138 292170 256208 292226
rect 255888 292102 256208 292170
rect 255888 292046 255958 292102
rect 256014 292046 256082 292102
rect 256138 292046 256208 292102
rect 255888 291978 256208 292046
rect 255888 291922 255958 291978
rect 256014 291922 256082 291978
rect 256138 291922 256208 291978
rect 255888 291888 256208 291922
rect 286608 292350 286928 292384
rect 286608 292294 286678 292350
rect 286734 292294 286802 292350
rect 286858 292294 286928 292350
rect 286608 292226 286928 292294
rect 286608 292170 286678 292226
rect 286734 292170 286802 292226
rect 286858 292170 286928 292226
rect 286608 292102 286928 292170
rect 286608 292046 286678 292102
rect 286734 292046 286802 292102
rect 286858 292046 286928 292102
rect 286608 291978 286928 292046
rect 286608 291922 286678 291978
rect 286734 291922 286802 291978
rect 286858 291922 286928 291978
rect 286608 291888 286928 291922
rect 317328 292350 317648 292384
rect 317328 292294 317398 292350
rect 317454 292294 317522 292350
rect 317578 292294 317648 292350
rect 317328 292226 317648 292294
rect 317328 292170 317398 292226
rect 317454 292170 317522 292226
rect 317578 292170 317648 292226
rect 317328 292102 317648 292170
rect 317328 292046 317398 292102
rect 317454 292046 317522 292102
rect 317578 292046 317648 292102
rect 317328 291978 317648 292046
rect 317328 291922 317398 291978
rect 317454 291922 317522 291978
rect 317578 291922 317648 291978
rect 317328 291888 317648 291922
rect 271248 280350 271568 280384
rect 271248 280294 271318 280350
rect 271374 280294 271442 280350
rect 271498 280294 271568 280350
rect 271248 280226 271568 280294
rect 271248 280170 271318 280226
rect 271374 280170 271442 280226
rect 271498 280170 271568 280226
rect 271248 280102 271568 280170
rect 271248 280046 271318 280102
rect 271374 280046 271442 280102
rect 271498 280046 271568 280102
rect 271248 279978 271568 280046
rect 271248 279922 271318 279978
rect 271374 279922 271442 279978
rect 271498 279922 271568 279978
rect 271248 279888 271568 279922
rect 301968 280350 302288 280384
rect 301968 280294 302038 280350
rect 302094 280294 302162 280350
rect 302218 280294 302288 280350
rect 301968 280226 302288 280294
rect 301968 280170 302038 280226
rect 302094 280170 302162 280226
rect 302218 280170 302288 280226
rect 301968 280102 302288 280170
rect 301968 280046 302038 280102
rect 302094 280046 302162 280102
rect 302218 280046 302288 280102
rect 301968 279978 302288 280046
rect 301968 279922 302038 279978
rect 302094 279922 302162 279978
rect 302218 279922 302288 279978
rect 301968 279888 302288 279922
rect 332688 280350 333008 280384
rect 332688 280294 332758 280350
rect 332814 280294 332882 280350
rect 332938 280294 333008 280350
rect 332688 280226 333008 280294
rect 332688 280170 332758 280226
rect 332814 280170 332882 280226
rect 332938 280170 333008 280226
rect 332688 280102 333008 280170
rect 332688 280046 332758 280102
rect 332814 280046 332882 280102
rect 332938 280046 333008 280102
rect 332688 279978 333008 280046
rect 332688 279922 332758 279978
rect 332814 279922 332882 279978
rect 332938 279922 333008 279978
rect 332688 279888 333008 279922
rect 255888 274350 256208 274384
rect 255888 274294 255958 274350
rect 256014 274294 256082 274350
rect 256138 274294 256208 274350
rect 255888 274226 256208 274294
rect 255888 274170 255958 274226
rect 256014 274170 256082 274226
rect 256138 274170 256208 274226
rect 255888 274102 256208 274170
rect 255888 274046 255958 274102
rect 256014 274046 256082 274102
rect 256138 274046 256208 274102
rect 255888 273978 256208 274046
rect 255888 273922 255958 273978
rect 256014 273922 256082 273978
rect 256138 273922 256208 273978
rect 255888 273888 256208 273922
rect 286608 274350 286928 274384
rect 286608 274294 286678 274350
rect 286734 274294 286802 274350
rect 286858 274294 286928 274350
rect 286608 274226 286928 274294
rect 286608 274170 286678 274226
rect 286734 274170 286802 274226
rect 286858 274170 286928 274226
rect 286608 274102 286928 274170
rect 286608 274046 286678 274102
rect 286734 274046 286802 274102
rect 286858 274046 286928 274102
rect 286608 273978 286928 274046
rect 286608 273922 286678 273978
rect 286734 273922 286802 273978
rect 286858 273922 286928 273978
rect 286608 273888 286928 273922
rect 317328 274350 317648 274384
rect 317328 274294 317398 274350
rect 317454 274294 317522 274350
rect 317578 274294 317648 274350
rect 317328 274226 317648 274294
rect 317328 274170 317398 274226
rect 317454 274170 317522 274226
rect 317578 274170 317648 274226
rect 317328 274102 317648 274170
rect 317328 274046 317398 274102
rect 317454 274046 317522 274102
rect 317578 274046 317648 274102
rect 317328 273978 317648 274046
rect 317328 273922 317398 273978
rect 317454 273922 317522 273978
rect 317578 273922 317648 273978
rect 317328 273888 317648 273922
rect 271248 262350 271568 262384
rect 271248 262294 271318 262350
rect 271374 262294 271442 262350
rect 271498 262294 271568 262350
rect 271248 262226 271568 262294
rect 271248 262170 271318 262226
rect 271374 262170 271442 262226
rect 271498 262170 271568 262226
rect 271248 262102 271568 262170
rect 271248 262046 271318 262102
rect 271374 262046 271442 262102
rect 271498 262046 271568 262102
rect 271248 261978 271568 262046
rect 271248 261922 271318 261978
rect 271374 261922 271442 261978
rect 271498 261922 271568 261978
rect 271248 261888 271568 261922
rect 301968 262350 302288 262384
rect 301968 262294 302038 262350
rect 302094 262294 302162 262350
rect 302218 262294 302288 262350
rect 301968 262226 302288 262294
rect 301968 262170 302038 262226
rect 302094 262170 302162 262226
rect 302218 262170 302288 262226
rect 301968 262102 302288 262170
rect 301968 262046 302038 262102
rect 302094 262046 302162 262102
rect 302218 262046 302288 262102
rect 301968 261978 302288 262046
rect 301968 261922 302038 261978
rect 302094 261922 302162 261978
rect 302218 261922 302288 261978
rect 301968 261888 302288 261922
rect 332688 262350 333008 262384
rect 332688 262294 332758 262350
rect 332814 262294 332882 262350
rect 332938 262294 333008 262350
rect 332688 262226 333008 262294
rect 332688 262170 332758 262226
rect 332814 262170 332882 262226
rect 332938 262170 333008 262226
rect 332688 262102 333008 262170
rect 332688 262046 332758 262102
rect 332814 262046 332882 262102
rect 332938 262046 333008 262102
rect 332688 261978 333008 262046
rect 332688 261922 332758 261978
rect 332814 261922 332882 261978
rect 332938 261922 333008 261978
rect 332688 261888 333008 261922
rect 255888 256350 256208 256384
rect 255888 256294 255958 256350
rect 256014 256294 256082 256350
rect 256138 256294 256208 256350
rect 255888 256226 256208 256294
rect 255888 256170 255958 256226
rect 256014 256170 256082 256226
rect 256138 256170 256208 256226
rect 255888 256102 256208 256170
rect 255888 256046 255958 256102
rect 256014 256046 256082 256102
rect 256138 256046 256208 256102
rect 255888 255978 256208 256046
rect 255888 255922 255958 255978
rect 256014 255922 256082 255978
rect 256138 255922 256208 255978
rect 255888 255888 256208 255922
rect 286608 256350 286928 256384
rect 286608 256294 286678 256350
rect 286734 256294 286802 256350
rect 286858 256294 286928 256350
rect 286608 256226 286928 256294
rect 286608 256170 286678 256226
rect 286734 256170 286802 256226
rect 286858 256170 286928 256226
rect 286608 256102 286928 256170
rect 286608 256046 286678 256102
rect 286734 256046 286802 256102
rect 286858 256046 286928 256102
rect 286608 255978 286928 256046
rect 286608 255922 286678 255978
rect 286734 255922 286802 255978
rect 286858 255922 286928 255978
rect 286608 255888 286928 255922
rect 317328 256350 317648 256384
rect 317328 256294 317398 256350
rect 317454 256294 317522 256350
rect 317578 256294 317648 256350
rect 317328 256226 317648 256294
rect 317328 256170 317398 256226
rect 317454 256170 317522 256226
rect 317578 256170 317648 256226
rect 317328 256102 317648 256170
rect 317328 256046 317398 256102
rect 317454 256046 317522 256102
rect 317578 256046 317648 256102
rect 317328 255978 317648 256046
rect 317328 255922 317398 255978
rect 317454 255922 317522 255978
rect 317578 255922 317648 255978
rect 317328 255888 317648 255922
rect 338156 250348 338212 342422
rect 338492 314188 338548 380402
rect 338604 317098 338660 380582
rect 339500 363300 339556 363310
rect 339276 347172 339332 347182
rect 339276 342478 339332 347116
rect 339276 342412 339332 342422
rect 338604 317044 339444 317098
rect 338604 317042 339388 317044
rect 339388 316978 339444 316988
rect 338268 314132 338548 314188
rect 338268 301978 338324 314132
rect 339276 309540 339332 309550
rect 339276 309148 339332 309484
rect 338716 309092 339332 309148
rect 338716 305788 338772 309092
rect 338268 301912 338324 301922
rect 338380 305732 338772 305788
rect 338380 253738 338436 305732
rect 339388 301978 339444 301988
rect 339388 298116 339444 301922
rect 339388 298050 339444 298060
rect 339276 286244 339332 286254
rect 339276 285958 339332 286188
rect 338380 253672 338436 253682
rect 338492 285902 339332 285958
rect 337932 250292 338212 250348
rect 337932 244918 337988 250292
rect 338380 249958 338436 249968
rect 337932 244852 337988 244862
rect 338044 249902 338380 249958
rect 271248 244350 271568 244384
rect 271248 244294 271318 244350
rect 271374 244294 271442 244350
rect 271498 244294 271568 244350
rect 271248 244226 271568 244294
rect 271248 244170 271318 244226
rect 271374 244170 271442 244226
rect 271498 244170 271568 244226
rect 271248 244102 271568 244170
rect 271248 244046 271318 244102
rect 271374 244046 271442 244102
rect 271498 244046 271568 244102
rect 271248 243978 271568 244046
rect 271248 243922 271318 243978
rect 271374 243922 271442 243978
rect 271498 243922 271568 243978
rect 271248 243888 271568 243922
rect 301968 244350 302288 244384
rect 301968 244294 302038 244350
rect 302094 244294 302162 244350
rect 302218 244294 302288 244350
rect 301968 244226 302288 244294
rect 301968 244170 302038 244226
rect 302094 244170 302162 244226
rect 302218 244170 302288 244226
rect 301968 244102 302288 244170
rect 301968 244046 302038 244102
rect 302094 244046 302162 244102
rect 302218 244046 302288 244102
rect 301968 243978 302288 244046
rect 301968 243922 302038 243978
rect 302094 243922 302162 243978
rect 302218 243922 302288 243978
rect 301968 243888 302288 243922
rect 332688 244350 333008 244384
rect 332688 244294 332758 244350
rect 332814 244294 332882 244350
rect 332938 244294 333008 244350
rect 332688 244226 333008 244294
rect 332688 244170 332758 244226
rect 332814 244170 332882 244226
rect 332938 244170 333008 244226
rect 332688 244102 333008 244170
rect 332688 244046 332758 244102
rect 332814 244046 332882 244102
rect 332938 244046 333008 244102
rect 332688 243978 333008 244046
rect 332688 243922 332758 243978
rect 332814 243922 332882 243978
rect 332938 243922 333008 243978
rect 332688 243888 333008 243922
rect 336924 241498 336980 241508
rect 289772 241138 289828 241148
rect 241836 239698 241892 239708
rect 244188 238532 244244 238542
rect 243404 237076 243460 237086
rect 241724 234546 241780 234556
rect 241836 236964 241892 236974
rect 241836 227998 241892 236908
rect 241836 227932 241892 227942
rect 243404 224578 243460 237020
rect 244188 236998 244244 238476
rect 245084 238532 245140 238542
rect 245084 237178 245140 238476
rect 245084 237112 245140 237122
rect 251178 238350 251798 240034
rect 281372 239764 281428 239774
rect 273980 239652 274036 239662
rect 251178 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 251798 238350
rect 272972 239540 273028 239550
rect 251178 238226 251798 238294
rect 251178 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 251798 238226
rect 251178 238102 251798 238170
rect 251178 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 251798 238102
rect 251178 237978 251798 238046
rect 251178 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 251798 237978
rect 243404 224512 243460 224522
rect 243516 236964 243572 236974
rect 244188 236932 244244 236942
rect 243516 224398 243572 236908
rect 243516 224332 243572 224342
rect 241052 211012 241108 211022
rect 251178 220350 251798 237922
rect 270508 238308 270564 238318
rect 269836 237178 269892 237188
rect 268716 237076 268772 237086
rect 267036 236964 267092 236974
rect 251178 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 251798 220350
rect 251178 220226 251798 220294
rect 251178 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 251798 220226
rect 251178 220102 251798 220170
rect 251178 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 251798 220102
rect 251178 219978 251798 220046
rect 251178 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 251798 219978
rect 251178 210574 251798 219922
rect 266924 234500 266980 234510
rect 189532 209794 189588 209804
rect 264796 210084 264852 210094
rect 186396 209682 186452 209692
rect 182700 209570 182756 209580
rect 181132 209458 181188 209468
rect 177996 209346 178052 209356
rect 264796 209076 264852 210028
rect 264796 209010 264852 209020
rect 44448 202350 44768 202384
rect 44448 202294 44518 202350
rect 44574 202294 44642 202350
rect 44698 202294 44768 202350
rect 44448 202226 44768 202294
rect 44448 202170 44518 202226
rect 44574 202170 44642 202226
rect 44698 202170 44768 202226
rect 44448 202102 44768 202170
rect 44448 202046 44518 202102
rect 44574 202046 44642 202102
rect 44698 202046 44768 202102
rect 44448 201978 44768 202046
rect 44448 201922 44518 201978
rect 44574 201922 44642 201978
rect 44698 201922 44768 201978
rect 44448 201888 44768 201922
rect 75168 202350 75488 202384
rect 75168 202294 75238 202350
rect 75294 202294 75362 202350
rect 75418 202294 75488 202350
rect 75168 202226 75488 202294
rect 75168 202170 75238 202226
rect 75294 202170 75362 202226
rect 75418 202170 75488 202226
rect 75168 202102 75488 202170
rect 75168 202046 75238 202102
rect 75294 202046 75362 202102
rect 75418 202046 75488 202102
rect 75168 201978 75488 202046
rect 75168 201922 75238 201978
rect 75294 201922 75362 201978
rect 75418 201922 75488 201978
rect 75168 201888 75488 201922
rect 105888 202350 106208 202384
rect 105888 202294 105958 202350
rect 106014 202294 106082 202350
rect 106138 202294 106208 202350
rect 105888 202226 106208 202294
rect 105888 202170 105958 202226
rect 106014 202170 106082 202226
rect 106138 202170 106208 202226
rect 105888 202102 106208 202170
rect 105888 202046 105958 202102
rect 106014 202046 106082 202102
rect 106138 202046 106208 202102
rect 105888 201978 106208 202046
rect 105888 201922 105958 201978
rect 106014 201922 106082 201978
rect 106138 201922 106208 201978
rect 105888 201888 106208 201922
rect 136608 202350 136928 202384
rect 136608 202294 136678 202350
rect 136734 202294 136802 202350
rect 136858 202294 136928 202350
rect 136608 202226 136928 202294
rect 136608 202170 136678 202226
rect 136734 202170 136802 202226
rect 136858 202170 136928 202226
rect 136608 202102 136928 202170
rect 136608 202046 136678 202102
rect 136734 202046 136802 202102
rect 136858 202046 136928 202102
rect 136608 201978 136928 202046
rect 136608 201922 136678 201978
rect 136734 201922 136802 201978
rect 136858 201922 136928 201978
rect 136608 201888 136928 201922
rect 167328 202350 167648 202384
rect 167328 202294 167398 202350
rect 167454 202294 167522 202350
rect 167578 202294 167648 202350
rect 167328 202226 167648 202294
rect 167328 202170 167398 202226
rect 167454 202170 167522 202226
rect 167578 202170 167648 202226
rect 167328 202102 167648 202170
rect 167328 202046 167398 202102
rect 167454 202046 167522 202102
rect 167578 202046 167648 202102
rect 167328 201978 167648 202046
rect 167328 201922 167398 201978
rect 167454 201922 167522 201978
rect 167578 201922 167648 201978
rect 167328 201888 167648 201922
rect 198048 202350 198368 202384
rect 198048 202294 198118 202350
rect 198174 202294 198242 202350
rect 198298 202294 198368 202350
rect 198048 202226 198368 202294
rect 198048 202170 198118 202226
rect 198174 202170 198242 202226
rect 198298 202170 198368 202226
rect 198048 202102 198368 202170
rect 198048 202046 198118 202102
rect 198174 202046 198242 202102
rect 198298 202046 198368 202102
rect 198048 201978 198368 202046
rect 198048 201922 198118 201978
rect 198174 201922 198242 201978
rect 198298 201922 198368 201978
rect 198048 201888 198368 201922
rect 228768 202350 229088 202384
rect 228768 202294 228838 202350
rect 228894 202294 228962 202350
rect 229018 202294 229088 202350
rect 228768 202226 229088 202294
rect 228768 202170 228838 202226
rect 228894 202170 228962 202226
rect 229018 202170 229088 202226
rect 228768 202102 229088 202170
rect 228768 202046 228838 202102
rect 228894 202046 228962 202102
rect 229018 202046 229088 202102
rect 228768 201978 229088 202046
rect 228768 201922 228838 201978
rect 228894 201922 228962 201978
rect 229018 201922 229088 201978
rect 228768 201888 229088 201922
rect 259488 202350 259808 202384
rect 259488 202294 259558 202350
rect 259614 202294 259682 202350
rect 259738 202294 259808 202350
rect 259488 202226 259808 202294
rect 259488 202170 259558 202226
rect 259614 202170 259682 202226
rect 259738 202170 259808 202226
rect 259488 202102 259808 202170
rect 259488 202046 259558 202102
rect 259614 202046 259682 202102
rect 259738 202046 259808 202102
rect 259488 201978 259808 202046
rect 259488 201922 259558 201978
rect 259614 201922 259682 201978
rect 259738 201922 259808 201978
rect 259488 201888 259808 201922
rect 59808 190350 60128 190384
rect 59808 190294 59878 190350
rect 59934 190294 60002 190350
rect 60058 190294 60128 190350
rect 59808 190226 60128 190294
rect 59808 190170 59878 190226
rect 59934 190170 60002 190226
rect 60058 190170 60128 190226
rect 59808 190102 60128 190170
rect 59808 190046 59878 190102
rect 59934 190046 60002 190102
rect 60058 190046 60128 190102
rect 59808 189978 60128 190046
rect 59808 189922 59878 189978
rect 59934 189922 60002 189978
rect 60058 189922 60128 189978
rect 59808 189888 60128 189922
rect 90528 190350 90848 190384
rect 90528 190294 90598 190350
rect 90654 190294 90722 190350
rect 90778 190294 90848 190350
rect 90528 190226 90848 190294
rect 90528 190170 90598 190226
rect 90654 190170 90722 190226
rect 90778 190170 90848 190226
rect 90528 190102 90848 190170
rect 90528 190046 90598 190102
rect 90654 190046 90722 190102
rect 90778 190046 90848 190102
rect 90528 189978 90848 190046
rect 90528 189922 90598 189978
rect 90654 189922 90722 189978
rect 90778 189922 90848 189978
rect 90528 189888 90848 189922
rect 121248 190350 121568 190384
rect 121248 190294 121318 190350
rect 121374 190294 121442 190350
rect 121498 190294 121568 190350
rect 121248 190226 121568 190294
rect 121248 190170 121318 190226
rect 121374 190170 121442 190226
rect 121498 190170 121568 190226
rect 121248 190102 121568 190170
rect 121248 190046 121318 190102
rect 121374 190046 121442 190102
rect 121498 190046 121568 190102
rect 121248 189978 121568 190046
rect 121248 189922 121318 189978
rect 121374 189922 121442 189978
rect 121498 189922 121568 189978
rect 121248 189888 121568 189922
rect 151968 190350 152288 190384
rect 151968 190294 152038 190350
rect 152094 190294 152162 190350
rect 152218 190294 152288 190350
rect 151968 190226 152288 190294
rect 151968 190170 152038 190226
rect 152094 190170 152162 190226
rect 152218 190170 152288 190226
rect 151968 190102 152288 190170
rect 151968 190046 152038 190102
rect 152094 190046 152162 190102
rect 152218 190046 152288 190102
rect 151968 189978 152288 190046
rect 151968 189922 152038 189978
rect 152094 189922 152162 189978
rect 152218 189922 152288 189978
rect 151968 189888 152288 189922
rect 182688 190350 183008 190384
rect 182688 190294 182758 190350
rect 182814 190294 182882 190350
rect 182938 190294 183008 190350
rect 182688 190226 183008 190294
rect 182688 190170 182758 190226
rect 182814 190170 182882 190226
rect 182938 190170 183008 190226
rect 182688 190102 183008 190170
rect 182688 190046 182758 190102
rect 182814 190046 182882 190102
rect 182938 190046 183008 190102
rect 182688 189978 183008 190046
rect 182688 189922 182758 189978
rect 182814 189922 182882 189978
rect 182938 189922 183008 189978
rect 182688 189888 183008 189922
rect 213408 190350 213728 190384
rect 213408 190294 213478 190350
rect 213534 190294 213602 190350
rect 213658 190294 213728 190350
rect 213408 190226 213728 190294
rect 213408 190170 213478 190226
rect 213534 190170 213602 190226
rect 213658 190170 213728 190226
rect 213408 190102 213728 190170
rect 213408 190046 213478 190102
rect 213534 190046 213602 190102
rect 213658 190046 213728 190102
rect 213408 189978 213728 190046
rect 213408 189922 213478 189978
rect 213534 189922 213602 189978
rect 213658 189922 213728 189978
rect 213408 189888 213728 189922
rect 244128 190350 244448 190384
rect 244128 190294 244198 190350
rect 244254 190294 244322 190350
rect 244378 190294 244448 190350
rect 244128 190226 244448 190294
rect 244128 190170 244198 190226
rect 244254 190170 244322 190226
rect 244378 190170 244448 190226
rect 244128 190102 244448 190170
rect 244128 190046 244198 190102
rect 244254 190046 244322 190102
rect 244378 190046 244448 190102
rect 244128 189978 244448 190046
rect 244128 189922 244198 189978
rect 244254 189922 244322 189978
rect 244378 189922 244448 189978
rect 244128 189888 244448 189922
rect 44448 184350 44768 184384
rect 44448 184294 44518 184350
rect 44574 184294 44642 184350
rect 44698 184294 44768 184350
rect 44448 184226 44768 184294
rect 44448 184170 44518 184226
rect 44574 184170 44642 184226
rect 44698 184170 44768 184226
rect 44448 184102 44768 184170
rect 44448 184046 44518 184102
rect 44574 184046 44642 184102
rect 44698 184046 44768 184102
rect 44448 183978 44768 184046
rect 44448 183922 44518 183978
rect 44574 183922 44642 183978
rect 44698 183922 44768 183978
rect 44448 183888 44768 183922
rect 75168 184350 75488 184384
rect 75168 184294 75238 184350
rect 75294 184294 75362 184350
rect 75418 184294 75488 184350
rect 75168 184226 75488 184294
rect 75168 184170 75238 184226
rect 75294 184170 75362 184226
rect 75418 184170 75488 184226
rect 75168 184102 75488 184170
rect 75168 184046 75238 184102
rect 75294 184046 75362 184102
rect 75418 184046 75488 184102
rect 75168 183978 75488 184046
rect 75168 183922 75238 183978
rect 75294 183922 75362 183978
rect 75418 183922 75488 183978
rect 75168 183888 75488 183922
rect 105888 184350 106208 184384
rect 105888 184294 105958 184350
rect 106014 184294 106082 184350
rect 106138 184294 106208 184350
rect 105888 184226 106208 184294
rect 105888 184170 105958 184226
rect 106014 184170 106082 184226
rect 106138 184170 106208 184226
rect 105888 184102 106208 184170
rect 105888 184046 105958 184102
rect 106014 184046 106082 184102
rect 106138 184046 106208 184102
rect 105888 183978 106208 184046
rect 105888 183922 105958 183978
rect 106014 183922 106082 183978
rect 106138 183922 106208 183978
rect 105888 183888 106208 183922
rect 136608 184350 136928 184384
rect 136608 184294 136678 184350
rect 136734 184294 136802 184350
rect 136858 184294 136928 184350
rect 136608 184226 136928 184294
rect 136608 184170 136678 184226
rect 136734 184170 136802 184226
rect 136858 184170 136928 184226
rect 136608 184102 136928 184170
rect 136608 184046 136678 184102
rect 136734 184046 136802 184102
rect 136858 184046 136928 184102
rect 136608 183978 136928 184046
rect 136608 183922 136678 183978
rect 136734 183922 136802 183978
rect 136858 183922 136928 183978
rect 136608 183888 136928 183922
rect 167328 184350 167648 184384
rect 167328 184294 167398 184350
rect 167454 184294 167522 184350
rect 167578 184294 167648 184350
rect 167328 184226 167648 184294
rect 167328 184170 167398 184226
rect 167454 184170 167522 184226
rect 167578 184170 167648 184226
rect 167328 184102 167648 184170
rect 167328 184046 167398 184102
rect 167454 184046 167522 184102
rect 167578 184046 167648 184102
rect 167328 183978 167648 184046
rect 167328 183922 167398 183978
rect 167454 183922 167522 183978
rect 167578 183922 167648 183978
rect 167328 183888 167648 183922
rect 198048 184350 198368 184384
rect 198048 184294 198118 184350
rect 198174 184294 198242 184350
rect 198298 184294 198368 184350
rect 198048 184226 198368 184294
rect 198048 184170 198118 184226
rect 198174 184170 198242 184226
rect 198298 184170 198368 184226
rect 198048 184102 198368 184170
rect 198048 184046 198118 184102
rect 198174 184046 198242 184102
rect 198298 184046 198368 184102
rect 198048 183978 198368 184046
rect 198048 183922 198118 183978
rect 198174 183922 198242 183978
rect 198298 183922 198368 183978
rect 198048 183888 198368 183922
rect 228768 184350 229088 184384
rect 228768 184294 228838 184350
rect 228894 184294 228962 184350
rect 229018 184294 229088 184350
rect 228768 184226 229088 184294
rect 228768 184170 228838 184226
rect 228894 184170 228962 184226
rect 229018 184170 229088 184226
rect 228768 184102 229088 184170
rect 228768 184046 228838 184102
rect 228894 184046 228962 184102
rect 229018 184046 229088 184102
rect 228768 183978 229088 184046
rect 228768 183922 228838 183978
rect 228894 183922 228962 183978
rect 229018 183922 229088 183978
rect 228768 183888 229088 183922
rect 259488 184350 259808 184384
rect 259488 184294 259558 184350
rect 259614 184294 259682 184350
rect 259738 184294 259808 184350
rect 259488 184226 259808 184294
rect 259488 184170 259558 184226
rect 259614 184170 259682 184226
rect 259738 184170 259808 184226
rect 259488 184102 259808 184170
rect 259488 184046 259558 184102
rect 259614 184046 259682 184102
rect 259738 184046 259808 184102
rect 259488 183978 259808 184046
rect 259488 183922 259558 183978
rect 259614 183922 259682 183978
rect 259738 183922 259808 183978
rect 259488 183888 259808 183922
rect 59808 172350 60128 172384
rect 59808 172294 59878 172350
rect 59934 172294 60002 172350
rect 60058 172294 60128 172350
rect 59808 172226 60128 172294
rect 59808 172170 59878 172226
rect 59934 172170 60002 172226
rect 60058 172170 60128 172226
rect 59808 172102 60128 172170
rect 59808 172046 59878 172102
rect 59934 172046 60002 172102
rect 60058 172046 60128 172102
rect 59808 171978 60128 172046
rect 59808 171922 59878 171978
rect 59934 171922 60002 171978
rect 60058 171922 60128 171978
rect 59808 171888 60128 171922
rect 90528 172350 90848 172384
rect 90528 172294 90598 172350
rect 90654 172294 90722 172350
rect 90778 172294 90848 172350
rect 90528 172226 90848 172294
rect 90528 172170 90598 172226
rect 90654 172170 90722 172226
rect 90778 172170 90848 172226
rect 90528 172102 90848 172170
rect 90528 172046 90598 172102
rect 90654 172046 90722 172102
rect 90778 172046 90848 172102
rect 90528 171978 90848 172046
rect 90528 171922 90598 171978
rect 90654 171922 90722 171978
rect 90778 171922 90848 171978
rect 90528 171888 90848 171922
rect 121248 172350 121568 172384
rect 121248 172294 121318 172350
rect 121374 172294 121442 172350
rect 121498 172294 121568 172350
rect 121248 172226 121568 172294
rect 121248 172170 121318 172226
rect 121374 172170 121442 172226
rect 121498 172170 121568 172226
rect 121248 172102 121568 172170
rect 121248 172046 121318 172102
rect 121374 172046 121442 172102
rect 121498 172046 121568 172102
rect 121248 171978 121568 172046
rect 121248 171922 121318 171978
rect 121374 171922 121442 171978
rect 121498 171922 121568 171978
rect 121248 171888 121568 171922
rect 151968 172350 152288 172384
rect 151968 172294 152038 172350
rect 152094 172294 152162 172350
rect 152218 172294 152288 172350
rect 151968 172226 152288 172294
rect 151968 172170 152038 172226
rect 152094 172170 152162 172226
rect 152218 172170 152288 172226
rect 151968 172102 152288 172170
rect 151968 172046 152038 172102
rect 152094 172046 152162 172102
rect 152218 172046 152288 172102
rect 151968 171978 152288 172046
rect 151968 171922 152038 171978
rect 152094 171922 152162 171978
rect 152218 171922 152288 171978
rect 151968 171888 152288 171922
rect 182688 172350 183008 172384
rect 182688 172294 182758 172350
rect 182814 172294 182882 172350
rect 182938 172294 183008 172350
rect 182688 172226 183008 172294
rect 182688 172170 182758 172226
rect 182814 172170 182882 172226
rect 182938 172170 183008 172226
rect 182688 172102 183008 172170
rect 182688 172046 182758 172102
rect 182814 172046 182882 172102
rect 182938 172046 183008 172102
rect 182688 171978 183008 172046
rect 182688 171922 182758 171978
rect 182814 171922 182882 171978
rect 182938 171922 183008 171978
rect 182688 171888 183008 171922
rect 213408 172350 213728 172384
rect 213408 172294 213478 172350
rect 213534 172294 213602 172350
rect 213658 172294 213728 172350
rect 213408 172226 213728 172294
rect 213408 172170 213478 172226
rect 213534 172170 213602 172226
rect 213658 172170 213728 172226
rect 213408 172102 213728 172170
rect 213408 172046 213478 172102
rect 213534 172046 213602 172102
rect 213658 172046 213728 172102
rect 213408 171978 213728 172046
rect 213408 171922 213478 171978
rect 213534 171922 213602 171978
rect 213658 171922 213728 171978
rect 213408 171888 213728 171922
rect 244128 172350 244448 172384
rect 244128 172294 244198 172350
rect 244254 172294 244322 172350
rect 244378 172294 244448 172350
rect 244128 172226 244448 172294
rect 244128 172170 244198 172226
rect 244254 172170 244322 172226
rect 244378 172170 244448 172226
rect 244128 172102 244448 172170
rect 244128 172046 244198 172102
rect 244254 172046 244322 172102
rect 244378 172046 244448 172102
rect 244128 171978 244448 172046
rect 244128 171922 244198 171978
rect 244254 171922 244322 171978
rect 244378 171922 244448 171978
rect 244128 171888 244448 171922
rect 44448 166350 44768 166384
rect 44448 166294 44518 166350
rect 44574 166294 44642 166350
rect 44698 166294 44768 166350
rect 44448 166226 44768 166294
rect 44448 166170 44518 166226
rect 44574 166170 44642 166226
rect 44698 166170 44768 166226
rect 44448 166102 44768 166170
rect 44448 166046 44518 166102
rect 44574 166046 44642 166102
rect 44698 166046 44768 166102
rect 44448 165978 44768 166046
rect 44448 165922 44518 165978
rect 44574 165922 44642 165978
rect 44698 165922 44768 165978
rect 44448 165888 44768 165922
rect 75168 166350 75488 166384
rect 75168 166294 75238 166350
rect 75294 166294 75362 166350
rect 75418 166294 75488 166350
rect 75168 166226 75488 166294
rect 75168 166170 75238 166226
rect 75294 166170 75362 166226
rect 75418 166170 75488 166226
rect 75168 166102 75488 166170
rect 75168 166046 75238 166102
rect 75294 166046 75362 166102
rect 75418 166046 75488 166102
rect 75168 165978 75488 166046
rect 75168 165922 75238 165978
rect 75294 165922 75362 165978
rect 75418 165922 75488 165978
rect 75168 165888 75488 165922
rect 105888 166350 106208 166384
rect 105888 166294 105958 166350
rect 106014 166294 106082 166350
rect 106138 166294 106208 166350
rect 105888 166226 106208 166294
rect 105888 166170 105958 166226
rect 106014 166170 106082 166226
rect 106138 166170 106208 166226
rect 105888 166102 106208 166170
rect 105888 166046 105958 166102
rect 106014 166046 106082 166102
rect 106138 166046 106208 166102
rect 105888 165978 106208 166046
rect 105888 165922 105958 165978
rect 106014 165922 106082 165978
rect 106138 165922 106208 165978
rect 105888 165888 106208 165922
rect 136608 166350 136928 166384
rect 136608 166294 136678 166350
rect 136734 166294 136802 166350
rect 136858 166294 136928 166350
rect 136608 166226 136928 166294
rect 136608 166170 136678 166226
rect 136734 166170 136802 166226
rect 136858 166170 136928 166226
rect 136608 166102 136928 166170
rect 136608 166046 136678 166102
rect 136734 166046 136802 166102
rect 136858 166046 136928 166102
rect 136608 165978 136928 166046
rect 136608 165922 136678 165978
rect 136734 165922 136802 165978
rect 136858 165922 136928 165978
rect 136608 165888 136928 165922
rect 167328 166350 167648 166384
rect 167328 166294 167398 166350
rect 167454 166294 167522 166350
rect 167578 166294 167648 166350
rect 167328 166226 167648 166294
rect 167328 166170 167398 166226
rect 167454 166170 167522 166226
rect 167578 166170 167648 166226
rect 167328 166102 167648 166170
rect 167328 166046 167398 166102
rect 167454 166046 167522 166102
rect 167578 166046 167648 166102
rect 167328 165978 167648 166046
rect 167328 165922 167398 165978
rect 167454 165922 167522 165978
rect 167578 165922 167648 165978
rect 167328 165888 167648 165922
rect 198048 166350 198368 166384
rect 198048 166294 198118 166350
rect 198174 166294 198242 166350
rect 198298 166294 198368 166350
rect 198048 166226 198368 166294
rect 198048 166170 198118 166226
rect 198174 166170 198242 166226
rect 198298 166170 198368 166226
rect 198048 166102 198368 166170
rect 198048 166046 198118 166102
rect 198174 166046 198242 166102
rect 198298 166046 198368 166102
rect 198048 165978 198368 166046
rect 198048 165922 198118 165978
rect 198174 165922 198242 165978
rect 198298 165922 198368 165978
rect 198048 165888 198368 165922
rect 228768 166350 229088 166384
rect 228768 166294 228838 166350
rect 228894 166294 228962 166350
rect 229018 166294 229088 166350
rect 228768 166226 229088 166294
rect 228768 166170 228838 166226
rect 228894 166170 228962 166226
rect 229018 166170 229088 166226
rect 228768 166102 229088 166170
rect 228768 166046 228838 166102
rect 228894 166046 228962 166102
rect 229018 166046 229088 166102
rect 228768 165978 229088 166046
rect 228768 165922 228838 165978
rect 228894 165922 228962 165978
rect 229018 165922 229088 165978
rect 228768 165888 229088 165922
rect 259488 166350 259808 166384
rect 259488 166294 259558 166350
rect 259614 166294 259682 166350
rect 259738 166294 259808 166350
rect 259488 166226 259808 166294
rect 259488 166170 259558 166226
rect 259614 166170 259682 166226
rect 259738 166170 259808 166226
rect 259488 166102 259808 166170
rect 259488 166046 259558 166102
rect 259614 166046 259682 166102
rect 259738 166046 259808 166102
rect 259488 165978 259808 166046
rect 259488 165922 259558 165978
rect 259614 165922 259682 165978
rect 259738 165922 259808 165978
rect 259488 165888 259808 165922
rect 59808 154350 60128 154384
rect 59808 154294 59878 154350
rect 59934 154294 60002 154350
rect 60058 154294 60128 154350
rect 59808 154226 60128 154294
rect 59808 154170 59878 154226
rect 59934 154170 60002 154226
rect 60058 154170 60128 154226
rect 59808 154102 60128 154170
rect 59808 154046 59878 154102
rect 59934 154046 60002 154102
rect 60058 154046 60128 154102
rect 59808 153978 60128 154046
rect 59808 153922 59878 153978
rect 59934 153922 60002 153978
rect 60058 153922 60128 153978
rect 59808 153888 60128 153922
rect 90528 154350 90848 154384
rect 90528 154294 90598 154350
rect 90654 154294 90722 154350
rect 90778 154294 90848 154350
rect 90528 154226 90848 154294
rect 90528 154170 90598 154226
rect 90654 154170 90722 154226
rect 90778 154170 90848 154226
rect 90528 154102 90848 154170
rect 90528 154046 90598 154102
rect 90654 154046 90722 154102
rect 90778 154046 90848 154102
rect 90528 153978 90848 154046
rect 90528 153922 90598 153978
rect 90654 153922 90722 153978
rect 90778 153922 90848 153978
rect 90528 153888 90848 153922
rect 121248 154350 121568 154384
rect 121248 154294 121318 154350
rect 121374 154294 121442 154350
rect 121498 154294 121568 154350
rect 121248 154226 121568 154294
rect 121248 154170 121318 154226
rect 121374 154170 121442 154226
rect 121498 154170 121568 154226
rect 121248 154102 121568 154170
rect 121248 154046 121318 154102
rect 121374 154046 121442 154102
rect 121498 154046 121568 154102
rect 121248 153978 121568 154046
rect 121248 153922 121318 153978
rect 121374 153922 121442 153978
rect 121498 153922 121568 153978
rect 121248 153888 121568 153922
rect 151968 154350 152288 154384
rect 151968 154294 152038 154350
rect 152094 154294 152162 154350
rect 152218 154294 152288 154350
rect 151968 154226 152288 154294
rect 151968 154170 152038 154226
rect 152094 154170 152162 154226
rect 152218 154170 152288 154226
rect 151968 154102 152288 154170
rect 151968 154046 152038 154102
rect 152094 154046 152162 154102
rect 152218 154046 152288 154102
rect 151968 153978 152288 154046
rect 151968 153922 152038 153978
rect 152094 153922 152162 153978
rect 152218 153922 152288 153978
rect 151968 153888 152288 153922
rect 182688 154350 183008 154384
rect 182688 154294 182758 154350
rect 182814 154294 182882 154350
rect 182938 154294 183008 154350
rect 182688 154226 183008 154294
rect 182688 154170 182758 154226
rect 182814 154170 182882 154226
rect 182938 154170 183008 154226
rect 182688 154102 183008 154170
rect 182688 154046 182758 154102
rect 182814 154046 182882 154102
rect 182938 154046 183008 154102
rect 182688 153978 183008 154046
rect 182688 153922 182758 153978
rect 182814 153922 182882 153978
rect 182938 153922 183008 153978
rect 182688 153888 183008 153922
rect 213408 154350 213728 154384
rect 213408 154294 213478 154350
rect 213534 154294 213602 154350
rect 213658 154294 213728 154350
rect 213408 154226 213728 154294
rect 213408 154170 213478 154226
rect 213534 154170 213602 154226
rect 213658 154170 213728 154226
rect 213408 154102 213728 154170
rect 213408 154046 213478 154102
rect 213534 154046 213602 154102
rect 213658 154046 213728 154102
rect 213408 153978 213728 154046
rect 213408 153922 213478 153978
rect 213534 153922 213602 153978
rect 213658 153922 213728 153978
rect 213408 153888 213728 153922
rect 244128 154350 244448 154384
rect 244128 154294 244198 154350
rect 244254 154294 244322 154350
rect 244378 154294 244448 154350
rect 244128 154226 244448 154294
rect 244128 154170 244198 154226
rect 244254 154170 244322 154226
rect 244378 154170 244448 154226
rect 244128 154102 244448 154170
rect 244128 154046 244198 154102
rect 244254 154046 244322 154102
rect 244378 154046 244448 154102
rect 244128 153978 244448 154046
rect 244128 153922 244198 153978
rect 244254 153922 244322 153978
rect 244378 153922 244448 153978
rect 244128 153888 244448 153922
rect 44448 148350 44768 148384
rect 44448 148294 44518 148350
rect 44574 148294 44642 148350
rect 44698 148294 44768 148350
rect 44448 148226 44768 148294
rect 44448 148170 44518 148226
rect 44574 148170 44642 148226
rect 44698 148170 44768 148226
rect 44448 148102 44768 148170
rect 44448 148046 44518 148102
rect 44574 148046 44642 148102
rect 44698 148046 44768 148102
rect 44448 147978 44768 148046
rect 44448 147922 44518 147978
rect 44574 147922 44642 147978
rect 44698 147922 44768 147978
rect 44448 147888 44768 147922
rect 75168 148350 75488 148384
rect 75168 148294 75238 148350
rect 75294 148294 75362 148350
rect 75418 148294 75488 148350
rect 75168 148226 75488 148294
rect 75168 148170 75238 148226
rect 75294 148170 75362 148226
rect 75418 148170 75488 148226
rect 75168 148102 75488 148170
rect 75168 148046 75238 148102
rect 75294 148046 75362 148102
rect 75418 148046 75488 148102
rect 75168 147978 75488 148046
rect 75168 147922 75238 147978
rect 75294 147922 75362 147978
rect 75418 147922 75488 147978
rect 75168 147888 75488 147922
rect 105888 148350 106208 148384
rect 105888 148294 105958 148350
rect 106014 148294 106082 148350
rect 106138 148294 106208 148350
rect 105888 148226 106208 148294
rect 105888 148170 105958 148226
rect 106014 148170 106082 148226
rect 106138 148170 106208 148226
rect 105888 148102 106208 148170
rect 105888 148046 105958 148102
rect 106014 148046 106082 148102
rect 106138 148046 106208 148102
rect 105888 147978 106208 148046
rect 105888 147922 105958 147978
rect 106014 147922 106082 147978
rect 106138 147922 106208 147978
rect 105888 147888 106208 147922
rect 136608 148350 136928 148384
rect 136608 148294 136678 148350
rect 136734 148294 136802 148350
rect 136858 148294 136928 148350
rect 136608 148226 136928 148294
rect 136608 148170 136678 148226
rect 136734 148170 136802 148226
rect 136858 148170 136928 148226
rect 136608 148102 136928 148170
rect 136608 148046 136678 148102
rect 136734 148046 136802 148102
rect 136858 148046 136928 148102
rect 136608 147978 136928 148046
rect 136608 147922 136678 147978
rect 136734 147922 136802 147978
rect 136858 147922 136928 147978
rect 136608 147888 136928 147922
rect 167328 148350 167648 148384
rect 167328 148294 167398 148350
rect 167454 148294 167522 148350
rect 167578 148294 167648 148350
rect 167328 148226 167648 148294
rect 167328 148170 167398 148226
rect 167454 148170 167522 148226
rect 167578 148170 167648 148226
rect 167328 148102 167648 148170
rect 167328 148046 167398 148102
rect 167454 148046 167522 148102
rect 167578 148046 167648 148102
rect 167328 147978 167648 148046
rect 167328 147922 167398 147978
rect 167454 147922 167522 147978
rect 167578 147922 167648 147978
rect 167328 147888 167648 147922
rect 198048 148350 198368 148384
rect 198048 148294 198118 148350
rect 198174 148294 198242 148350
rect 198298 148294 198368 148350
rect 198048 148226 198368 148294
rect 198048 148170 198118 148226
rect 198174 148170 198242 148226
rect 198298 148170 198368 148226
rect 198048 148102 198368 148170
rect 198048 148046 198118 148102
rect 198174 148046 198242 148102
rect 198298 148046 198368 148102
rect 198048 147978 198368 148046
rect 198048 147922 198118 147978
rect 198174 147922 198242 147978
rect 198298 147922 198368 147978
rect 198048 147888 198368 147922
rect 228768 148350 229088 148384
rect 228768 148294 228838 148350
rect 228894 148294 228962 148350
rect 229018 148294 229088 148350
rect 228768 148226 229088 148294
rect 228768 148170 228838 148226
rect 228894 148170 228962 148226
rect 229018 148170 229088 148226
rect 228768 148102 229088 148170
rect 228768 148046 228838 148102
rect 228894 148046 228962 148102
rect 229018 148046 229088 148102
rect 228768 147978 229088 148046
rect 228768 147922 228838 147978
rect 228894 147922 228962 147978
rect 229018 147922 229088 147978
rect 228768 147888 229088 147922
rect 259488 148350 259808 148384
rect 259488 148294 259558 148350
rect 259614 148294 259682 148350
rect 259738 148294 259808 148350
rect 259488 148226 259808 148294
rect 259488 148170 259558 148226
rect 259614 148170 259682 148226
rect 259738 148170 259808 148226
rect 259488 148102 259808 148170
rect 259488 148046 259558 148102
rect 259614 148046 259682 148102
rect 259738 148046 259808 148102
rect 259488 147978 259808 148046
rect 259488 147922 259558 147978
rect 259614 147922 259682 147978
rect 259738 147922 259808 147978
rect 259488 147888 259808 147922
rect 59808 136350 60128 136384
rect 59808 136294 59878 136350
rect 59934 136294 60002 136350
rect 60058 136294 60128 136350
rect 59808 136226 60128 136294
rect 59808 136170 59878 136226
rect 59934 136170 60002 136226
rect 60058 136170 60128 136226
rect 59808 136102 60128 136170
rect 59808 136046 59878 136102
rect 59934 136046 60002 136102
rect 60058 136046 60128 136102
rect 59808 135978 60128 136046
rect 59808 135922 59878 135978
rect 59934 135922 60002 135978
rect 60058 135922 60128 135978
rect 59808 135888 60128 135922
rect 90528 136350 90848 136384
rect 90528 136294 90598 136350
rect 90654 136294 90722 136350
rect 90778 136294 90848 136350
rect 90528 136226 90848 136294
rect 90528 136170 90598 136226
rect 90654 136170 90722 136226
rect 90778 136170 90848 136226
rect 90528 136102 90848 136170
rect 90528 136046 90598 136102
rect 90654 136046 90722 136102
rect 90778 136046 90848 136102
rect 90528 135978 90848 136046
rect 90528 135922 90598 135978
rect 90654 135922 90722 135978
rect 90778 135922 90848 135978
rect 90528 135888 90848 135922
rect 121248 136350 121568 136384
rect 121248 136294 121318 136350
rect 121374 136294 121442 136350
rect 121498 136294 121568 136350
rect 121248 136226 121568 136294
rect 121248 136170 121318 136226
rect 121374 136170 121442 136226
rect 121498 136170 121568 136226
rect 121248 136102 121568 136170
rect 121248 136046 121318 136102
rect 121374 136046 121442 136102
rect 121498 136046 121568 136102
rect 121248 135978 121568 136046
rect 121248 135922 121318 135978
rect 121374 135922 121442 135978
rect 121498 135922 121568 135978
rect 121248 135888 121568 135922
rect 151968 136350 152288 136384
rect 151968 136294 152038 136350
rect 152094 136294 152162 136350
rect 152218 136294 152288 136350
rect 151968 136226 152288 136294
rect 151968 136170 152038 136226
rect 152094 136170 152162 136226
rect 152218 136170 152288 136226
rect 151968 136102 152288 136170
rect 151968 136046 152038 136102
rect 152094 136046 152162 136102
rect 152218 136046 152288 136102
rect 151968 135978 152288 136046
rect 151968 135922 152038 135978
rect 152094 135922 152162 135978
rect 152218 135922 152288 135978
rect 151968 135888 152288 135922
rect 182688 136350 183008 136384
rect 182688 136294 182758 136350
rect 182814 136294 182882 136350
rect 182938 136294 183008 136350
rect 182688 136226 183008 136294
rect 182688 136170 182758 136226
rect 182814 136170 182882 136226
rect 182938 136170 183008 136226
rect 182688 136102 183008 136170
rect 182688 136046 182758 136102
rect 182814 136046 182882 136102
rect 182938 136046 183008 136102
rect 182688 135978 183008 136046
rect 182688 135922 182758 135978
rect 182814 135922 182882 135978
rect 182938 135922 183008 135978
rect 182688 135888 183008 135922
rect 213408 136350 213728 136384
rect 213408 136294 213478 136350
rect 213534 136294 213602 136350
rect 213658 136294 213728 136350
rect 213408 136226 213728 136294
rect 213408 136170 213478 136226
rect 213534 136170 213602 136226
rect 213658 136170 213728 136226
rect 213408 136102 213728 136170
rect 213408 136046 213478 136102
rect 213534 136046 213602 136102
rect 213658 136046 213728 136102
rect 213408 135978 213728 136046
rect 213408 135922 213478 135978
rect 213534 135922 213602 135978
rect 213658 135922 213728 135978
rect 213408 135888 213728 135922
rect 244128 136350 244448 136384
rect 244128 136294 244198 136350
rect 244254 136294 244322 136350
rect 244378 136294 244448 136350
rect 244128 136226 244448 136294
rect 244128 136170 244198 136226
rect 244254 136170 244322 136226
rect 244378 136170 244448 136226
rect 244128 136102 244448 136170
rect 244128 136046 244198 136102
rect 244254 136046 244322 136102
rect 244378 136046 244448 136102
rect 244128 135978 244448 136046
rect 244128 135922 244198 135978
rect 244254 135922 244322 135978
rect 244378 135922 244448 135978
rect 244128 135888 244448 135922
rect 44448 130350 44768 130384
rect 44448 130294 44518 130350
rect 44574 130294 44642 130350
rect 44698 130294 44768 130350
rect 44448 130226 44768 130294
rect 44448 130170 44518 130226
rect 44574 130170 44642 130226
rect 44698 130170 44768 130226
rect 44448 130102 44768 130170
rect 44448 130046 44518 130102
rect 44574 130046 44642 130102
rect 44698 130046 44768 130102
rect 44448 129978 44768 130046
rect 44448 129922 44518 129978
rect 44574 129922 44642 129978
rect 44698 129922 44768 129978
rect 44448 129888 44768 129922
rect 75168 130350 75488 130384
rect 75168 130294 75238 130350
rect 75294 130294 75362 130350
rect 75418 130294 75488 130350
rect 75168 130226 75488 130294
rect 75168 130170 75238 130226
rect 75294 130170 75362 130226
rect 75418 130170 75488 130226
rect 75168 130102 75488 130170
rect 75168 130046 75238 130102
rect 75294 130046 75362 130102
rect 75418 130046 75488 130102
rect 75168 129978 75488 130046
rect 75168 129922 75238 129978
rect 75294 129922 75362 129978
rect 75418 129922 75488 129978
rect 75168 129888 75488 129922
rect 105888 130350 106208 130384
rect 105888 130294 105958 130350
rect 106014 130294 106082 130350
rect 106138 130294 106208 130350
rect 105888 130226 106208 130294
rect 105888 130170 105958 130226
rect 106014 130170 106082 130226
rect 106138 130170 106208 130226
rect 105888 130102 106208 130170
rect 105888 130046 105958 130102
rect 106014 130046 106082 130102
rect 106138 130046 106208 130102
rect 105888 129978 106208 130046
rect 105888 129922 105958 129978
rect 106014 129922 106082 129978
rect 106138 129922 106208 129978
rect 105888 129888 106208 129922
rect 136608 130350 136928 130384
rect 136608 130294 136678 130350
rect 136734 130294 136802 130350
rect 136858 130294 136928 130350
rect 136608 130226 136928 130294
rect 136608 130170 136678 130226
rect 136734 130170 136802 130226
rect 136858 130170 136928 130226
rect 136608 130102 136928 130170
rect 136608 130046 136678 130102
rect 136734 130046 136802 130102
rect 136858 130046 136928 130102
rect 136608 129978 136928 130046
rect 136608 129922 136678 129978
rect 136734 129922 136802 129978
rect 136858 129922 136928 129978
rect 136608 129888 136928 129922
rect 167328 130350 167648 130384
rect 167328 130294 167398 130350
rect 167454 130294 167522 130350
rect 167578 130294 167648 130350
rect 167328 130226 167648 130294
rect 167328 130170 167398 130226
rect 167454 130170 167522 130226
rect 167578 130170 167648 130226
rect 167328 130102 167648 130170
rect 167328 130046 167398 130102
rect 167454 130046 167522 130102
rect 167578 130046 167648 130102
rect 167328 129978 167648 130046
rect 167328 129922 167398 129978
rect 167454 129922 167522 129978
rect 167578 129922 167648 129978
rect 167328 129888 167648 129922
rect 198048 130350 198368 130384
rect 198048 130294 198118 130350
rect 198174 130294 198242 130350
rect 198298 130294 198368 130350
rect 198048 130226 198368 130294
rect 198048 130170 198118 130226
rect 198174 130170 198242 130226
rect 198298 130170 198368 130226
rect 198048 130102 198368 130170
rect 198048 130046 198118 130102
rect 198174 130046 198242 130102
rect 198298 130046 198368 130102
rect 198048 129978 198368 130046
rect 198048 129922 198118 129978
rect 198174 129922 198242 129978
rect 198298 129922 198368 129978
rect 198048 129888 198368 129922
rect 228768 130350 229088 130384
rect 228768 130294 228838 130350
rect 228894 130294 228962 130350
rect 229018 130294 229088 130350
rect 228768 130226 229088 130294
rect 228768 130170 228838 130226
rect 228894 130170 228962 130226
rect 229018 130170 229088 130226
rect 228768 130102 229088 130170
rect 228768 130046 228838 130102
rect 228894 130046 228962 130102
rect 229018 130046 229088 130102
rect 228768 129978 229088 130046
rect 228768 129922 228838 129978
rect 228894 129922 228962 129978
rect 229018 129922 229088 129978
rect 228768 129888 229088 129922
rect 259488 130350 259808 130384
rect 259488 130294 259558 130350
rect 259614 130294 259682 130350
rect 259738 130294 259808 130350
rect 259488 130226 259808 130294
rect 259488 130170 259558 130226
rect 259614 130170 259682 130226
rect 259738 130170 259808 130226
rect 259488 130102 259808 130170
rect 259488 130046 259558 130102
rect 259614 130046 259682 130102
rect 259738 130046 259808 130102
rect 259488 129978 259808 130046
rect 259488 129922 259558 129978
rect 259614 129922 259682 129978
rect 259738 129922 259808 129978
rect 259488 129888 259808 129922
rect 59808 118350 60128 118384
rect 59808 118294 59878 118350
rect 59934 118294 60002 118350
rect 60058 118294 60128 118350
rect 59808 118226 60128 118294
rect 59808 118170 59878 118226
rect 59934 118170 60002 118226
rect 60058 118170 60128 118226
rect 59808 118102 60128 118170
rect 59808 118046 59878 118102
rect 59934 118046 60002 118102
rect 60058 118046 60128 118102
rect 59808 117978 60128 118046
rect 59808 117922 59878 117978
rect 59934 117922 60002 117978
rect 60058 117922 60128 117978
rect 59808 117888 60128 117922
rect 90528 118350 90848 118384
rect 90528 118294 90598 118350
rect 90654 118294 90722 118350
rect 90778 118294 90848 118350
rect 90528 118226 90848 118294
rect 90528 118170 90598 118226
rect 90654 118170 90722 118226
rect 90778 118170 90848 118226
rect 90528 118102 90848 118170
rect 90528 118046 90598 118102
rect 90654 118046 90722 118102
rect 90778 118046 90848 118102
rect 90528 117978 90848 118046
rect 90528 117922 90598 117978
rect 90654 117922 90722 117978
rect 90778 117922 90848 117978
rect 90528 117888 90848 117922
rect 121248 118350 121568 118384
rect 121248 118294 121318 118350
rect 121374 118294 121442 118350
rect 121498 118294 121568 118350
rect 121248 118226 121568 118294
rect 121248 118170 121318 118226
rect 121374 118170 121442 118226
rect 121498 118170 121568 118226
rect 121248 118102 121568 118170
rect 121248 118046 121318 118102
rect 121374 118046 121442 118102
rect 121498 118046 121568 118102
rect 121248 117978 121568 118046
rect 121248 117922 121318 117978
rect 121374 117922 121442 117978
rect 121498 117922 121568 117978
rect 121248 117888 121568 117922
rect 151968 118350 152288 118384
rect 151968 118294 152038 118350
rect 152094 118294 152162 118350
rect 152218 118294 152288 118350
rect 151968 118226 152288 118294
rect 151968 118170 152038 118226
rect 152094 118170 152162 118226
rect 152218 118170 152288 118226
rect 151968 118102 152288 118170
rect 151968 118046 152038 118102
rect 152094 118046 152162 118102
rect 152218 118046 152288 118102
rect 151968 117978 152288 118046
rect 151968 117922 152038 117978
rect 152094 117922 152162 117978
rect 152218 117922 152288 117978
rect 151968 117888 152288 117922
rect 182688 118350 183008 118384
rect 182688 118294 182758 118350
rect 182814 118294 182882 118350
rect 182938 118294 183008 118350
rect 182688 118226 183008 118294
rect 182688 118170 182758 118226
rect 182814 118170 182882 118226
rect 182938 118170 183008 118226
rect 182688 118102 183008 118170
rect 182688 118046 182758 118102
rect 182814 118046 182882 118102
rect 182938 118046 183008 118102
rect 182688 117978 183008 118046
rect 182688 117922 182758 117978
rect 182814 117922 182882 117978
rect 182938 117922 183008 117978
rect 182688 117888 183008 117922
rect 213408 118350 213728 118384
rect 213408 118294 213478 118350
rect 213534 118294 213602 118350
rect 213658 118294 213728 118350
rect 213408 118226 213728 118294
rect 213408 118170 213478 118226
rect 213534 118170 213602 118226
rect 213658 118170 213728 118226
rect 213408 118102 213728 118170
rect 213408 118046 213478 118102
rect 213534 118046 213602 118102
rect 213658 118046 213728 118102
rect 213408 117978 213728 118046
rect 213408 117922 213478 117978
rect 213534 117922 213602 117978
rect 213658 117922 213728 117978
rect 213408 117888 213728 117922
rect 244128 118350 244448 118384
rect 244128 118294 244198 118350
rect 244254 118294 244322 118350
rect 244378 118294 244448 118350
rect 244128 118226 244448 118294
rect 244128 118170 244198 118226
rect 244254 118170 244322 118226
rect 244378 118170 244448 118226
rect 244128 118102 244448 118170
rect 244128 118046 244198 118102
rect 244254 118046 244322 118102
rect 244378 118046 244448 118102
rect 244128 117978 244448 118046
rect 244128 117922 244198 117978
rect 244254 117922 244322 117978
rect 244378 117922 244448 117978
rect 244128 117888 244448 117922
rect 44448 112350 44768 112384
rect 44448 112294 44518 112350
rect 44574 112294 44642 112350
rect 44698 112294 44768 112350
rect 44448 112226 44768 112294
rect 44448 112170 44518 112226
rect 44574 112170 44642 112226
rect 44698 112170 44768 112226
rect 44448 112102 44768 112170
rect 44448 112046 44518 112102
rect 44574 112046 44642 112102
rect 44698 112046 44768 112102
rect 44448 111978 44768 112046
rect 44448 111922 44518 111978
rect 44574 111922 44642 111978
rect 44698 111922 44768 111978
rect 44448 111888 44768 111922
rect 75168 112350 75488 112384
rect 75168 112294 75238 112350
rect 75294 112294 75362 112350
rect 75418 112294 75488 112350
rect 75168 112226 75488 112294
rect 75168 112170 75238 112226
rect 75294 112170 75362 112226
rect 75418 112170 75488 112226
rect 75168 112102 75488 112170
rect 75168 112046 75238 112102
rect 75294 112046 75362 112102
rect 75418 112046 75488 112102
rect 75168 111978 75488 112046
rect 75168 111922 75238 111978
rect 75294 111922 75362 111978
rect 75418 111922 75488 111978
rect 75168 111888 75488 111922
rect 105888 112350 106208 112384
rect 105888 112294 105958 112350
rect 106014 112294 106082 112350
rect 106138 112294 106208 112350
rect 105888 112226 106208 112294
rect 105888 112170 105958 112226
rect 106014 112170 106082 112226
rect 106138 112170 106208 112226
rect 105888 112102 106208 112170
rect 105888 112046 105958 112102
rect 106014 112046 106082 112102
rect 106138 112046 106208 112102
rect 105888 111978 106208 112046
rect 105888 111922 105958 111978
rect 106014 111922 106082 111978
rect 106138 111922 106208 111978
rect 105888 111888 106208 111922
rect 136608 112350 136928 112384
rect 136608 112294 136678 112350
rect 136734 112294 136802 112350
rect 136858 112294 136928 112350
rect 136608 112226 136928 112294
rect 136608 112170 136678 112226
rect 136734 112170 136802 112226
rect 136858 112170 136928 112226
rect 136608 112102 136928 112170
rect 136608 112046 136678 112102
rect 136734 112046 136802 112102
rect 136858 112046 136928 112102
rect 136608 111978 136928 112046
rect 136608 111922 136678 111978
rect 136734 111922 136802 111978
rect 136858 111922 136928 111978
rect 136608 111888 136928 111922
rect 167328 112350 167648 112384
rect 167328 112294 167398 112350
rect 167454 112294 167522 112350
rect 167578 112294 167648 112350
rect 167328 112226 167648 112294
rect 167328 112170 167398 112226
rect 167454 112170 167522 112226
rect 167578 112170 167648 112226
rect 167328 112102 167648 112170
rect 167328 112046 167398 112102
rect 167454 112046 167522 112102
rect 167578 112046 167648 112102
rect 167328 111978 167648 112046
rect 167328 111922 167398 111978
rect 167454 111922 167522 111978
rect 167578 111922 167648 111978
rect 167328 111888 167648 111922
rect 198048 112350 198368 112384
rect 198048 112294 198118 112350
rect 198174 112294 198242 112350
rect 198298 112294 198368 112350
rect 198048 112226 198368 112294
rect 198048 112170 198118 112226
rect 198174 112170 198242 112226
rect 198298 112170 198368 112226
rect 198048 112102 198368 112170
rect 198048 112046 198118 112102
rect 198174 112046 198242 112102
rect 198298 112046 198368 112102
rect 198048 111978 198368 112046
rect 198048 111922 198118 111978
rect 198174 111922 198242 111978
rect 198298 111922 198368 111978
rect 198048 111888 198368 111922
rect 228768 112350 229088 112384
rect 228768 112294 228838 112350
rect 228894 112294 228962 112350
rect 229018 112294 229088 112350
rect 228768 112226 229088 112294
rect 228768 112170 228838 112226
rect 228894 112170 228962 112226
rect 229018 112170 229088 112226
rect 228768 112102 229088 112170
rect 228768 112046 228838 112102
rect 228894 112046 228962 112102
rect 229018 112046 229088 112102
rect 228768 111978 229088 112046
rect 228768 111922 228838 111978
rect 228894 111922 228962 111978
rect 229018 111922 229088 111978
rect 228768 111888 229088 111922
rect 259488 112350 259808 112384
rect 259488 112294 259558 112350
rect 259614 112294 259682 112350
rect 259738 112294 259808 112350
rect 259488 112226 259808 112294
rect 259488 112170 259558 112226
rect 259614 112170 259682 112226
rect 259738 112170 259808 112226
rect 259488 112102 259808 112170
rect 259488 112046 259558 112102
rect 259614 112046 259682 112102
rect 259738 112046 259808 112102
rect 259488 111978 259808 112046
rect 259488 111922 259558 111978
rect 259614 111922 259682 111978
rect 259738 111922 259808 111978
rect 259488 111888 259808 111922
rect 59808 100350 60128 100384
rect 59808 100294 59878 100350
rect 59934 100294 60002 100350
rect 60058 100294 60128 100350
rect 59808 100226 60128 100294
rect 59808 100170 59878 100226
rect 59934 100170 60002 100226
rect 60058 100170 60128 100226
rect 59808 100102 60128 100170
rect 59808 100046 59878 100102
rect 59934 100046 60002 100102
rect 60058 100046 60128 100102
rect 59808 99978 60128 100046
rect 59808 99922 59878 99978
rect 59934 99922 60002 99978
rect 60058 99922 60128 99978
rect 59808 99888 60128 99922
rect 90528 100350 90848 100384
rect 90528 100294 90598 100350
rect 90654 100294 90722 100350
rect 90778 100294 90848 100350
rect 90528 100226 90848 100294
rect 90528 100170 90598 100226
rect 90654 100170 90722 100226
rect 90778 100170 90848 100226
rect 90528 100102 90848 100170
rect 90528 100046 90598 100102
rect 90654 100046 90722 100102
rect 90778 100046 90848 100102
rect 90528 99978 90848 100046
rect 90528 99922 90598 99978
rect 90654 99922 90722 99978
rect 90778 99922 90848 99978
rect 90528 99888 90848 99922
rect 121248 100350 121568 100384
rect 121248 100294 121318 100350
rect 121374 100294 121442 100350
rect 121498 100294 121568 100350
rect 121248 100226 121568 100294
rect 121248 100170 121318 100226
rect 121374 100170 121442 100226
rect 121498 100170 121568 100226
rect 121248 100102 121568 100170
rect 121248 100046 121318 100102
rect 121374 100046 121442 100102
rect 121498 100046 121568 100102
rect 121248 99978 121568 100046
rect 121248 99922 121318 99978
rect 121374 99922 121442 99978
rect 121498 99922 121568 99978
rect 121248 99888 121568 99922
rect 151968 100350 152288 100384
rect 151968 100294 152038 100350
rect 152094 100294 152162 100350
rect 152218 100294 152288 100350
rect 151968 100226 152288 100294
rect 151968 100170 152038 100226
rect 152094 100170 152162 100226
rect 152218 100170 152288 100226
rect 151968 100102 152288 100170
rect 151968 100046 152038 100102
rect 152094 100046 152162 100102
rect 152218 100046 152288 100102
rect 151968 99978 152288 100046
rect 151968 99922 152038 99978
rect 152094 99922 152162 99978
rect 152218 99922 152288 99978
rect 151968 99888 152288 99922
rect 182688 100350 183008 100384
rect 182688 100294 182758 100350
rect 182814 100294 182882 100350
rect 182938 100294 183008 100350
rect 182688 100226 183008 100294
rect 182688 100170 182758 100226
rect 182814 100170 182882 100226
rect 182938 100170 183008 100226
rect 182688 100102 183008 100170
rect 182688 100046 182758 100102
rect 182814 100046 182882 100102
rect 182938 100046 183008 100102
rect 182688 99978 183008 100046
rect 182688 99922 182758 99978
rect 182814 99922 182882 99978
rect 182938 99922 183008 99978
rect 182688 99888 183008 99922
rect 213408 100350 213728 100384
rect 213408 100294 213478 100350
rect 213534 100294 213602 100350
rect 213658 100294 213728 100350
rect 213408 100226 213728 100294
rect 213408 100170 213478 100226
rect 213534 100170 213602 100226
rect 213658 100170 213728 100226
rect 213408 100102 213728 100170
rect 213408 100046 213478 100102
rect 213534 100046 213602 100102
rect 213658 100046 213728 100102
rect 213408 99978 213728 100046
rect 213408 99922 213478 99978
rect 213534 99922 213602 99978
rect 213658 99922 213728 99978
rect 213408 99888 213728 99922
rect 244128 100350 244448 100384
rect 244128 100294 244198 100350
rect 244254 100294 244322 100350
rect 244378 100294 244448 100350
rect 244128 100226 244448 100294
rect 244128 100170 244198 100226
rect 244254 100170 244322 100226
rect 244378 100170 244448 100226
rect 244128 100102 244448 100170
rect 244128 100046 244198 100102
rect 244254 100046 244322 100102
rect 244378 100046 244448 100102
rect 244128 99978 244448 100046
rect 244128 99922 244198 99978
rect 244254 99922 244322 99978
rect 244378 99922 244448 99978
rect 244128 99888 244448 99922
rect 44448 94350 44768 94384
rect 44448 94294 44518 94350
rect 44574 94294 44642 94350
rect 44698 94294 44768 94350
rect 44448 94226 44768 94294
rect 44448 94170 44518 94226
rect 44574 94170 44642 94226
rect 44698 94170 44768 94226
rect 44448 94102 44768 94170
rect 44448 94046 44518 94102
rect 44574 94046 44642 94102
rect 44698 94046 44768 94102
rect 44448 93978 44768 94046
rect 44448 93922 44518 93978
rect 44574 93922 44642 93978
rect 44698 93922 44768 93978
rect 44448 93888 44768 93922
rect 75168 94350 75488 94384
rect 75168 94294 75238 94350
rect 75294 94294 75362 94350
rect 75418 94294 75488 94350
rect 75168 94226 75488 94294
rect 75168 94170 75238 94226
rect 75294 94170 75362 94226
rect 75418 94170 75488 94226
rect 75168 94102 75488 94170
rect 75168 94046 75238 94102
rect 75294 94046 75362 94102
rect 75418 94046 75488 94102
rect 75168 93978 75488 94046
rect 75168 93922 75238 93978
rect 75294 93922 75362 93978
rect 75418 93922 75488 93978
rect 75168 93888 75488 93922
rect 105888 94350 106208 94384
rect 105888 94294 105958 94350
rect 106014 94294 106082 94350
rect 106138 94294 106208 94350
rect 105888 94226 106208 94294
rect 105888 94170 105958 94226
rect 106014 94170 106082 94226
rect 106138 94170 106208 94226
rect 105888 94102 106208 94170
rect 105888 94046 105958 94102
rect 106014 94046 106082 94102
rect 106138 94046 106208 94102
rect 105888 93978 106208 94046
rect 105888 93922 105958 93978
rect 106014 93922 106082 93978
rect 106138 93922 106208 93978
rect 105888 93888 106208 93922
rect 136608 94350 136928 94384
rect 136608 94294 136678 94350
rect 136734 94294 136802 94350
rect 136858 94294 136928 94350
rect 136608 94226 136928 94294
rect 136608 94170 136678 94226
rect 136734 94170 136802 94226
rect 136858 94170 136928 94226
rect 136608 94102 136928 94170
rect 136608 94046 136678 94102
rect 136734 94046 136802 94102
rect 136858 94046 136928 94102
rect 136608 93978 136928 94046
rect 136608 93922 136678 93978
rect 136734 93922 136802 93978
rect 136858 93922 136928 93978
rect 136608 93888 136928 93922
rect 167328 94350 167648 94384
rect 167328 94294 167398 94350
rect 167454 94294 167522 94350
rect 167578 94294 167648 94350
rect 167328 94226 167648 94294
rect 167328 94170 167398 94226
rect 167454 94170 167522 94226
rect 167578 94170 167648 94226
rect 167328 94102 167648 94170
rect 167328 94046 167398 94102
rect 167454 94046 167522 94102
rect 167578 94046 167648 94102
rect 167328 93978 167648 94046
rect 167328 93922 167398 93978
rect 167454 93922 167522 93978
rect 167578 93922 167648 93978
rect 167328 93888 167648 93922
rect 198048 94350 198368 94384
rect 198048 94294 198118 94350
rect 198174 94294 198242 94350
rect 198298 94294 198368 94350
rect 198048 94226 198368 94294
rect 198048 94170 198118 94226
rect 198174 94170 198242 94226
rect 198298 94170 198368 94226
rect 198048 94102 198368 94170
rect 198048 94046 198118 94102
rect 198174 94046 198242 94102
rect 198298 94046 198368 94102
rect 198048 93978 198368 94046
rect 198048 93922 198118 93978
rect 198174 93922 198242 93978
rect 198298 93922 198368 93978
rect 198048 93888 198368 93922
rect 228768 94350 229088 94384
rect 228768 94294 228838 94350
rect 228894 94294 228962 94350
rect 229018 94294 229088 94350
rect 228768 94226 229088 94294
rect 228768 94170 228838 94226
rect 228894 94170 228962 94226
rect 229018 94170 229088 94226
rect 228768 94102 229088 94170
rect 228768 94046 228838 94102
rect 228894 94046 228962 94102
rect 229018 94046 229088 94102
rect 228768 93978 229088 94046
rect 228768 93922 228838 93978
rect 228894 93922 228962 93978
rect 229018 93922 229088 93978
rect 228768 93888 229088 93922
rect 259488 94350 259808 94384
rect 259488 94294 259558 94350
rect 259614 94294 259682 94350
rect 259738 94294 259808 94350
rect 259488 94226 259808 94294
rect 259488 94170 259558 94226
rect 259614 94170 259682 94226
rect 259738 94170 259808 94226
rect 259488 94102 259808 94170
rect 259488 94046 259558 94102
rect 259614 94046 259682 94102
rect 259738 94046 259808 94102
rect 259488 93978 259808 94046
rect 259488 93922 259558 93978
rect 259614 93922 259682 93978
rect 259738 93922 259808 93978
rect 259488 93888 259808 93922
rect 59808 82350 60128 82384
rect 59808 82294 59878 82350
rect 59934 82294 60002 82350
rect 60058 82294 60128 82350
rect 59808 82226 60128 82294
rect 59808 82170 59878 82226
rect 59934 82170 60002 82226
rect 60058 82170 60128 82226
rect 59808 82102 60128 82170
rect 59808 82046 59878 82102
rect 59934 82046 60002 82102
rect 60058 82046 60128 82102
rect 59808 81978 60128 82046
rect 59808 81922 59878 81978
rect 59934 81922 60002 81978
rect 60058 81922 60128 81978
rect 59808 81888 60128 81922
rect 90528 82350 90848 82384
rect 90528 82294 90598 82350
rect 90654 82294 90722 82350
rect 90778 82294 90848 82350
rect 90528 82226 90848 82294
rect 90528 82170 90598 82226
rect 90654 82170 90722 82226
rect 90778 82170 90848 82226
rect 90528 82102 90848 82170
rect 90528 82046 90598 82102
rect 90654 82046 90722 82102
rect 90778 82046 90848 82102
rect 90528 81978 90848 82046
rect 90528 81922 90598 81978
rect 90654 81922 90722 81978
rect 90778 81922 90848 81978
rect 90528 81888 90848 81922
rect 121248 82350 121568 82384
rect 121248 82294 121318 82350
rect 121374 82294 121442 82350
rect 121498 82294 121568 82350
rect 121248 82226 121568 82294
rect 121248 82170 121318 82226
rect 121374 82170 121442 82226
rect 121498 82170 121568 82226
rect 121248 82102 121568 82170
rect 121248 82046 121318 82102
rect 121374 82046 121442 82102
rect 121498 82046 121568 82102
rect 121248 81978 121568 82046
rect 121248 81922 121318 81978
rect 121374 81922 121442 81978
rect 121498 81922 121568 81978
rect 121248 81888 121568 81922
rect 151968 82350 152288 82384
rect 151968 82294 152038 82350
rect 152094 82294 152162 82350
rect 152218 82294 152288 82350
rect 151968 82226 152288 82294
rect 151968 82170 152038 82226
rect 152094 82170 152162 82226
rect 152218 82170 152288 82226
rect 151968 82102 152288 82170
rect 151968 82046 152038 82102
rect 152094 82046 152162 82102
rect 152218 82046 152288 82102
rect 151968 81978 152288 82046
rect 151968 81922 152038 81978
rect 152094 81922 152162 81978
rect 152218 81922 152288 81978
rect 151968 81888 152288 81922
rect 182688 82350 183008 82384
rect 182688 82294 182758 82350
rect 182814 82294 182882 82350
rect 182938 82294 183008 82350
rect 182688 82226 183008 82294
rect 182688 82170 182758 82226
rect 182814 82170 182882 82226
rect 182938 82170 183008 82226
rect 182688 82102 183008 82170
rect 182688 82046 182758 82102
rect 182814 82046 182882 82102
rect 182938 82046 183008 82102
rect 182688 81978 183008 82046
rect 182688 81922 182758 81978
rect 182814 81922 182882 81978
rect 182938 81922 183008 81978
rect 182688 81888 183008 81922
rect 213408 82350 213728 82384
rect 213408 82294 213478 82350
rect 213534 82294 213602 82350
rect 213658 82294 213728 82350
rect 213408 82226 213728 82294
rect 213408 82170 213478 82226
rect 213534 82170 213602 82226
rect 213658 82170 213728 82226
rect 213408 82102 213728 82170
rect 213408 82046 213478 82102
rect 213534 82046 213602 82102
rect 213658 82046 213728 82102
rect 213408 81978 213728 82046
rect 213408 81922 213478 81978
rect 213534 81922 213602 81978
rect 213658 81922 213728 81978
rect 213408 81888 213728 81922
rect 244128 82350 244448 82384
rect 244128 82294 244198 82350
rect 244254 82294 244322 82350
rect 244378 82294 244448 82350
rect 244128 82226 244448 82294
rect 244128 82170 244198 82226
rect 244254 82170 244322 82226
rect 244378 82170 244448 82226
rect 244128 82102 244448 82170
rect 244128 82046 244198 82102
rect 244254 82046 244322 82102
rect 244378 82046 244448 82102
rect 244128 81978 244448 82046
rect 244128 81922 244198 81978
rect 244254 81922 244322 81978
rect 244378 81922 244448 81978
rect 244128 81888 244448 81922
rect 44448 76350 44768 76384
rect 44448 76294 44518 76350
rect 44574 76294 44642 76350
rect 44698 76294 44768 76350
rect 44448 76226 44768 76294
rect 44448 76170 44518 76226
rect 44574 76170 44642 76226
rect 44698 76170 44768 76226
rect 44448 76102 44768 76170
rect 44448 76046 44518 76102
rect 44574 76046 44642 76102
rect 44698 76046 44768 76102
rect 44448 75978 44768 76046
rect 44448 75922 44518 75978
rect 44574 75922 44642 75978
rect 44698 75922 44768 75978
rect 44448 75888 44768 75922
rect 75168 76350 75488 76384
rect 75168 76294 75238 76350
rect 75294 76294 75362 76350
rect 75418 76294 75488 76350
rect 75168 76226 75488 76294
rect 75168 76170 75238 76226
rect 75294 76170 75362 76226
rect 75418 76170 75488 76226
rect 75168 76102 75488 76170
rect 75168 76046 75238 76102
rect 75294 76046 75362 76102
rect 75418 76046 75488 76102
rect 75168 75978 75488 76046
rect 75168 75922 75238 75978
rect 75294 75922 75362 75978
rect 75418 75922 75488 75978
rect 75168 75888 75488 75922
rect 105888 76350 106208 76384
rect 105888 76294 105958 76350
rect 106014 76294 106082 76350
rect 106138 76294 106208 76350
rect 105888 76226 106208 76294
rect 105888 76170 105958 76226
rect 106014 76170 106082 76226
rect 106138 76170 106208 76226
rect 105888 76102 106208 76170
rect 105888 76046 105958 76102
rect 106014 76046 106082 76102
rect 106138 76046 106208 76102
rect 105888 75978 106208 76046
rect 105888 75922 105958 75978
rect 106014 75922 106082 75978
rect 106138 75922 106208 75978
rect 105888 75888 106208 75922
rect 136608 76350 136928 76384
rect 136608 76294 136678 76350
rect 136734 76294 136802 76350
rect 136858 76294 136928 76350
rect 136608 76226 136928 76294
rect 136608 76170 136678 76226
rect 136734 76170 136802 76226
rect 136858 76170 136928 76226
rect 136608 76102 136928 76170
rect 136608 76046 136678 76102
rect 136734 76046 136802 76102
rect 136858 76046 136928 76102
rect 136608 75978 136928 76046
rect 136608 75922 136678 75978
rect 136734 75922 136802 75978
rect 136858 75922 136928 75978
rect 136608 75888 136928 75922
rect 167328 76350 167648 76384
rect 167328 76294 167398 76350
rect 167454 76294 167522 76350
rect 167578 76294 167648 76350
rect 167328 76226 167648 76294
rect 167328 76170 167398 76226
rect 167454 76170 167522 76226
rect 167578 76170 167648 76226
rect 167328 76102 167648 76170
rect 167328 76046 167398 76102
rect 167454 76046 167522 76102
rect 167578 76046 167648 76102
rect 167328 75978 167648 76046
rect 167328 75922 167398 75978
rect 167454 75922 167522 75978
rect 167578 75922 167648 75978
rect 167328 75888 167648 75922
rect 198048 76350 198368 76384
rect 198048 76294 198118 76350
rect 198174 76294 198242 76350
rect 198298 76294 198368 76350
rect 198048 76226 198368 76294
rect 198048 76170 198118 76226
rect 198174 76170 198242 76226
rect 198298 76170 198368 76226
rect 198048 76102 198368 76170
rect 198048 76046 198118 76102
rect 198174 76046 198242 76102
rect 198298 76046 198368 76102
rect 198048 75978 198368 76046
rect 198048 75922 198118 75978
rect 198174 75922 198242 75978
rect 198298 75922 198368 75978
rect 198048 75888 198368 75922
rect 228768 76350 229088 76384
rect 228768 76294 228838 76350
rect 228894 76294 228962 76350
rect 229018 76294 229088 76350
rect 228768 76226 229088 76294
rect 228768 76170 228838 76226
rect 228894 76170 228962 76226
rect 229018 76170 229088 76226
rect 228768 76102 229088 76170
rect 228768 76046 228838 76102
rect 228894 76046 228962 76102
rect 229018 76046 229088 76102
rect 228768 75978 229088 76046
rect 228768 75922 228838 75978
rect 228894 75922 228962 75978
rect 229018 75922 229088 75978
rect 228768 75888 229088 75922
rect 259488 76350 259808 76384
rect 259488 76294 259558 76350
rect 259614 76294 259682 76350
rect 259738 76294 259808 76350
rect 259488 76226 259808 76294
rect 259488 76170 259558 76226
rect 259614 76170 259682 76226
rect 259738 76170 259808 76226
rect 259488 76102 259808 76170
rect 259488 76046 259558 76102
rect 259614 76046 259682 76102
rect 259738 76046 259808 76102
rect 259488 75978 259808 76046
rect 259488 75922 259558 75978
rect 259614 75922 259682 75978
rect 259738 75922 259808 75978
rect 259488 75888 259808 75922
rect 59808 64350 60128 64384
rect 59808 64294 59878 64350
rect 59934 64294 60002 64350
rect 60058 64294 60128 64350
rect 59808 64226 60128 64294
rect 59808 64170 59878 64226
rect 59934 64170 60002 64226
rect 60058 64170 60128 64226
rect 59808 64102 60128 64170
rect 59808 64046 59878 64102
rect 59934 64046 60002 64102
rect 60058 64046 60128 64102
rect 59808 63978 60128 64046
rect 59808 63922 59878 63978
rect 59934 63922 60002 63978
rect 60058 63922 60128 63978
rect 59808 63888 60128 63922
rect 90528 64350 90848 64384
rect 90528 64294 90598 64350
rect 90654 64294 90722 64350
rect 90778 64294 90848 64350
rect 90528 64226 90848 64294
rect 90528 64170 90598 64226
rect 90654 64170 90722 64226
rect 90778 64170 90848 64226
rect 90528 64102 90848 64170
rect 90528 64046 90598 64102
rect 90654 64046 90722 64102
rect 90778 64046 90848 64102
rect 90528 63978 90848 64046
rect 90528 63922 90598 63978
rect 90654 63922 90722 63978
rect 90778 63922 90848 63978
rect 90528 63888 90848 63922
rect 121248 64350 121568 64384
rect 121248 64294 121318 64350
rect 121374 64294 121442 64350
rect 121498 64294 121568 64350
rect 121248 64226 121568 64294
rect 121248 64170 121318 64226
rect 121374 64170 121442 64226
rect 121498 64170 121568 64226
rect 121248 64102 121568 64170
rect 121248 64046 121318 64102
rect 121374 64046 121442 64102
rect 121498 64046 121568 64102
rect 121248 63978 121568 64046
rect 121248 63922 121318 63978
rect 121374 63922 121442 63978
rect 121498 63922 121568 63978
rect 121248 63888 121568 63922
rect 151968 64350 152288 64384
rect 151968 64294 152038 64350
rect 152094 64294 152162 64350
rect 152218 64294 152288 64350
rect 151968 64226 152288 64294
rect 151968 64170 152038 64226
rect 152094 64170 152162 64226
rect 152218 64170 152288 64226
rect 151968 64102 152288 64170
rect 151968 64046 152038 64102
rect 152094 64046 152162 64102
rect 152218 64046 152288 64102
rect 151968 63978 152288 64046
rect 151968 63922 152038 63978
rect 152094 63922 152162 63978
rect 152218 63922 152288 63978
rect 151968 63888 152288 63922
rect 182688 64350 183008 64384
rect 182688 64294 182758 64350
rect 182814 64294 182882 64350
rect 182938 64294 183008 64350
rect 182688 64226 183008 64294
rect 182688 64170 182758 64226
rect 182814 64170 182882 64226
rect 182938 64170 183008 64226
rect 182688 64102 183008 64170
rect 182688 64046 182758 64102
rect 182814 64046 182882 64102
rect 182938 64046 183008 64102
rect 182688 63978 183008 64046
rect 182688 63922 182758 63978
rect 182814 63922 182882 63978
rect 182938 63922 183008 63978
rect 182688 63888 183008 63922
rect 213408 64350 213728 64384
rect 213408 64294 213478 64350
rect 213534 64294 213602 64350
rect 213658 64294 213728 64350
rect 213408 64226 213728 64294
rect 213408 64170 213478 64226
rect 213534 64170 213602 64226
rect 213658 64170 213728 64226
rect 213408 64102 213728 64170
rect 213408 64046 213478 64102
rect 213534 64046 213602 64102
rect 213658 64046 213728 64102
rect 213408 63978 213728 64046
rect 213408 63922 213478 63978
rect 213534 63922 213602 63978
rect 213658 63922 213728 63978
rect 213408 63888 213728 63922
rect 244128 64350 244448 64384
rect 244128 64294 244198 64350
rect 244254 64294 244322 64350
rect 244378 64294 244448 64350
rect 244128 64226 244448 64294
rect 244128 64170 244198 64226
rect 244254 64170 244322 64226
rect 244378 64170 244448 64226
rect 244128 64102 244448 64170
rect 244128 64046 244198 64102
rect 244254 64046 244322 64102
rect 244378 64046 244448 64102
rect 244128 63978 244448 64046
rect 244128 63922 244198 63978
rect 244254 63922 244322 63978
rect 244378 63922 244448 63978
rect 244128 63888 244448 63922
rect 44448 58350 44768 58384
rect 44448 58294 44518 58350
rect 44574 58294 44642 58350
rect 44698 58294 44768 58350
rect 44448 58226 44768 58294
rect 44448 58170 44518 58226
rect 44574 58170 44642 58226
rect 44698 58170 44768 58226
rect 44448 58102 44768 58170
rect 44448 58046 44518 58102
rect 44574 58046 44642 58102
rect 44698 58046 44768 58102
rect 44448 57978 44768 58046
rect 44448 57922 44518 57978
rect 44574 57922 44642 57978
rect 44698 57922 44768 57978
rect 44448 57888 44768 57922
rect 75168 58350 75488 58384
rect 75168 58294 75238 58350
rect 75294 58294 75362 58350
rect 75418 58294 75488 58350
rect 75168 58226 75488 58294
rect 75168 58170 75238 58226
rect 75294 58170 75362 58226
rect 75418 58170 75488 58226
rect 75168 58102 75488 58170
rect 75168 58046 75238 58102
rect 75294 58046 75362 58102
rect 75418 58046 75488 58102
rect 75168 57978 75488 58046
rect 75168 57922 75238 57978
rect 75294 57922 75362 57978
rect 75418 57922 75488 57978
rect 75168 57888 75488 57922
rect 105888 58350 106208 58384
rect 105888 58294 105958 58350
rect 106014 58294 106082 58350
rect 106138 58294 106208 58350
rect 105888 58226 106208 58294
rect 105888 58170 105958 58226
rect 106014 58170 106082 58226
rect 106138 58170 106208 58226
rect 105888 58102 106208 58170
rect 105888 58046 105958 58102
rect 106014 58046 106082 58102
rect 106138 58046 106208 58102
rect 105888 57978 106208 58046
rect 105888 57922 105958 57978
rect 106014 57922 106082 57978
rect 106138 57922 106208 57978
rect 105888 57888 106208 57922
rect 136608 58350 136928 58384
rect 136608 58294 136678 58350
rect 136734 58294 136802 58350
rect 136858 58294 136928 58350
rect 136608 58226 136928 58294
rect 136608 58170 136678 58226
rect 136734 58170 136802 58226
rect 136858 58170 136928 58226
rect 136608 58102 136928 58170
rect 136608 58046 136678 58102
rect 136734 58046 136802 58102
rect 136858 58046 136928 58102
rect 136608 57978 136928 58046
rect 136608 57922 136678 57978
rect 136734 57922 136802 57978
rect 136858 57922 136928 57978
rect 136608 57888 136928 57922
rect 167328 58350 167648 58384
rect 167328 58294 167398 58350
rect 167454 58294 167522 58350
rect 167578 58294 167648 58350
rect 167328 58226 167648 58294
rect 167328 58170 167398 58226
rect 167454 58170 167522 58226
rect 167578 58170 167648 58226
rect 167328 58102 167648 58170
rect 167328 58046 167398 58102
rect 167454 58046 167522 58102
rect 167578 58046 167648 58102
rect 167328 57978 167648 58046
rect 167328 57922 167398 57978
rect 167454 57922 167522 57978
rect 167578 57922 167648 57978
rect 167328 57888 167648 57922
rect 198048 58350 198368 58384
rect 198048 58294 198118 58350
rect 198174 58294 198242 58350
rect 198298 58294 198368 58350
rect 198048 58226 198368 58294
rect 198048 58170 198118 58226
rect 198174 58170 198242 58226
rect 198298 58170 198368 58226
rect 198048 58102 198368 58170
rect 198048 58046 198118 58102
rect 198174 58046 198242 58102
rect 198298 58046 198368 58102
rect 198048 57978 198368 58046
rect 198048 57922 198118 57978
rect 198174 57922 198242 57978
rect 198298 57922 198368 57978
rect 198048 57888 198368 57922
rect 228768 58350 229088 58384
rect 228768 58294 228838 58350
rect 228894 58294 228962 58350
rect 229018 58294 229088 58350
rect 228768 58226 229088 58294
rect 228768 58170 228838 58226
rect 228894 58170 228962 58226
rect 229018 58170 229088 58226
rect 228768 58102 229088 58170
rect 228768 58046 228838 58102
rect 228894 58046 228962 58102
rect 229018 58046 229088 58102
rect 228768 57978 229088 58046
rect 228768 57922 228838 57978
rect 228894 57922 228962 57978
rect 229018 57922 229088 57978
rect 228768 57888 229088 57922
rect 259488 58350 259808 58384
rect 259488 58294 259558 58350
rect 259614 58294 259682 58350
rect 259738 58294 259808 58350
rect 259488 58226 259808 58294
rect 259488 58170 259558 58226
rect 259614 58170 259682 58226
rect 259738 58170 259808 58226
rect 259488 58102 259808 58170
rect 259488 58046 259558 58102
rect 259614 58046 259682 58102
rect 259738 58046 259808 58102
rect 259488 57978 259808 58046
rect 259488 57922 259558 57978
rect 259614 57922 259682 57978
rect 259738 57922 259808 57978
rect 259488 57888 259808 57922
rect 66858 40350 67478 48914
rect 66858 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 67478 40350
rect 66858 40226 67478 40294
rect 66858 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 67478 40226
rect 66858 40102 67478 40170
rect 66858 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 67478 40102
rect 66858 39978 67478 40046
rect 66858 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 67478 39978
rect 66858 22350 67478 39922
rect 66858 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 67478 22350
rect 66858 22226 67478 22294
rect 66858 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 67478 22226
rect 66858 22102 67478 22170
rect 66858 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 67478 22102
rect 66858 21978 67478 22046
rect 66858 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 67478 21978
rect 57148 4978 57204 4988
rect 43596 4610 43652 4620
rect 55132 4798 55188 4808
rect 41020 4162 41076 4172
rect 55132 3444 55188 4742
rect 55132 3378 55188 3388
rect 57148 3444 57204 4922
rect 57148 3378 57204 3388
rect 66858 4350 67478 21922
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 46350 71198 48914
rect 70578 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 71198 46350
rect 70578 46226 71198 46294
rect 70578 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 71198 46226
rect 70578 46102 71198 46170
rect 70578 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 71198 46102
rect 70578 45978 71198 46046
rect 70578 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 71198 45978
rect 70578 28350 71198 45922
rect 90636 47818 90692 47828
rect 70578 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 71198 28350
rect 70578 28226 71198 28294
rect 70578 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 71198 28226
rect 70578 28102 71198 28170
rect 70578 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 71198 28102
rect 70578 27978 71198 28046
rect 70578 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 71198 27978
rect 70578 10350 71198 27922
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 70578 -1120 71198 9922
rect 75516 41158 75572 41168
rect 75516 4116 75572 41102
rect 75516 4050 75572 4060
rect 90636 4116 90692 47762
rect 90636 4050 90692 4060
rect 97578 40350 98198 48914
rect 97578 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 98198 40350
rect 97578 40226 98198 40294
rect 97578 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 98198 40226
rect 97578 40102 98198 40170
rect 97578 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 98198 40102
rect 97578 39978 98198 40046
rect 97578 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 98198 39978
rect 97578 22350 98198 39922
rect 97578 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 98198 22350
rect 97578 22226 98198 22294
rect 97578 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 98198 22226
rect 97578 22102 98198 22170
rect 97578 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 98198 22102
rect 97578 21978 98198 22046
rect 97578 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 98198 21978
rect 97578 4350 98198 21922
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 46350 101918 48914
rect 101298 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 101918 46350
rect 101298 46226 101918 46294
rect 101298 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 101918 46226
rect 101298 46102 101918 46170
rect 101298 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 101918 46102
rect 101298 45978 101918 46046
rect 101298 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 101918 45978
rect 101298 28350 101918 45922
rect 110796 47998 110852 48008
rect 101298 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 101918 28350
rect 101298 28226 101918 28294
rect 101298 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 101918 28226
rect 101298 28102 101918 28170
rect 101298 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 101918 28102
rect 101298 27978 101918 28046
rect 101298 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 101918 27978
rect 101298 10350 101918 27922
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 101298 -1120 101918 9922
rect 104076 44578 104132 44588
rect 104076 4228 104132 44522
rect 104076 4162 104132 4172
rect 110796 4228 110852 47942
rect 110796 4162 110852 4172
rect 128298 40350 128918 48914
rect 128298 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 128918 40350
rect 128298 40226 128918 40294
rect 128298 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 128918 40226
rect 128298 40102 128918 40170
rect 128298 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 128918 40102
rect 128298 39978 128918 40046
rect 128298 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 128918 39978
rect 128298 22350 128918 39922
rect 128298 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 128918 22350
rect 128298 22226 128918 22294
rect 128298 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 128918 22226
rect 128298 22102 128918 22170
rect 128298 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 128918 22102
rect 128298 21978 128918 22046
rect 128298 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 128918 21978
rect 128298 4350 128918 21922
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 46350 132638 48914
rect 132018 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 132638 46350
rect 132018 46226 132638 46294
rect 132018 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 132638 46226
rect 132018 46102 132638 46170
rect 132018 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 132638 46102
rect 132018 45978 132638 46046
rect 132018 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 132638 45978
rect 132018 28350 132638 45922
rect 132018 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 132638 28350
rect 132018 28226 132638 28294
rect 132018 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 132638 28226
rect 132018 28102 132638 28170
rect 132018 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 132638 28102
rect 132018 27978 132638 28046
rect 132018 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 132638 27978
rect 132018 10350 132638 27922
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 132018 -1120 132638 9922
rect 154476 44758 154532 44768
rect 137228 4978 137284 4988
rect 137228 3444 137284 4922
rect 137228 3378 137284 3388
rect 148652 4798 148708 4808
rect 148652 3444 148708 4742
rect 154476 4116 154532 44702
rect 154476 4050 154532 4060
rect 159018 40350 159638 48914
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 159018 22350 159638 39922
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 159018 4350 159638 21922
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 159018 4102 159638 4170
rect 148652 3378 148708 3388
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 46350 163358 48914
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 162738 28350 163358 45922
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 162738 10350 163358 27922
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 162738 -1120 163358 9922
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 40350 190358 48914
rect 189738 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 190358 40350
rect 189738 40226 190358 40294
rect 189738 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 190358 40226
rect 189738 40102 190358 40170
rect 189738 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 190358 40102
rect 189738 39978 190358 40046
rect 189738 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 190358 39978
rect 189738 22350 190358 39922
rect 189738 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 190358 22350
rect 189738 22226 190358 22294
rect 189738 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 190358 22226
rect 189738 22102 190358 22170
rect 189738 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 190358 22102
rect 189738 21978 190358 22046
rect 189738 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 190358 21978
rect 189738 4350 190358 21922
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 189738 4102 190358 4170
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 46350 194078 48914
rect 193458 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 194078 46350
rect 193458 46226 194078 46294
rect 193458 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 194078 46226
rect 193458 46102 194078 46170
rect 193458 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 194078 46102
rect 193458 45978 194078 46046
rect 193458 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 194078 45978
rect 193458 28350 194078 45922
rect 193458 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 194078 28350
rect 193458 28226 194078 28294
rect 193458 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 194078 28226
rect 193458 28102 194078 28170
rect 193458 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 194078 28102
rect 193458 27978 194078 28046
rect 193458 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 194078 27978
rect 193458 10350 194078 27922
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 193458 -1120 194078 9922
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 40350 221078 48914
rect 220458 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 221078 40350
rect 220458 40226 221078 40294
rect 220458 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 221078 40226
rect 220458 40102 221078 40170
rect 220458 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 221078 40102
rect 220458 39978 221078 40046
rect 220458 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 221078 39978
rect 220458 22350 221078 39922
rect 220458 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 221078 22350
rect 220458 22226 221078 22294
rect 220458 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 221078 22226
rect 220458 22102 221078 22170
rect 220458 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 221078 22102
rect 220458 21978 221078 22046
rect 220458 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 221078 21978
rect 220458 4350 221078 21922
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 46350 224798 48914
rect 224178 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 224798 46350
rect 224178 46226 224798 46294
rect 224178 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 224798 46226
rect 224178 46102 224798 46170
rect 224178 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 224798 46102
rect 224178 45978 224798 46046
rect 224178 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 224798 45978
rect 224178 28350 224798 45922
rect 224178 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 224798 28350
rect 224178 28226 224798 28294
rect 224178 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 224798 28226
rect 224178 28102 224798 28170
rect 224178 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 224798 28102
rect 224178 27978 224798 28046
rect 224178 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 224798 27978
rect 224178 10350 224798 27922
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 224178 -1120 224798 9922
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 40350 251798 48914
rect 251178 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 251798 40350
rect 251178 40226 251798 40294
rect 251178 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 251798 40226
rect 251178 40102 251798 40170
rect 251178 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 251798 40102
rect 251178 39978 251798 40046
rect 251178 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 251798 39978
rect 251178 22350 251798 39922
rect 251178 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 251798 22350
rect 251178 22226 251798 22294
rect 251178 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 251798 22226
rect 251178 22102 251798 22170
rect 251178 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 251798 22102
rect 251178 21978 251798 22046
rect 251178 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 251798 21978
rect 251178 4350 251798 21922
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 251178 4102 251798 4170
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 251178 -160 251798 3922
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 46350 255518 48914
rect 266924 48580 266980 234444
rect 267036 209098 267092 236908
rect 268604 236964 268660 236974
rect 267260 231812 267316 231822
rect 267036 209032 267092 209042
rect 267148 231058 267204 231068
rect 266924 48514 266980 48524
rect 254898 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 255518 46350
rect 254898 46226 255518 46294
rect 254898 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 255518 46226
rect 254898 46102 255518 46170
rect 254898 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 255518 46102
rect 254898 45978 255518 46046
rect 254898 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 255518 45978
rect 254898 28350 255518 45922
rect 254898 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 255518 28350
rect 254898 28226 255518 28294
rect 254898 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 255518 28226
rect 254898 28102 255518 28170
rect 254898 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 255518 28102
rect 254898 27978 255518 28046
rect 254898 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 255518 27978
rect 254898 10350 255518 27922
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 254898 -1120 255518 9922
rect 267148 4228 267204 231002
rect 267260 4340 267316 231756
rect 267484 231588 267540 231598
rect 267372 224578 267428 224588
rect 267372 38276 267428 224522
rect 267484 47998 267540 231532
rect 267484 47932 267540 47942
rect 267596 211438 267652 211448
rect 267596 47796 267652 211382
rect 268604 110098 268660 236908
rect 268604 110032 268660 110042
rect 268716 106678 268772 237020
rect 269500 231700 269556 231710
rect 269388 230916 269444 230926
rect 269164 211258 269220 211268
rect 269164 196588 269220 211202
rect 269276 209636 269332 209646
rect 269276 201236 269332 209580
rect 269276 201170 269332 201180
rect 269164 196532 269332 196588
rect 268716 106612 268772 106622
rect 269276 96404 269332 196532
rect 269276 96338 269332 96348
rect 269388 48132 269444 230860
rect 269388 48066 269444 48076
rect 269500 48020 269556 231644
rect 269500 47954 269556 47964
rect 269612 231476 269668 231486
rect 269612 47908 269668 231420
rect 269724 231238 269780 231248
rect 269724 49588 269780 231182
rect 269724 49522 269780 49532
rect 269612 47842 269668 47852
rect 267596 47730 267652 47740
rect 267372 38210 267428 38220
rect 269836 5908 269892 237122
rect 270060 234276 270116 234286
rect 269948 231418 270004 231428
rect 269948 44548 270004 231362
rect 270060 47818 270116 234220
rect 270060 47752 270116 47762
rect 269948 44482 270004 44492
rect 270508 29428 270564 238252
rect 270620 232932 270676 232942
rect 270620 41748 270676 232876
rect 271068 232820 271124 232830
rect 270732 227998 270788 228008
rect 270732 41972 270788 227942
rect 270732 41906 270788 41916
rect 270844 227818 270900 227828
rect 270620 41682 270676 41692
rect 270844 41636 270900 227762
rect 270956 227638 271012 227648
rect 270956 44660 271012 227582
rect 271068 49700 271124 232764
rect 272860 224980 272916 224990
rect 271180 219716 271236 219726
rect 271180 160468 271236 219660
rect 272524 218148 272580 218158
rect 272300 214900 272356 214910
rect 271292 211428 271348 211438
rect 271292 169204 271348 211372
rect 272188 211316 272244 211326
rect 272188 209636 272244 211260
rect 272188 209570 272244 209580
rect 272300 208348 272356 214844
rect 272412 212996 272468 213006
rect 272412 211316 272468 212940
rect 272412 211250 272468 211260
rect 272524 208348 272580 218092
rect 272636 216132 272692 216142
rect 272636 209524 272692 216076
rect 272636 209458 272692 209468
rect 272748 211092 272804 211102
rect 272300 208292 272468 208348
rect 272524 208292 272692 208348
rect 271292 169138 271348 169148
rect 272188 202468 272244 202478
rect 271180 160402 271236 160412
rect 272188 110964 272244 202412
rect 272412 186676 272468 208292
rect 272636 192500 272692 208292
rect 272748 204148 272804 211036
rect 272860 208348 272916 224924
rect 272972 209860 273028 239484
rect 273868 224218 273924 224228
rect 272972 209794 273028 209804
rect 273196 210532 273252 210542
rect 273084 209412 273140 209422
rect 272860 208292 273028 208348
rect 272748 204082 272804 204092
rect 272748 202580 272916 202618
rect 272748 202562 272860 202580
rect 272748 195412 272804 202562
rect 272860 202514 272916 202524
rect 272972 202258 273028 208292
rect 272748 195346 272804 195356
rect 272860 202202 273028 202258
rect 272636 192434 272692 192444
rect 272860 189588 272916 202202
rect 272860 189522 272916 189532
rect 272972 199892 273028 199902
rect 272412 186610 272468 186620
rect 272300 153658 272356 153674
rect 272300 153570 272356 153580
rect 272188 110898 272244 110908
rect 272972 108052 273028 199836
rect 273084 198324 273140 209356
rect 273196 202580 273252 210476
rect 273196 202514 273252 202524
rect 273420 209636 273476 209646
rect 273084 198258 273140 198268
rect 273420 183764 273476 209580
rect 273420 183698 273476 183708
rect 272972 107986 273028 107996
rect 271068 49634 271124 49644
rect 270956 44594 271012 44604
rect 270844 41570 270900 41580
rect 273868 37828 273924 224162
rect 273980 163380 274036 239596
rect 277228 236998 277284 237008
rect 275548 224398 275604 224408
rect 274428 221396 274484 221406
rect 274316 211204 274372 211214
rect 273980 163314 274036 163324
rect 274092 210178 274148 210188
rect 274092 154196 274148 210122
rect 274204 208738 274260 208748
rect 274204 154420 274260 208682
rect 274316 154644 274372 211148
rect 274428 172116 274484 221340
rect 274428 172050 274484 172060
rect 274652 216468 274708 216478
rect 274316 154578 274372 154588
rect 274204 154354 274260 154364
rect 274092 154130 274148 154140
rect 274652 153478 274708 216412
rect 274652 144564 274708 153422
rect 274652 144498 274708 144508
rect 275548 38164 275604 224342
rect 275548 38098 275604 38108
rect 276332 213108 276388 213118
rect 273868 37762 273924 37772
rect 270508 29362 270564 29372
rect 276332 7140 276388 213052
rect 277228 44772 277284 236942
rect 277340 212884 277396 212894
rect 277340 151732 277396 212828
rect 277340 151666 277396 151676
rect 277228 44706 277284 44716
rect 276332 7074 276388 7084
rect 269836 5842 269892 5852
rect 281372 4798 281428 239708
rect 281372 4732 281428 4742
rect 281898 238350 282518 240034
rect 281898 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 282518 238350
rect 281898 238226 282518 238294
rect 281898 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 282518 238226
rect 281898 238102 282518 238170
rect 281898 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 282518 238102
rect 281898 237978 282518 238046
rect 281898 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 282518 237978
rect 281898 220350 282518 237922
rect 281898 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 282518 220350
rect 281898 220226 282518 220294
rect 281898 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 282518 220226
rect 281898 220102 282518 220170
rect 281898 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 282518 220102
rect 281898 219978 282518 220046
rect 281898 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 282518 219978
rect 281898 202350 282518 219922
rect 281898 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 282518 202350
rect 281898 202226 282518 202294
rect 281898 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 282518 202226
rect 281898 202102 282518 202170
rect 281898 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 282518 202102
rect 281898 201978 282518 202046
rect 281898 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 282518 201978
rect 281898 184350 282518 201922
rect 281898 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 282518 184350
rect 281898 184226 282518 184294
rect 281898 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 282518 184226
rect 281898 184102 282518 184170
rect 281898 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 282518 184102
rect 281898 183978 282518 184046
rect 281898 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 282518 183978
rect 281898 166350 282518 183922
rect 281898 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 282518 166350
rect 281898 166226 282518 166294
rect 281898 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 282518 166226
rect 281898 166102 282518 166170
rect 281898 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 282518 166102
rect 281898 165978 282518 166046
rect 281898 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 282518 165978
rect 281898 148350 282518 165922
rect 281898 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 282518 148350
rect 281898 148226 282518 148294
rect 281898 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 282518 148226
rect 281898 148102 282518 148170
rect 281898 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 282518 148102
rect 281898 147978 282518 148046
rect 281898 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 282518 147978
rect 281898 130350 282518 147922
rect 281898 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 282518 130350
rect 281898 130226 282518 130294
rect 281898 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 282518 130226
rect 281898 130102 282518 130170
rect 281898 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 282518 130102
rect 281898 129978 282518 130046
rect 281898 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 282518 129978
rect 281898 112350 282518 129922
rect 281898 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 282518 112350
rect 281898 112226 282518 112294
rect 281898 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 282518 112226
rect 281898 112102 282518 112170
rect 281898 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 282518 112102
rect 281898 111978 282518 112046
rect 281898 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 282518 111978
rect 281898 94350 282518 111922
rect 281898 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 282518 94350
rect 281898 94226 282518 94294
rect 281898 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 282518 94226
rect 281898 94102 282518 94170
rect 281898 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 282518 94102
rect 281898 93978 282518 94046
rect 281898 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 282518 93978
rect 281898 76350 282518 93922
rect 281898 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 282518 76350
rect 281898 76226 282518 76294
rect 281898 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 282518 76226
rect 281898 76102 282518 76170
rect 281898 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 282518 76102
rect 281898 75978 282518 76046
rect 281898 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 282518 75978
rect 281898 58350 282518 75922
rect 281898 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 282518 58350
rect 281898 58226 282518 58294
rect 281898 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 282518 58226
rect 281898 58102 282518 58170
rect 281898 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 282518 58102
rect 281898 57978 282518 58046
rect 281898 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 282518 57978
rect 281898 40350 282518 57922
rect 283052 234612 283108 234622
rect 283052 44758 283108 234556
rect 283052 44692 283108 44702
rect 285618 226350 286238 240034
rect 285618 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 286238 226350
rect 285618 226226 286238 226294
rect 285618 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 286238 226226
rect 285618 226102 286238 226170
rect 285618 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 286238 226102
rect 285618 225978 286238 226046
rect 285618 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 286238 225978
rect 285618 208350 286238 225922
rect 285618 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 286238 208350
rect 285618 208226 286238 208294
rect 285618 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 286238 208226
rect 285618 208102 286238 208170
rect 285618 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 286238 208102
rect 285618 207978 286238 208046
rect 285618 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 286238 207978
rect 285618 190350 286238 207922
rect 285618 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 286238 190350
rect 285618 190226 286238 190294
rect 285618 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 286238 190226
rect 285618 190102 286238 190170
rect 285618 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 286238 190102
rect 285618 189978 286238 190046
rect 285618 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 286238 189978
rect 285618 172350 286238 189922
rect 285618 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 286238 172350
rect 285618 172226 286238 172294
rect 285618 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 286238 172226
rect 285618 172102 286238 172170
rect 285618 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 286238 172102
rect 285618 171978 286238 172046
rect 285618 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 286238 171978
rect 285618 154350 286238 171922
rect 285618 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 286238 154350
rect 285618 154226 286238 154294
rect 285618 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 286238 154226
rect 285618 154102 286238 154170
rect 285618 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 286238 154102
rect 285618 153978 286238 154046
rect 285618 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 286238 153978
rect 285618 136350 286238 153922
rect 285618 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 286238 136350
rect 285618 136226 286238 136294
rect 285618 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 286238 136226
rect 285618 136102 286238 136170
rect 285618 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 286238 136102
rect 285618 135978 286238 136046
rect 285618 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 286238 135978
rect 285618 118350 286238 135922
rect 285618 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 286238 118350
rect 285618 118226 286238 118294
rect 285618 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 286238 118226
rect 285618 118102 286238 118170
rect 285618 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 286238 118102
rect 285618 117978 286238 118046
rect 285618 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 286238 117978
rect 285618 100350 286238 117922
rect 285618 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 286238 100350
rect 285618 100226 286238 100294
rect 285618 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 286238 100226
rect 285618 100102 286238 100170
rect 285618 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 286238 100102
rect 285618 99978 286238 100046
rect 285618 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 286238 99978
rect 285618 82350 286238 99922
rect 285618 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 286238 82350
rect 285618 82226 286238 82294
rect 285618 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 286238 82226
rect 285618 82102 286238 82170
rect 285618 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 286238 82102
rect 285618 81978 286238 82046
rect 285618 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 286238 81978
rect 285618 64350 286238 81922
rect 285618 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 286238 64350
rect 285618 64226 286238 64294
rect 285618 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 286238 64226
rect 285618 64102 286238 64170
rect 285618 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 286238 64102
rect 285618 63978 286238 64046
rect 285618 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 286238 63978
rect 285618 46350 286238 63922
rect 285618 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 286238 46350
rect 285618 46226 286238 46294
rect 285618 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 286238 46226
rect 285618 46102 286238 46170
rect 285618 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 286238 46102
rect 285618 45978 286238 46046
rect 285618 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 286238 45978
rect 281898 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 282518 40350
rect 281898 40226 282518 40294
rect 281898 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 282518 40226
rect 281898 40102 282518 40170
rect 281898 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 282518 40102
rect 281898 39978 282518 40046
rect 281898 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 282518 39978
rect 281898 22350 282518 39922
rect 281898 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 282518 22350
rect 281898 22226 282518 22294
rect 281898 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 282518 22226
rect 281898 22102 282518 22170
rect 281898 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 282518 22102
rect 281898 21978 282518 22046
rect 281898 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 282518 21978
rect 267260 4274 267316 4284
rect 281898 4350 282518 21922
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 267148 4162 267204 4172
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 285618 28350 286238 45922
rect 285618 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 286238 28350
rect 285618 28226 286238 28294
rect 285618 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 286238 28226
rect 285618 28102 286238 28170
rect 285618 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 286238 28102
rect 285618 27978 286238 28046
rect 285618 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 286238 27978
rect 285618 10350 286238 27922
rect 285618 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 286238 10350
rect 285618 10226 286238 10294
rect 285618 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 286238 10226
rect 285618 10102 286238 10170
rect 285618 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 286238 10102
rect 285618 9978 286238 10046
rect 285618 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 286238 9978
rect 285618 -1120 286238 9922
rect 288316 239092 288372 239102
rect 288316 4978 288372 239036
rect 288316 4912 288372 4922
rect 289772 4564 289828 241082
rect 312618 238350 313238 240034
rect 312618 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 313238 238350
rect 312618 238226 313238 238294
rect 312618 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 313238 238226
rect 312618 238102 313238 238170
rect 312618 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 313238 238102
rect 312618 237978 313238 238046
rect 312618 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 313238 237978
rect 302316 236964 302372 236974
rect 296604 223076 296660 223086
rect 296492 210756 296548 210766
rect 293132 209076 293188 209086
rect 293132 104158 293188 209020
rect 293244 141958 293300 141968
rect 293244 125524 293300 141902
rect 293244 125458 293300 125468
rect 293132 104092 293188 104102
rect 296492 103978 296548 210700
rect 296604 152758 296660 223020
rect 301532 222740 301588 222750
rect 296604 152692 296660 152702
rect 298172 209098 298228 209108
rect 298172 106820 298228 209042
rect 300636 199332 300692 199342
rect 298956 198100 299012 198110
rect 298956 157438 299012 198044
rect 300524 195972 300580 195982
rect 300524 160468 300580 195916
rect 300636 160580 300692 199276
rect 300636 160514 300692 160524
rect 300524 160402 300580 160412
rect 298956 157372 299012 157382
rect 298172 106754 298228 106764
rect 296492 103912 296548 103922
rect 301532 99988 301588 222684
rect 301644 219940 301700 219950
rect 301644 142772 301700 219884
rect 302316 159124 302372 236908
rect 302316 159058 302372 159068
rect 303436 236964 303492 236974
rect 303436 152068 303492 236908
rect 307356 236964 307412 236974
rect 305468 184350 305788 184384
rect 305468 184294 305538 184350
rect 305594 184294 305662 184350
rect 305718 184294 305788 184350
rect 305468 184226 305788 184294
rect 305468 184170 305538 184226
rect 305594 184170 305662 184226
rect 305718 184170 305788 184226
rect 305468 184102 305788 184170
rect 305468 184046 305538 184102
rect 305594 184046 305662 184102
rect 305718 184046 305788 184102
rect 305468 183978 305788 184046
rect 305468 183922 305538 183978
rect 305594 183922 305662 183978
rect 305718 183922 305788 183978
rect 305468 183888 305788 183922
rect 305468 166350 305788 166384
rect 305468 166294 305538 166350
rect 305594 166294 305662 166350
rect 305718 166294 305788 166350
rect 305468 166226 305788 166294
rect 305468 166170 305538 166226
rect 305594 166170 305662 166226
rect 305718 166170 305788 166226
rect 305468 166102 305788 166170
rect 305468 166046 305538 166102
rect 305594 166046 305662 166102
rect 305718 166046 305788 166102
rect 305468 165978 305788 166046
rect 305468 165922 305538 165978
rect 305594 165922 305662 165978
rect 305718 165922 305788 165978
rect 305468 165888 305788 165922
rect 303996 160804 304052 160814
rect 303996 160468 304052 160748
rect 307356 160580 307412 236908
rect 309036 236964 309092 236974
rect 309036 197578 309092 236908
rect 309036 197512 309092 197522
rect 310716 236964 310772 236974
rect 310716 197398 310772 236908
rect 310716 197332 310772 197342
rect 312618 220350 313238 237922
rect 312618 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 313238 220350
rect 312618 220226 313238 220294
rect 312618 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 313238 220226
rect 312618 220102 313238 220170
rect 312618 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 313238 220102
rect 312618 219978 313238 220046
rect 312618 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 313238 219978
rect 312618 202350 313238 219922
rect 312618 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 313238 202350
rect 312618 202226 313238 202294
rect 312618 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 313238 202226
rect 312618 202102 313238 202170
rect 312618 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 313238 202102
rect 312618 201978 313238 202046
rect 312618 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 313238 201978
rect 312618 193230 313238 201922
rect 316338 226350 316958 240034
rect 336812 238618 336868 238628
rect 316338 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 316958 226350
rect 316338 226226 316958 226294
rect 316338 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 316958 226226
rect 316338 226102 316958 226170
rect 316338 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 316958 226102
rect 316338 225978 316958 226046
rect 316338 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 316958 225978
rect 316338 208350 316958 225922
rect 316338 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 316958 208350
rect 316338 208226 316958 208294
rect 316338 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 316958 208226
rect 316338 208102 316958 208170
rect 316338 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 316958 208102
rect 316338 207978 316958 208046
rect 316338 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 316958 207978
rect 316338 193230 316958 207922
rect 319116 236964 319172 236974
rect 318556 197204 318612 197214
rect 318556 195860 318612 197148
rect 318556 195794 318612 195804
rect 319116 193978 319172 236908
rect 334236 236964 334292 236974
rect 325276 197204 325332 197214
rect 323820 196532 323876 196542
rect 323820 196308 323876 196476
rect 323820 196242 323876 196252
rect 325276 195748 325332 197148
rect 325276 195682 325332 195692
rect 319116 193912 319172 193922
rect 334236 192358 334292 236908
rect 335916 236964 335972 236974
rect 335916 193258 335972 236908
rect 335916 193202 336084 193258
rect 336028 192538 336084 193202
rect 336028 192500 336420 192538
rect 336028 192482 336364 192500
rect 336364 192434 336420 192444
rect 334236 192292 334292 192302
rect 309752 190350 310072 190384
rect 309752 190294 309822 190350
rect 309878 190294 309946 190350
rect 310002 190294 310072 190350
rect 309752 190226 310072 190294
rect 309752 190170 309822 190226
rect 309878 190170 309946 190226
rect 310002 190170 310072 190226
rect 309752 190102 310072 190170
rect 309752 190046 309822 190102
rect 309878 190046 309946 190102
rect 310002 190046 310072 190102
rect 309752 189978 310072 190046
rect 309752 189922 309822 189978
rect 309878 189922 309946 189978
rect 310002 189922 310072 189978
rect 309752 189888 310072 189922
rect 318320 190350 318640 190384
rect 318320 190294 318390 190350
rect 318446 190294 318514 190350
rect 318570 190294 318640 190350
rect 318320 190226 318640 190294
rect 318320 190170 318390 190226
rect 318446 190170 318514 190226
rect 318570 190170 318640 190226
rect 318320 190102 318640 190170
rect 318320 190046 318390 190102
rect 318446 190046 318514 190102
rect 318570 190046 318640 190102
rect 318320 189978 318640 190046
rect 318320 189922 318390 189978
rect 318446 189922 318514 189978
rect 318570 189922 318640 189978
rect 318320 189888 318640 189922
rect 326888 190350 327208 190384
rect 326888 190294 326958 190350
rect 327014 190294 327082 190350
rect 327138 190294 327208 190350
rect 326888 190226 327208 190294
rect 326888 190170 326958 190226
rect 327014 190170 327082 190226
rect 327138 190170 327208 190226
rect 326888 190102 327208 190170
rect 326888 190046 326958 190102
rect 327014 190046 327082 190102
rect 327138 190046 327208 190102
rect 326888 189978 327208 190046
rect 326888 189922 326958 189978
rect 327014 189922 327082 189978
rect 327138 189922 327208 189978
rect 326888 189888 327208 189922
rect 335456 190350 335776 190384
rect 335456 190294 335526 190350
rect 335582 190294 335650 190350
rect 335706 190294 335776 190350
rect 335456 190226 335776 190294
rect 335456 190170 335526 190226
rect 335582 190170 335650 190226
rect 335706 190170 335776 190226
rect 335456 190102 335776 190170
rect 335456 190046 335526 190102
rect 335582 190046 335650 190102
rect 335706 190046 335776 190102
rect 335456 189978 335776 190046
rect 335456 189922 335526 189978
rect 335582 189922 335650 189978
rect 335706 189922 335776 189978
rect 335456 189888 335776 189922
rect 314036 184350 314356 184384
rect 314036 184294 314106 184350
rect 314162 184294 314230 184350
rect 314286 184294 314356 184350
rect 314036 184226 314356 184294
rect 314036 184170 314106 184226
rect 314162 184170 314230 184226
rect 314286 184170 314356 184226
rect 314036 184102 314356 184170
rect 314036 184046 314106 184102
rect 314162 184046 314230 184102
rect 314286 184046 314356 184102
rect 314036 183978 314356 184046
rect 314036 183922 314106 183978
rect 314162 183922 314230 183978
rect 314286 183922 314356 183978
rect 314036 183888 314356 183922
rect 322604 184350 322924 184384
rect 322604 184294 322674 184350
rect 322730 184294 322798 184350
rect 322854 184294 322924 184350
rect 322604 184226 322924 184294
rect 322604 184170 322674 184226
rect 322730 184170 322798 184226
rect 322854 184170 322924 184226
rect 322604 184102 322924 184170
rect 322604 184046 322674 184102
rect 322730 184046 322798 184102
rect 322854 184046 322924 184102
rect 322604 183978 322924 184046
rect 322604 183922 322674 183978
rect 322730 183922 322798 183978
rect 322854 183922 322924 183978
rect 322604 183888 322924 183922
rect 331172 184350 331492 184384
rect 331172 184294 331242 184350
rect 331298 184294 331366 184350
rect 331422 184294 331492 184350
rect 331172 184226 331492 184294
rect 331172 184170 331242 184226
rect 331298 184170 331366 184226
rect 331422 184170 331492 184226
rect 331172 184102 331492 184170
rect 331172 184046 331242 184102
rect 331298 184046 331366 184102
rect 331422 184046 331492 184102
rect 331172 183978 331492 184046
rect 331172 183922 331242 183978
rect 331298 183922 331366 183978
rect 331422 183922 331492 183978
rect 331172 183888 331492 183922
rect 309752 172350 310072 172384
rect 309752 172294 309822 172350
rect 309878 172294 309946 172350
rect 310002 172294 310072 172350
rect 309752 172226 310072 172294
rect 309752 172170 309822 172226
rect 309878 172170 309946 172226
rect 310002 172170 310072 172226
rect 309752 172102 310072 172170
rect 309752 172046 309822 172102
rect 309878 172046 309946 172102
rect 310002 172046 310072 172102
rect 309752 171978 310072 172046
rect 309752 171922 309822 171978
rect 309878 171922 309946 171978
rect 310002 171922 310072 171978
rect 309752 171888 310072 171922
rect 318320 172350 318640 172384
rect 318320 172294 318390 172350
rect 318446 172294 318514 172350
rect 318570 172294 318640 172350
rect 318320 172226 318640 172294
rect 318320 172170 318390 172226
rect 318446 172170 318514 172226
rect 318570 172170 318640 172226
rect 318320 172102 318640 172170
rect 318320 172046 318390 172102
rect 318446 172046 318514 172102
rect 318570 172046 318640 172102
rect 318320 171978 318640 172046
rect 318320 171922 318390 171978
rect 318446 171922 318514 171978
rect 318570 171922 318640 171978
rect 318320 171888 318640 171922
rect 326888 172350 327208 172384
rect 326888 172294 326958 172350
rect 327014 172294 327082 172350
rect 327138 172294 327208 172350
rect 326888 172226 327208 172294
rect 326888 172170 326958 172226
rect 327014 172170 327082 172226
rect 327138 172170 327208 172226
rect 326888 172102 327208 172170
rect 326888 172046 326958 172102
rect 327014 172046 327082 172102
rect 327138 172046 327208 172102
rect 326888 171978 327208 172046
rect 326888 171922 326958 171978
rect 327014 171922 327082 171978
rect 327138 171922 327208 171978
rect 326888 171888 327208 171922
rect 335456 172350 335776 172384
rect 335456 172294 335526 172350
rect 335582 172294 335650 172350
rect 335706 172294 335776 172350
rect 335456 172226 335776 172294
rect 335456 172170 335526 172226
rect 335582 172170 335650 172226
rect 335706 172170 335776 172226
rect 335456 172102 335776 172170
rect 335456 172046 335526 172102
rect 335582 172046 335650 172102
rect 335706 172046 335776 172102
rect 335456 171978 335776 172046
rect 335456 171922 335526 171978
rect 335582 171922 335650 171978
rect 335706 171922 335776 171978
rect 335456 171888 335776 171922
rect 314036 166350 314356 166384
rect 314036 166294 314106 166350
rect 314162 166294 314230 166350
rect 314286 166294 314356 166350
rect 314036 166226 314356 166294
rect 314036 166170 314106 166226
rect 314162 166170 314230 166226
rect 314286 166170 314356 166226
rect 314036 166102 314356 166170
rect 314036 166046 314106 166102
rect 314162 166046 314230 166102
rect 314286 166046 314356 166102
rect 314036 165978 314356 166046
rect 314036 165922 314106 165978
rect 314162 165922 314230 165978
rect 314286 165922 314356 165978
rect 314036 165888 314356 165922
rect 322604 166350 322924 166384
rect 322604 166294 322674 166350
rect 322730 166294 322798 166350
rect 322854 166294 322924 166350
rect 322604 166226 322924 166294
rect 322604 166170 322674 166226
rect 322730 166170 322798 166226
rect 322854 166170 322924 166226
rect 322604 166102 322924 166170
rect 322604 166046 322674 166102
rect 322730 166046 322798 166102
rect 322854 166046 322924 166102
rect 322604 165978 322924 166046
rect 322604 165922 322674 165978
rect 322730 165922 322798 165978
rect 322854 165922 322924 165978
rect 322604 165888 322924 165922
rect 331172 166350 331492 166384
rect 331172 166294 331242 166350
rect 331298 166294 331366 166350
rect 331422 166294 331492 166350
rect 331172 166226 331492 166294
rect 331172 166170 331242 166226
rect 331298 166170 331366 166226
rect 331422 166170 331492 166226
rect 331172 166102 331492 166170
rect 331172 166046 331242 166102
rect 331298 166046 331366 166102
rect 331422 166046 331492 166102
rect 331172 165978 331492 166046
rect 331172 165922 331242 165978
rect 331298 165922 331366 165978
rect 331422 165922 331492 165978
rect 331172 165888 331492 165922
rect 307356 160514 307412 160524
rect 303996 160402 304052 160412
rect 306572 157892 306628 157902
rect 306572 157438 306628 157836
rect 306572 157372 306628 157382
rect 303436 152002 303492 152012
rect 312618 148350 313238 163170
rect 312618 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 313238 148350
rect 312618 148226 313238 148294
rect 312618 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 313238 148226
rect 312618 148102 313238 148170
rect 312618 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 313238 148102
rect 312618 147978 313238 148046
rect 312618 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 313238 147978
rect 301644 142706 301700 142716
rect 311612 146998 311668 147008
rect 311612 119700 311668 146942
rect 311612 119634 311668 119644
rect 312618 130350 313238 147922
rect 312618 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 313238 130350
rect 312618 130226 313238 130294
rect 312618 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 313238 130226
rect 312618 130102 313238 130170
rect 312618 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 313238 130102
rect 312618 129978 313238 130046
rect 312618 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 313238 129978
rect 301532 99922 301588 99932
rect 312618 112350 313238 129922
rect 312618 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 313238 112350
rect 312618 112226 313238 112294
rect 312618 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 313238 112226
rect 312618 112102 313238 112170
rect 312618 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 313238 112102
rect 312618 111978 313238 112046
rect 312618 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 313238 111978
rect 312618 94350 313238 111922
rect 312618 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 313238 94350
rect 312618 94226 313238 94294
rect 312618 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 313238 94226
rect 312618 94102 313238 94170
rect 312618 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 313238 94102
rect 312618 93978 313238 94046
rect 312618 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 313238 93978
rect 299500 82147 299820 82204
rect 299500 82091 299528 82147
rect 299584 82091 299632 82147
rect 299688 82091 299736 82147
rect 299792 82091 299820 82147
rect 299500 82043 299820 82091
rect 299500 81987 299528 82043
rect 299584 81987 299632 82043
rect 299688 81987 299736 82043
rect 299792 81987 299820 82043
rect 299500 81939 299820 81987
rect 299500 81883 299528 81939
rect 299584 81883 299632 81939
rect 299688 81883 299736 81939
rect 299792 81883 299820 81939
rect 299500 81826 299820 81883
rect 307816 82147 308136 82204
rect 307816 82091 307844 82147
rect 307900 82091 307948 82147
rect 308004 82091 308052 82147
rect 308108 82091 308136 82147
rect 307816 82043 308136 82091
rect 307816 81987 307844 82043
rect 307900 81987 307948 82043
rect 308004 81987 308052 82043
rect 308108 81987 308136 82043
rect 307816 81939 308136 81987
rect 307816 81883 307844 81939
rect 307900 81883 307948 81939
rect 308004 81883 308052 81939
rect 308108 81883 308136 81939
rect 307816 81826 308136 81883
rect 295342 76350 295662 76384
rect 295342 76294 295412 76350
rect 295468 76294 295536 76350
rect 295592 76294 295662 76350
rect 295342 76226 295662 76294
rect 295342 76170 295412 76226
rect 295468 76170 295536 76226
rect 295592 76170 295662 76226
rect 295342 76102 295662 76170
rect 295342 76046 295412 76102
rect 295468 76046 295536 76102
rect 295592 76046 295662 76102
rect 295342 75978 295662 76046
rect 295342 75922 295412 75978
rect 295468 75922 295536 75978
rect 295592 75922 295662 75978
rect 295342 75888 295662 75922
rect 303658 76350 303978 76384
rect 303658 76294 303728 76350
rect 303784 76294 303852 76350
rect 303908 76294 303978 76350
rect 303658 76226 303978 76294
rect 303658 76170 303728 76226
rect 303784 76170 303852 76226
rect 303908 76170 303978 76226
rect 303658 76102 303978 76170
rect 303658 76046 303728 76102
rect 303784 76046 303852 76102
rect 303908 76046 303978 76102
rect 303658 75978 303978 76046
rect 303658 75922 303728 75978
rect 303784 75922 303852 75978
rect 303908 75922 303978 75978
rect 303658 75888 303978 75922
rect 311974 76350 312294 76384
rect 311974 76294 312044 76350
rect 312100 76294 312168 76350
rect 312224 76294 312294 76350
rect 311974 76226 312294 76294
rect 311974 76170 312044 76226
rect 312100 76170 312168 76226
rect 312224 76170 312294 76226
rect 311974 76102 312294 76170
rect 311974 76046 312044 76102
rect 312100 76046 312168 76102
rect 312224 76046 312294 76102
rect 311974 75978 312294 76046
rect 311974 75922 312044 75978
rect 312100 75922 312168 75978
rect 312224 75922 312294 75978
rect 311974 75888 312294 75922
rect 312618 76350 313238 93922
rect 316338 154350 316958 163170
rect 316338 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 316958 154350
rect 316338 154226 316958 154294
rect 316338 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 316958 154226
rect 316338 154102 316958 154170
rect 316338 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 316958 154102
rect 316338 153978 316958 154046
rect 316338 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 316958 153978
rect 316338 136350 316958 153922
rect 316338 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 316958 136350
rect 316338 136226 316958 136294
rect 316338 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 316958 136226
rect 316338 136102 316958 136170
rect 316338 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 316958 136102
rect 316338 135978 316958 136046
rect 316338 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 316958 135978
rect 316338 118350 316958 135922
rect 316338 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 316958 118350
rect 316338 118226 316958 118294
rect 316338 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 316958 118226
rect 316338 118102 316958 118170
rect 316338 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 316958 118102
rect 316338 117978 316958 118046
rect 316338 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 316958 117978
rect 316338 100350 316958 117922
rect 316338 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 316958 100350
rect 316338 100226 316958 100294
rect 316338 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 316958 100226
rect 316338 100102 316958 100170
rect 316338 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 316958 100102
rect 316338 99978 316958 100046
rect 316338 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 316958 99978
rect 316338 84316 316958 99922
rect 316132 82147 316452 82204
rect 316132 82091 316160 82147
rect 316216 82091 316264 82147
rect 316320 82091 316368 82147
rect 316424 82091 316452 82147
rect 316132 82043 316452 82091
rect 316132 81987 316160 82043
rect 316216 81987 316264 82043
rect 316320 81987 316368 82043
rect 316424 81987 316452 82043
rect 316132 81939 316452 81987
rect 316132 81883 316160 81939
rect 316216 81883 316264 81939
rect 316320 81883 316368 81939
rect 316424 81883 316452 81939
rect 316132 81826 316452 81883
rect 324448 82147 324768 82204
rect 324448 82091 324476 82147
rect 324532 82091 324580 82147
rect 324636 82091 324684 82147
rect 324740 82091 324768 82147
rect 324448 82043 324768 82091
rect 324448 81987 324476 82043
rect 324532 81987 324580 82043
rect 324636 81987 324684 82043
rect 324740 81987 324768 82043
rect 324448 81939 324768 81987
rect 324448 81883 324476 81939
rect 324532 81883 324580 81939
rect 324636 81883 324684 81939
rect 324740 81883 324768 81939
rect 324448 81826 324768 81883
rect 312618 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 313238 76350
rect 312618 76226 313238 76294
rect 312618 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 313238 76226
rect 312618 76102 313238 76170
rect 312618 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 313238 76102
rect 312618 75978 313238 76046
rect 312618 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 313238 75978
rect 299500 64350 299820 64384
rect 299500 64294 299570 64350
rect 299626 64294 299694 64350
rect 299750 64294 299820 64350
rect 299500 64226 299820 64294
rect 299500 64170 299570 64226
rect 299626 64170 299694 64226
rect 299750 64170 299820 64226
rect 299500 64102 299820 64170
rect 299500 64046 299570 64102
rect 299626 64046 299694 64102
rect 299750 64046 299820 64102
rect 299500 63978 299820 64046
rect 299500 63922 299570 63978
rect 299626 63922 299694 63978
rect 299750 63922 299820 63978
rect 299500 63888 299820 63922
rect 307816 64350 308136 64384
rect 307816 64294 307886 64350
rect 307942 64294 308010 64350
rect 308066 64294 308136 64350
rect 307816 64226 308136 64294
rect 307816 64170 307886 64226
rect 307942 64170 308010 64226
rect 308066 64170 308136 64226
rect 307816 64102 308136 64170
rect 307816 64046 307886 64102
rect 307942 64046 308010 64102
rect 308066 64046 308136 64102
rect 307816 63978 308136 64046
rect 307816 63922 307886 63978
rect 307942 63922 308010 63978
rect 308066 63922 308136 63978
rect 307816 63888 308136 63922
rect 295342 58350 295662 58384
rect 295342 58294 295412 58350
rect 295468 58294 295536 58350
rect 295592 58294 295662 58350
rect 295342 58226 295662 58294
rect 295342 58170 295412 58226
rect 295468 58170 295536 58226
rect 295592 58170 295662 58226
rect 295342 58102 295662 58170
rect 295342 58046 295412 58102
rect 295468 58046 295536 58102
rect 295592 58046 295662 58102
rect 295342 57978 295662 58046
rect 295342 57922 295412 57978
rect 295468 57922 295536 57978
rect 295592 57922 295662 57978
rect 295342 57888 295662 57922
rect 303658 58350 303978 58384
rect 303658 58294 303728 58350
rect 303784 58294 303852 58350
rect 303908 58294 303978 58350
rect 303658 58226 303978 58294
rect 303658 58170 303728 58226
rect 303784 58170 303852 58226
rect 303908 58170 303978 58226
rect 303658 58102 303978 58170
rect 303658 58046 303728 58102
rect 303784 58046 303852 58102
rect 303908 58046 303978 58102
rect 303658 57978 303978 58046
rect 303658 57922 303728 57978
rect 303784 57922 303852 57978
rect 303908 57922 303978 57978
rect 303658 57888 303978 57922
rect 311974 58350 312294 58384
rect 311974 58294 312044 58350
rect 312100 58294 312168 58350
rect 312224 58294 312294 58350
rect 311974 58226 312294 58294
rect 311974 58170 312044 58226
rect 312100 58170 312168 58226
rect 312224 58170 312294 58226
rect 311974 58102 312294 58170
rect 311974 58046 312044 58102
rect 312100 58046 312168 58102
rect 312224 58046 312294 58102
rect 311974 57978 312294 58046
rect 311974 57922 312044 57978
rect 312100 57922 312168 57978
rect 312224 57922 312294 57978
rect 311974 57888 312294 57922
rect 312618 58350 313238 75922
rect 320290 76350 320610 76384
rect 320290 76294 320360 76350
rect 320416 76294 320484 76350
rect 320540 76294 320610 76350
rect 320290 76226 320610 76294
rect 320290 76170 320360 76226
rect 320416 76170 320484 76226
rect 320540 76170 320610 76226
rect 320290 76102 320610 76170
rect 320290 76046 320360 76102
rect 320416 76046 320484 76102
rect 320540 76046 320610 76102
rect 320290 75978 320610 76046
rect 320290 75922 320360 75978
rect 320416 75922 320484 75978
rect 320540 75922 320610 75978
rect 320290 75888 320610 75922
rect 316132 64350 316452 64384
rect 316132 64294 316202 64350
rect 316258 64294 316326 64350
rect 316382 64294 316452 64350
rect 316132 64226 316452 64294
rect 316132 64170 316202 64226
rect 316258 64170 316326 64226
rect 316382 64170 316452 64226
rect 316132 64102 316452 64170
rect 316132 64046 316202 64102
rect 316258 64046 316326 64102
rect 316382 64046 316452 64102
rect 316132 63978 316452 64046
rect 316132 63922 316202 63978
rect 316258 63922 316326 63978
rect 316382 63922 316452 63978
rect 316132 63888 316452 63922
rect 324448 64350 324768 64384
rect 324448 64294 324518 64350
rect 324574 64294 324642 64350
rect 324698 64294 324768 64350
rect 324448 64226 324768 64294
rect 324448 64170 324518 64226
rect 324574 64170 324642 64226
rect 324698 64170 324768 64226
rect 324448 64102 324768 64170
rect 324448 64046 324518 64102
rect 324574 64046 324642 64102
rect 324698 64046 324768 64102
rect 324448 63978 324768 64046
rect 324448 63922 324518 63978
rect 324574 63922 324642 63978
rect 324698 63922 324768 63978
rect 324448 63888 324768 63922
rect 312618 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 313238 58350
rect 312618 58226 313238 58294
rect 312618 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 313238 58226
rect 312618 58102 313238 58170
rect 312618 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 313238 58102
rect 312618 57978 313238 58046
rect 312618 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 313238 57978
rect 289772 4498 289828 4508
rect 312618 40350 313238 57922
rect 320290 58350 320610 58384
rect 320290 58294 320360 58350
rect 320416 58294 320484 58350
rect 320540 58294 320610 58350
rect 320290 58226 320610 58294
rect 320290 58170 320360 58226
rect 320416 58170 320484 58226
rect 320540 58170 320610 58226
rect 320290 58102 320610 58170
rect 320290 58046 320360 58102
rect 320416 58046 320484 58102
rect 320540 58046 320610 58102
rect 320290 57978 320610 58046
rect 320290 57922 320360 57978
rect 320416 57922 320484 57978
rect 320540 57922 320610 57978
rect 320290 57888 320610 57922
rect 312618 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 313238 40350
rect 312618 40226 313238 40294
rect 312618 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 313238 40226
rect 312618 40102 313238 40170
rect 312618 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 313238 40102
rect 312618 39978 313238 40046
rect 312618 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 313238 39978
rect 312618 22350 313238 39922
rect 312618 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 313238 22350
rect 312618 22226 313238 22294
rect 312618 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 313238 22226
rect 312618 22102 313238 22170
rect 312618 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 313238 22102
rect 312618 21978 313238 22046
rect 312618 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 313238 21978
rect 285618 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 286238 -1120
rect 285618 -1244 286238 -1176
rect 285618 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 286238 -1244
rect 285618 -1368 286238 -1300
rect 285618 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 286238 -1368
rect 285618 -1492 286238 -1424
rect 285618 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 286238 -1492
rect 285618 -1644 286238 -1548
rect 312618 4350 313238 21922
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 316338 46350 316958 50964
rect 316338 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 316958 46350
rect 316338 46226 316958 46294
rect 316338 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 316958 46226
rect 316338 46102 316958 46170
rect 316338 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 316958 46102
rect 316338 45978 316958 46046
rect 316338 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 316958 45978
rect 316338 28350 316958 45922
rect 336812 41860 336868 238562
rect 336924 46228 336980 241442
rect 337260 241318 337316 241328
rect 337148 240238 337204 240248
rect 337036 219268 337092 219278
rect 337036 164638 337092 219212
rect 337036 164572 337092 164582
rect 337148 46452 337204 240182
rect 337260 113876 337316 241262
rect 337372 214564 337428 214574
rect 337372 165732 337428 214508
rect 337372 165666 337428 165676
rect 337260 113810 337316 113820
rect 338044 50372 338100 249902
rect 338380 249892 338436 249902
rect 338492 249508 338548 285902
rect 339276 269220 339332 269230
rect 339276 259498 339332 269164
rect 339276 259442 339444 259498
rect 339276 259364 339332 259374
rect 339276 258598 339332 259308
rect 338716 258542 339332 258598
rect 338268 249452 338548 249508
rect 338604 258418 338660 258428
rect 338268 245458 338324 249452
rect 338492 247078 338548 247088
rect 338268 245392 338324 245402
rect 338380 247022 338492 247078
rect 338380 220948 338436 247022
rect 338492 247012 338548 247022
rect 338380 220882 338436 220892
rect 338492 245098 338548 245108
rect 338380 197578 338436 197588
rect 338380 141092 338436 197522
rect 338380 141026 338436 141036
rect 338044 50306 338100 50316
rect 337148 46386 337204 46396
rect 336924 46162 336980 46172
rect 336812 41794 336868 41804
rect 338492 38052 338548 245042
rect 338604 42980 338660 258362
rect 338716 256798 338772 258542
rect 339276 258468 339332 258478
rect 339276 258352 339332 258362
rect 339276 257572 339332 257582
rect 338716 256742 338996 256798
rect 338716 256618 338772 256628
rect 338716 44578 338772 256562
rect 338940 254818 338996 256742
rect 339276 256078 339332 257516
rect 339388 256900 339444 259442
rect 339388 256834 339444 256844
rect 339388 256676 339444 256686
rect 339388 256618 339444 256620
rect 339388 256552 339444 256562
rect 339276 256022 339444 256078
rect 338716 44512 338772 44522
rect 338828 254762 338996 254818
rect 338828 43092 338884 254762
rect 339388 254098 339444 256022
rect 338828 43026 338884 43036
rect 338940 254042 339444 254098
rect 338604 42914 338660 42924
rect 338940 41524 338996 254042
rect 338940 41458 338996 41468
rect 339052 253862 339444 253918
rect 338492 37986 338548 37996
rect 339052 37940 339108 253862
rect 339388 253764 339444 253862
rect 339276 253738 339332 253748
rect 339388 253698 339444 253708
rect 339276 247978 339332 253682
rect 339276 247940 339444 247978
rect 339276 247922 339388 247940
rect 339388 247874 339444 247884
rect 339276 247716 339332 247726
rect 339276 247078 339332 247660
rect 339276 247012 339332 247022
rect 339276 246820 339332 246830
rect 339276 232708 339332 246764
rect 339388 245458 339444 245468
rect 339388 245364 339444 245402
rect 339388 245298 339444 245308
rect 339388 245140 339444 245150
rect 339388 245032 339444 245042
rect 339388 244918 339444 244954
rect 339388 244850 339444 244860
rect 339388 242004 339444 242014
rect 339388 236852 339444 241948
rect 339388 236786 339444 236796
rect 339276 232642 339332 232652
rect 339164 201236 339220 201246
rect 339164 139438 339220 201180
rect 339500 157798 339556 363244
rect 339612 291620 339668 407762
rect 339612 291554 339668 291564
rect 339724 407638 339780 407648
rect 339724 288932 339780 407582
rect 343338 400350 343958 408466
rect 343338 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 343958 400350
rect 343338 400226 343958 400294
rect 343338 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 343958 400226
rect 343338 400102 343958 400170
rect 343338 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 343958 400102
rect 343338 399978 343958 400046
rect 343338 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 343958 399978
rect 339948 397378 340004 397388
rect 339724 288866 339780 288876
rect 339836 296996 339892 297006
rect 339724 281764 339780 281774
rect 339612 261156 339668 261166
rect 339612 240238 339668 261100
rect 339724 241678 339780 281708
rect 339724 241612 339780 241622
rect 339612 240172 339668 240182
rect 339724 240660 339780 240670
rect 339724 240212 339780 240604
rect 339724 240146 339780 240156
rect 339724 210898 339780 210908
rect 339724 165060 339780 210842
rect 339724 164994 339780 165004
rect 339500 157732 339556 157742
rect 339164 139372 339220 139382
rect 339836 118916 339892 296940
rect 339948 295652 340004 397322
rect 343196 395218 343252 395228
rect 342860 392532 342916 392542
rect 342748 390718 342804 390728
rect 341852 380818 341908 380828
rect 340620 369572 340676 369582
rect 339948 295586 340004 295596
rect 340060 329364 340116 329374
rect 339948 277508 340004 277518
rect 339948 242004 340004 277452
rect 340060 262108 340116 329308
rect 340396 311332 340452 311342
rect 340060 262052 340340 262108
rect 340060 256900 340116 256910
rect 340060 253764 340116 256844
rect 340060 253698 340116 253708
rect 340172 252084 340228 252094
rect 340060 250068 340116 250078
rect 340060 249958 340116 250012
rect 340060 249892 340116 249902
rect 339948 241938 340004 241948
rect 339948 240212 340004 240222
rect 339948 238798 340004 240156
rect 339948 238732 340004 238742
rect 340060 238532 340116 238542
rect 339948 236852 340004 236862
rect 339948 194628 340004 236796
rect 340060 234478 340116 238476
rect 340060 234412 340116 234422
rect 339948 193284 340004 194572
rect 339948 193218 340004 193228
rect 339836 118850 339892 118860
rect 340172 41158 340228 252028
rect 340284 246596 340340 262052
rect 340396 247044 340452 311276
rect 340396 246978 340452 246988
rect 340284 246530 340340 246540
rect 340284 193978 340340 193988
rect 340284 160498 340340 193922
rect 340396 193284 340452 193294
rect 340396 183204 340452 193228
rect 340396 183138 340452 183148
rect 340620 161218 340676 369516
rect 341852 349468 341908 380762
rect 341852 349412 342468 349468
rect 342076 326564 342132 326574
rect 341964 325668 342020 325678
rect 341068 321188 341124 321198
rect 340620 161152 340676 161162
rect 340732 296100 340788 296110
rect 340284 160432 340340 160442
rect 340732 115892 340788 296044
rect 341068 256228 341124 321132
rect 341180 319396 341236 319406
rect 341180 277284 341236 319340
rect 341292 314020 341348 314030
rect 341292 280532 341348 313964
rect 341404 310436 341460 310446
rect 341404 299012 341460 310380
rect 341404 298946 341460 298956
rect 341292 280466 341348 280476
rect 341852 298788 341908 298798
rect 341180 277218 341236 277228
rect 341404 279972 341460 279982
rect 341068 256162 341124 256172
rect 341292 246932 341348 246942
rect 340956 242004 341012 242014
rect 340844 240212 340900 240222
rect 340844 238618 340900 240156
rect 340844 238552 340900 238562
rect 340732 115826 340788 115836
rect 340956 48580 341012 241948
rect 341292 241498 341348 246876
rect 341292 241432 341348 241442
rect 341404 243684 341460 279916
rect 341404 239988 341460 243628
rect 341404 239922 341460 239932
rect 341068 192358 341124 192368
rect 341068 157892 341124 192302
rect 341068 157826 341124 157836
rect 341852 124740 341908 298732
rect 341964 156178 342020 325612
rect 342076 160678 342132 326508
rect 342412 320964 342468 349412
rect 342300 305060 342356 305070
rect 342076 160612 342132 160622
rect 342188 302372 342244 302382
rect 341964 156112 342020 156122
rect 342076 151172 342132 151182
rect 342076 149698 342132 151116
rect 342076 149632 342132 149642
rect 342188 136388 342244 302316
rect 342300 145124 342356 305004
rect 342412 241318 342468 320908
rect 342748 289828 342804 390662
rect 342860 344484 342916 392476
rect 343196 374052 343252 395162
rect 343196 373986 343252 373996
rect 343338 382350 343958 399922
rect 347058 406350 347678 408466
rect 352492 408100 352548 408110
rect 347058 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 347678 406350
rect 347058 406226 347678 406294
rect 347058 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 347678 406226
rect 347058 406102 347678 406170
rect 347058 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 347678 406102
rect 347058 405978 347678 406046
rect 347058 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 347678 405978
rect 343338 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 343958 382350
rect 343338 382226 343958 382294
rect 343338 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 343958 382226
rect 343338 382102 343958 382170
rect 343338 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 343958 382102
rect 343338 381978 343958 382046
rect 343338 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 343958 381978
rect 342860 344418 342916 344428
rect 343338 364350 343958 381922
rect 344092 398638 344148 398648
rect 344092 373156 344148 398582
rect 344092 373090 344148 373100
rect 344204 395398 344260 395408
rect 344204 371364 344260 395342
rect 344204 371298 344260 371308
rect 347058 388350 347678 405922
rect 347058 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 347678 388350
rect 347058 388226 347678 388294
rect 347058 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 347678 388226
rect 347058 388102 347678 388170
rect 347058 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 347678 388102
rect 347058 387978 347678 388046
rect 347058 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 347678 387978
rect 347058 370350 347678 387922
rect 348572 407278 348628 407288
rect 348572 384244 348628 407222
rect 352492 406644 352548 408044
rect 348572 384178 348628 384188
rect 352044 385028 352100 385038
rect 347058 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 347678 370350
rect 347058 370226 347678 370294
rect 347058 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 347678 370226
rect 347058 370102 347678 370170
rect 347058 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 347678 370102
rect 347058 369978 347678 370046
rect 347058 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 347678 369978
rect 343338 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 343958 364350
rect 343338 364226 343958 364294
rect 343338 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 343958 364226
rect 343338 364102 343958 364170
rect 343338 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 343958 364102
rect 343338 363978 343958 364046
rect 343338 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 343958 363978
rect 343338 346350 343958 363922
rect 343338 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 343958 346350
rect 343338 346226 343958 346294
rect 343338 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 343958 346226
rect 343338 346102 343958 346170
rect 343338 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 343958 346102
rect 343338 345978 343958 346046
rect 343338 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 343958 345978
rect 342748 289762 342804 289772
rect 343338 328350 343958 345922
rect 346892 368676 346948 368686
rect 346780 335524 346836 335534
rect 346556 334628 346612 334638
rect 346108 332836 346164 332846
rect 345548 331044 345604 331054
rect 343338 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 343958 328350
rect 343338 328226 343958 328294
rect 343338 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 343958 328226
rect 343338 328102 343958 328170
rect 343338 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 343958 328102
rect 343338 327978 343958 328046
rect 343338 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 343958 327978
rect 343338 310350 343958 327922
rect 344988 328356 345044 328366
rect 343338 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 343958 310350
rect 343338 310226 343958 310294
rect 343338 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 343958 310226
rect 343338 310102 343958 310170
rect 343338 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 343958 310102
rect 343338 309978 343958 310046
rect 343338 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 343958 309978
rect 343338 292350 343958 309922
rect 343338 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 343958 292350
rect 343338 292226 343958 292294
rect 343338 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 343958 292226
rect 343338 292102 343958 292170
rect 343338 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 343958 292102
rect 343338 291978 343958 292046
rect 343338 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 343958 291978
rect 343338 274350 343958 291922
rect 343338 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 343958 274350
rect 343338 274226 343958 274294
rect 343338 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 343958 274226
rect 343338 274102 343958 274170
rect 343338 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 343958 274102
rect 343338 273978 343958 274046
rect 343338 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 343958 273978
rect 343084 266532 343140 266542
rect 342860 265636 342916 265646
rect 342636 257012 342692 257022
rect 342524 247044 342580 247054
rect 342524 242004 342580 246988
rect 342636 243628 342692 256956
rect 342636 243572 342804 243628
rect 342524 241938 342580 241948
rect 342412 241252 342468 241262
rect 342748 240418 342804 243572
rect 342860 241138 342916 265580
rect 342860 241072 342916 241082
rect 342972 262052 343028 262062
rect 342524 240362 342804 240418
rect 342524 147812 342580 240362
rect 342636 239540 342692 239550
rect 342636 238978 342692 239484
rect 342972 239092 343028 261996
rect 343084 239652 343140 266476
rect 343338 256350 343958 273922
rect 344092 320292 344148 320302
rect 344092 262164 344148 320236
rect 344876 317604 344932 317614
rect 344652 316708 344708 316718
rect 344540 315812 344596 315822
rect 344428 307748 344484 307758
rect 344428 299124 344484 307692
rect 344428 299058 344484 299068
rect 344316 287140 344372 287150
rect 344092 262098 344148 262108
rect 344204 280868 344260 280878
rect 343338 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 343958 256350
rect 343338 256226 343958 256294
rect 343338 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 343958 256226
rect 343338 256102 343958 256170
rect 343338 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 343958 256102
rect 343338 255978 343958 256046
rect 343338 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 343958 255978
rect 343084 239586 343140 239596
rect 343196 248612 343252 248622
rect 342972 239026 343028 239036
rect 342636 238912 342692 238922
rect 343196 236180 343252 248556
rect 343196 236114 343252 236124
rect 343338 238350 343958 255922
rect 344204 255388 344260 280812
rect 344316 262918 344372 287084
rect 344316 262852 344372 262862
rect 344540 258692 344596 315756
rect 344652 262388 344708 316652
rect 344764 312228 344820 312238
rect 344764 283892 344820 312172
rect 344764 283826 344820 283836
rect 344652 262322 344708 262332
rect 344764 282660 344820 282670
rect 344540 258626 344596 258636
rect 344204 255332 344596 255388
rect 344428 253092 344484 253102
rect 344428 238756 344484 253036
rect 344540 246708 344596 255332
rect 344540 239204 344596 246652
rect 344652 251300 344708 251310
rect 344652 245252 344708 251244
rect 344652 245186 344708 245196
rect 344764 241858 344820 282604
rect 344876 282212 344932 317548
rect 344876 282146 344932 282156
rect 344988 257012 345044 328300
rect 345324 324772 345380 324782
rect 345212 299684 345268 299694
rect 344988 256946 345044 256956
rect 345100 262164 345156 262174
rect 345100 252980 345156 262108
rect 345100 252914 345156 252924
rect 344764 240418 344820 241802
rect 344764 240352 344820 240362
rect 344540 239138 344596 239148
rect 344428 238690 344484 238700
rect 343338 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 343958 238350
rect 343338 238226 343958 238294
rect 343338 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 343958 238226
rect 343338 238102 343958 238170
rect 343338 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 343958 238102
rect 343338 237978 343958 238046
rect 343338 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 343958 237978
rect 342524 147746 342580 147756
rect 343338 220350 343958 237922
rect 343338 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 343958 220350
rect 343338 220226 343958 220294
rect 343338 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 343958 220226
rect 343338 220102 343958 220170
rect 343338 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 343958 220102
rect 343338 219978 343958 220046
rect 343338 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 343958 219978
rect 343338 202350 343958 219922
rect 343338 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 343958 202350
rect 343338 202226 343958 202294
rect 343338 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 343958 202226
rect 343338 202102 343958 202170
rect 343338 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 343958 202102
rect 343338 201978 343958 202046
rect 343338 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 343958 201978
rect 343338 184350 343958 201922
rect 344316 234388 344372 234398
rect 344204 201012 344260 201022
rect 343338 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 343958 184350
rect 343338 184226 343958 184294
rect 343338 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 343958 184226
rect 343338 184102 343958 184170
rect 343338 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 343958 184102
rect 343338 183978 343958 184046
rect 343338 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 343958 183978
rect 343338 166350 343958 183922
rect 343338 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 343958 166350
rect 343338 166226 343958 166294
rect 343338 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 343958 166226
rect 343338 166102 343958 166170
rect 343338 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 343958 166102
rect 343338 165978 343958 166046
rect 343338 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 343958 165978
rect 343338 148350 343958 165922
rect 343338 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 343958 148350
rect 343338 148226 343958 148294
rect 343338 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 343958 148226
rect 343338 148102 343958 148170
rect 343338 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 343958 148102
rect 343338 147978 343958 148046
rect 343338 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 343958 147978
rect 342300 145058 342356 145068
rect 342188 136322 342244 136332
rect 341852 124674 341908 124684
rect 343338 130350 343958 147922
rect 344092 197398 344148 197408
rect 344092 139188 344148 197342
rect 344204 158698 344260 200956
rect 344204 158632 344260 158642
rect 344092 139122 344148 139132
rect 343338 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 343958 130350
rect 343338 130226 343958 130294
rect 343338 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 343958 130226
rect 343338 130102 343958 130170
rect 343338 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 343958 130102
rect 343338 129978 343958 130046
rect 343338 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 343958 129978
rect 343338 112350 343958 129922
rect 343338 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 343958 112350
rect 343338 112226 343958 112294
rect 343338 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 343958 112226
rect 343338 112102 343958 112170
rect 343338 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 343958 112102
rect 343338 111978 343958 112046
rect 343338 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 343958 111978
rect 342524 95732 342580 95742
rect 342524 94978 342580 95676
rect 342524 94912 342580 94922
rect 340956 48514 341012 48524
rect 343338 94350 343958 111922
rect 344316 98308 344372 234332
rect 345212 127652 345268 299628
rect 345324 155458 345380 324716
rect 345324 155392 345380 155402
rect 345436 301476 345492 301486
rect 345436 133476 345492 301420
rect 345548 252756 345604 330988
rect 346108 280532 346164 332780
rect 346108 280466 346164 280476
rect 346220 279076 346276 279086
rect 346220 267148 346276 279020
rect 346108 267092 346276 267148
rect 346108 258598 346164 267092
rect 345548 252690 345604 252700
rect 345660 258542 346164 258598
rect 345436 133410 345492 133420
rect 345548 240418 345604 240428
rect 345212 127586 345268 127596
rect 345548 98420 345604 240362
rect 345660 236628 345716 258542
rect 345996 257012 346052 257022
rect 345660 189252 345716 236572
rect 345884 245252 345940 245262
rect 345660 189186 345716 189196
rect 345772 211078 345828 211088
rect 345772 166180 345828 211022
rect 345772 166114 345828 166124
rect 345884 113092 345940 245196
rect 345884 113026 345940 113036
rect 345548 98354 345604 98364
rect 344316 98242 344372 98252
rect 343338 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 343958 94350
rect 343338 94226 343958 94294
rect 343338 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 343958 94226
rect 343338 94102 343958 94170
rect 343338 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 343958 94102
rect 343338 93978 343958 94046
rect 343338 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 343958 93978
rect 343338 76350 343958 93922
rect 343338 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 343958 76350
rect 343338 76226 343958 76294
rect 343338 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 343958 76226
rect 343338 76102 343958 76170
rect 343338 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 343958 76102
rect 343338 75978 343958 76046
rect 343338 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 343958 75978
rect 343338 58350 343958 75922
rect 343338 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 343958 58350
rect 343338 58226 343958 58294
rect 343338 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 343958 58226
rect 343338 58102 343958 58170
rect 343338 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 343958 58102
rect 343338 57978 343958 58046
rect 343338 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 343958 57978
rect 340172 41092 340228 41102
rect 339052 37874 339108 37884
rect 343338 40350 343958 57922
rect 345996 48356 346052 256956
rect 346108 245924 346164 245934
rect 346108 234298 346164 245868
rect 346108 234232 346164 234242
rect 346332 161028 346388 161038
rect 346332 160858 346388 160972
rect 346332 160792 346388 160802
rect 346108 157892 346164 157902
rect 346108 157438 346164 157836
rect 346108 157372 346164 157382
rect 346556 150418 346612 334572
rect 346668 331940 346724 331950
rect 346668 156100 346724 331884
rect 346668 156034 346724 156044
rect 346556 150352 346612 150362
rect 346780 148618 346836 335468
rect 346892 162838 346948 368620
rect 346892 162772 346948 162782
rect 347058 352350 347678 369922
rect 347058 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 347678 352350
rect 347058 352226 347678 352294
rect 347058 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 347678 352226
rect 347058 352102 347678 352170
rect 347058 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 347678 352102
rect 347058 351978 347678 352046
rect 347058 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 347678 351978
rect 347058 334350 347678 351922
rect 351932 340452 351988 340462
rect 347058 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 347678 334350
rect 347058 334226 347678 334294
rect 347058 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 347678 334226
rect 347058 334102 347678 334170
rect 347058 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 347678 334102
rect 347058 333978 347678 334046
rect 347058 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 347678 333978
rect 347058 316350 347678 333922
rect 350028 334404 350084 334414
rect 347058 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 347678 316350
rect 347058 316226 347678 316294
rect 347058 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 347678 316226
rect 347058 316102 347678 316170
rect 347058 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 347678 316102
rect 347058 315978 347678 316046
rect 347058 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 347678 315978
rect 347058 298350 347678 315922
rect 347058 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 347678 298350
rect 347058 298226 347678 298294
rect 347058 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 347678 298226
rect 347058 298102 347678 298170
rect 347058 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 347678 298102
rect 347058 297978 347678 298046
rect 347058 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 347678 297978
rect 347058 280350 347678 297922
rect 348684 333732 348740 333742
rect 348012 295204 348068 295214
rect 347058 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 347678 280350
rect 347058 280226 347678 280294
rect 347058 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 347678 280226
rect 347058 280102 347678 280170
rect 347058 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 347678 280102
rect 347058 279978 347678 280046
rect 347058 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 347678 279978
rect 347058 262350 347678 279922
rect 347058 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 347678 262350
rect 347058 262226 347678 262294
rect 347058 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 347678 262226
rect 347058 262102 347678 262170
rect 347058 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 347678 262102
rect 347058 261978 347678 262046
rect 347058 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 347678 261978
rect 347058 244350 347678 261922
rect 347788 291620 347844 291630
rect 347788 246932 347844 291564
rect 347788 246866 347844 246876
rect 347900 283556 347956 283566
rect 347058 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 347678 244350
rect 347058 244226 347678 244294
rect 347058 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 347678 244226
rect 347058 244102 347678 244170
rect 347058 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 347678 244102
rect 347058 243978 347678 244046
rect 347058 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 347678 243978
rect 347058 226350 347678 243922
rect 347900 240660 347956 283500
rect 348012 273028 348068 295148
rect 348012 272962 348068 272972
rect 348572 288932 348628 288942
rect 347900 240324 347956 240604
rect 347900 240258 347956 240268
rect 348460 246596 348516 246606
rect 347058 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 347678 226350
rect 347058 226226 347678 226294
rect 347058 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 347678 226226
rect 347058 226102 347678 226170
rect 347058 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 347678 226102
rect 347058 225978 347678 226046
rect 347058 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 347678 225978
rect 347058 208350 347678 225922
rect 347058 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 347678 208350
rect 347058 208226 347678 208294
rect 347058 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 347678 208226
rect 347058 208102 347678 208170
rect 347058 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 347678 208102
rect 347058 207978 347678 208046
rect 347058 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 347678 207978
rect 347058 190350 347678 207922
rect 347058 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 347678 190350
rect 347058 190226 347678 190294
rect 347058 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 347678 190226
rect 347058 190102 347678 190170
rect 347058 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 347678 190102
rect 347058 189978 347678 190046
rect 347058 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 347678 189978
rect 347058 172350 347678 189922
rect 347058 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 347678 172350
rect 347058 172226 347678 172294
rect 347058 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 347678 172226
rect 347058 172102 347678 172170
rect 347058 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 347678 172102
rect 347058 171978 347678 172046
rect 347058 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 347678 171978
rect 346892 159572 346948 159582
rect 346892 157978 346948 159516
rect 346892 157912 346948 157922
rect 346780 148552 346836 148562
rect 347058 154350 347678 171922
rect 348460 162118 348516 246540
rect 348460 162052 348516 162062
rect 347058 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 347678 154350
rect 347058 154226 347678 154294
rect 347058 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 347678 154226
rect 347058 154102 347678 154170
rect 347058 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 347678 154102
rect 347058 153978 347678 154046
rect 347058 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 347678 153978
rect 345996 48290 346052 48300
rect 347058 136350 347678 153922
rect 347058 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 347678 136350
rect 347058 136226 347678 136294
rect 347058 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 347678 136226
rect 347058 136102 347678 136170
rect 347058 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 347678 136102
rect 347058 135978 347678 136046
rect 347058 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 347678 135978
rect 347058 118350 347678 135922
rect 347058 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 347678 118350
rect 347058 118226 347678 118294
rect 347058 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 347678 118226
rect 347058 118102 347678 118170
rect 347058 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 347678 118102
rect 347058 117978 347678 118046
rect 347058 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 347678 117978
rect 347058 100350 347678 117922
rect 347058 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 347678 100350
rect 347058 100226 347678 100294
rect 347058 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 347678 100226
rect 347058 100102 347678 100170
rect 347058 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 347678 100102
rect 347058 99978 347678 100046
rect 347058 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 347678 99978
rect 347058 82350 347678 99922
rect 348572 98756 348628 288876
rect 348684 152578 348740 333676
rect 348908 327460 348964 327470
rect 348684 152512 348740 152522
rect 348796 243684 348852 243694
rect 348572 98690 348628 98700
rect 348796 98532 348852 243628
rect 348908 147476 348964 327404
rect 349020 322084 349076 322094
rect 349020 149380 349076 322028
rect 349132 318500 349188 318510
rect 349132 157892 349188 318444
rect 349580 294308 349636 294318
rect 349468 292404 349524 292414
rect 349468 249508 349524 292348
rect 349580 252084 349636 294252
rect 349580 252018 349636 252028
rect 349692 289828 349748 289838
rect 349468 249442 349524 249452
rect 349692 247828 349748 289772
rect 349692 247762 349748 247772
rect 349132 157826 349188 157836
rect 349244 240324 349300 240334
rect 349020 149314 349076 149324
rect 348908 147410 348964 147420
rect 349244 98644 349300 240268
rect 349356 181188 349412 181198
rect 349356 145738 349412 181132
rect 350028 147718 350084 334348
rect 350588 323876 350644 323886
rect 350364 322980 350420 322990
rect 350140 252756 350196 252766
rect 350140 152038 350196 252700
rect 350140 151972 350196 151982
rect 350252 246820 350308 246830
rect 350028 147652 350084 147662
rect 349356 145672 349412 145682
rect 350252 98868 350308 246764
rect 350364 150598 350420 322924
rect 350364 150532 350420 150542
rect 350476 303268 350532 303278
rect 350476 139300 350532 303212
rect 350588 152218 350644 323820
rect 350812 313124 350868 313134
rect 350588 152152 350644 152162
rect 350700 246708 350756 246718
rect 350476 139234 350532 139244
rect 350700 98980 350756 246652
rect 350812 163738 350868 313068
rect 351148 297892 351204 297902
rect 351148 196588 351204 297836
rect 351260 275492 351316 275502
rect 351260 261268 351316 275436
rect 351260 261202 351316 261212
rect 351820 257012 351876 257022
rect 351820 245252 351876 256956
rect 351820 245186 351876 245196
rect 350812 163672 350868 163682
rect 350924 196532 351204 196588
rect 351820 231588 351876 231598
rect 350812 152516 350868 152526
rect 350812 151284 350868 152460
rect 350812 146098 350868 151228
rect 350812 146032 350868 146042
rect 350924 121828 350980 196532
rect 351820 183876 351876 231532
rect 351820 183316 351876 183820
rect 351820 183250 351876 183260
rect 351820 167748 351876 167758
rect 351820 167338 351876 167692
rect 351820 167272 351876 167282
rect 351036 146244 351092 146254
rect 351036 141058 351092 146188
rect 351932 146244 351988 340396
rect 352044 292068 352100 384972
rect 352268 366212 352324 366222
rect 352268 364644 352324 366156
rect 352268 361228 352324 364588
rect 352044 292002 352100 292012
rect 352156 361172 352324 361228
rect 352044 268772 352100 268782
rect 352044 267876 352100 268716
rect 352044 151172 352100 267820
rect 352156 153860 352212 361172
rect 352156 153794 352212 153804
rect 352268 261828 352324 261838
rect 352268 152516 352324 261772
rect 352492 257012 352548 406588
rect 352492 256946 352548 256956
rect 352604 407540 352660 407550
rect 352604 249732 352660 407484
rect 353836 406918 353892 406928
rect 353612 406738 353668 406748
rect 353612 387716 353668 406682
rect 353612 387650 353668 387660
rect 353836 387604 353892 406862
rect 354396 406644 354452 409742
rect 354396 406578 354452 406588
rect 355292 407098 355348 407108
rect 355180 397378 355236 397388
rect 355068 397198 355124 397208
rect 353836 387538 353892 387548
rect 354956 395220 355012 395230
rect 354956 386036 355012 395164
rect 355068 390516 355124 397142
rect 355180 391412 355236 397322
rect 355292 395220 355348 407042
rect 355292 395154 355348 395164
rect 355180 391346 355236 391356
rect 355292 395038 355348 395048
rect 355292 391300 355348 394982
rect 355292 391234 355348 391244
rect 355404 390852 355460 410060
rect 357756 409618 357812 409628
rect 356076 409078 356132 409088
rect 356076 407428 356132 409022
rect 356748 408548 356804 408558
rect 356524 408212 356580 408222
rect 356076 407362 356132 407372
rect 356412 407428 356468 407438
rect 355404 390786 355460 390796
rect 355516 401604 355572 401614
rect 355068 390450 355124 390460
rect 354956 385970 355012 385980
rect 355516 383012 355572 401548
rect 355740 400618 355796 400628
rect 355740 396508 355796 400562
rect 355628 396452 355796 396508
rect 356076 397018 356132 397028
rect 355628 389508 355684 396452
rect 356076 391078 356132 396962
rect 356412 392518 356468 407372
rect 356412 392452 356468 392462
rect 356524 392338 356580 408156
rect 356524 392272 356580 392282
rect 356636 395108 356692 395118
rect 356076 391012 356132 391022
rect 356636 390898 356692 395052
rect 356636 390832 356692 390842
rect 355628 389442 355684 389452
rect 355516 382946 355572 382956
rect 355292 367780 355348 367790
rect 353612 360612 353668 360622
rect 352492 245252 352548 245262
rect 352492 243684 352548 245196
rect 352268 152450 352324 152460
rect 352380 198212 352436 198222
rect 352044 151106 352100 151116
rect 352380 149548 352436 198156
rect 351932 146178 351988 146188
rect 352044 149492 352436 149548
rect 351036 140992 351092 141002
rect 351932 143938 351988 143948
rect 350924 121762 350980 121772
rect 350700 98914 350756 98924
rect 350252 98802 350308 98812
rect 349244 98578 349300 98588
rect 348796 98466 348852 98476
rect 351932 91588 351988 143882
rect 352044 140878 352100 149492
rect 352044 128548 352100 140822
rect 352044 128482 352100 128492
rect 352492 144298 352548 243628
rect 352492 126028 352548 144242
rect 352604 144478 352660 249676
rect 352604 143938 352660 144422
rect 352604 143872 352660 143882
rect 352716 346500 352772 346510
rect 352716 142678 352772 346444
rect 353388 293188 353444 293198
rect 352828 291508 352884 291518
rect 352828 252084 352884 291452
rect 353388 284788 353444 293132
rect 353388 284722 353444 284732
rect 353500 286020 353556 286030
rect 352828 252018 352884 252028
rect 352940 262918 352996 262928
rect 352940 236628 352996 262862
rect 352940 236562 352996 236572
rect 353500 234658 353556 285964
rect 353500 162478 353556 234602
rect 353500 162412 353556 162422
rect 353612 157618 353668 360556
rect 353612 157552 353668 157562
rect 353724 329252 353780 329262
rect 352716 142612 352772 142622
rect 353724 140980 353780 329196
rect 355068 328356 355124 328366
rect 354396 322308 354452 322318
rect 354396 320964 354452 322252
rect 354060 305956 354116 305966
rect 353948 300580 354004 300590
rect 353724 140914 353780 140924
rect 353836 278964 353892 278974
rect 352156 125972 352548 126028
rect 352156 107156 352212 125972
rect 352156 107090 352212 107100
rect 353836 105140 353892 278908
rect 353948 130564 354004 300524
rect 354060 147364 354116 305900
rect 354172 252980 354228 252990
rect 354172 158878 354228 252924
rect 354284 236852 354340 236862
rect 354284 165538 354340 236796
rect 354284 165472 354340 165482
rect 354396 162298 354452 320908
rect 354508 306852 354564 306862
rect 354508 183428 354564 306796
rect 354508 183362 354564 183372
rect 354732 304276 354788 304286
rect 354396 162232 354452 162242
rect 354172 158812 354228 158822
rect 354060 147298 354116 147308
rect 354732 142212 354788 304220
rect 354844 304164 354900 304174
rect 354844 302428 354900 304108
rect 354844 302372 355012 302428
rect 354732 142146 354788 142156
rect 354844 189252 354900 189262
rect 353948 130498 354004 130508
rect 353836 105074 353892 105084
rect 353948 99092 354004 99102
rect 353948 98218 354004 99036
rect 354844 99092 354900 189196
rect 354956 164098 355012 302372
rect 354956 164032 355012 164042
rect 355068 163918 355124 328300
rect 355068 163852 355124 163862
rect 355180 292068 355236 292078
rect 355180 155638 355236 292012
rect 355292 159598 355348 367724
rect 355628 285684 355684 285694
rect 355516 281764 355572 281774
rect 355404 236638 355460 236648
rect 355404 236544 355460 236572
rect 355404 213598 355460 213608
rect 355404 213444 355460 213542
rect 355404 213378 355460 213388
rect 355292 159532 355348 159542
rect 355404 183204 355460 183214
rect 355180 155572 355236 155582
rect 354844 99026 354900 99036
rect 353948 98152 354004 98162
rect 355404 98196 355460 183148
rect 355516 101668 355572 281708
rect 355628 110068 355684 285628
rect 356636 236638 356692 236648
rect 356524 167338 356580 167348
rect 356076 166292 356132 166302
rect 356076 164818 356132 166236
rect 356076 164752 356132 164762
rect 356524 156996 356580 167282
rect 356524 156930 356580 156940
rect 355628 110002 355684 110012
rect 355516 101602 355572 101612
rect 355404 98130 355460 98140
rect 356636 97300 356692 236582
rect 356748 213598 356804 408492
rect 357756 407204 357812 409562
rect 444332 409444 444388 590156
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 466218 562350 466838 579922
rect 466218 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 466838 562350
rect 466218 562226 466838 562294
rect 466218 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 466838 562226
rect 466218 562102 466838 562170
rect 466218 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 466838 562102
rect 466218 561978 466838 562046
rect 466218 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 466838 561978
rect 455568 550350 455888 550384
rect 455568 550294 455638 550350
rect 455694 550294 455762 550350
rect 455818 550294 455888 550350
rect 455568 550226 455888 550294
rect 455568 550170 455638 550226
rect 455694 550170 455762 550226
rect 455818 550170 455888 550226
rect 455568 550102 455888 550170
rect 455568 550046 455638 550102
rect 455694 550046 455762 550102
rect 455818 550046 455888 550102
rect 455568 549978 455888 550046
rect 455568 549922 455638 549978
rect 455694 549922 455762 549978
rect 455818 549922 455888 549978
rect 455568 549888 455888 549922
rect 466218 544350 466838 561922
rect 466218 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 466838 544350
rect 466218 544226 466838 544294
rect 466218 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 466838 544226
rect 466218 544102 466838 544170
rect 466218 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 466838 544102
rect 466218 543978 466838 544046
rect 466218 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 466838 543978
rect 455568 532350 455888 532384
rect 455568 532294 455638 532350
rect 455694 532294 455762 532350
rect 455818 532294 455888 532350
rect 455568 532226 455888 532294
rect 455568 532170 455638 532226
rect 455694 532170 455762 532226
rect 455818 532170 455888 532226
rect 455568 532102 455888 532170
rect 455568 532046 455638 532102
rect 455694 532046 455762 532102
rect 455818 532046 455888 532102
rect 455568 531978 455888 532046
rect 455568 531922 455638 531978
rect 455694 531922 455762 531978
rect 455818 531922 455888 531978
rect 455568 531888 455888 531922
rect 466218 526350 466838 543922
rect 466218 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 466838 526350
rect 466218 526226 466838 526294
rect 466218 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 466838 526226
rect 466218 526102 466838 526170
rect 466218 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 466838 526102
rect 466218 525978 466838 526046
rect 466218 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 466838 525978
rect 455568 514350 455888 514384
rect 455568 514294 455638 514350
rect 455694 514294 455762 514350
rect 455818 514294 455888 514350
rect 455568 514226 455888 514294
rect 455568 514170 455638 514226
rect 455694 514170 455762 514226
rect 455818 514170 455888 514226
rect 455568 514102 455888 514170
rect 455568 514046 455638 514102
rect 455694 514046 455762 514102
rect 455818 514046 455888 514102
rect 455568 513978 455888 514046
rect 455568 513922 455638 513978
rect 455694 513922 455762 513978
rect 455818 513922 455888 513978
rect 455568 513888 455888 513922
rect 466218 508350 466838 525922
rect 466218 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 466838 508350
rect 466218 508226 466838 508294
rect 466218 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 466838 508226
rect 466218 508102 466838 508170
rect 466218 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 466838 508102
rect 466218 507978 466838 508046
rect 466218 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 466838 507978
rect 455568 496350 455888 496384
rect 455568 496294 455638 496350
rect 455694 496294 455762 496350
rect 455818 496294 455888 496350
rect 455568 496226 455888 496294
rect 455568 496170 455638 496226
rect 455694 496170 455762 496226
rect 455818 496170 455888 496226
rect 455568 496102 455888 496170
rect 455568 496046 455638 496102
rect 455694 496046 455762 496102
rect 455818 496046 455888 496102
rect 455568 495978 455888 496046
rect 455568 495922 455638 495978
rect 455694 495922 455762 495978
rect 455818 495922 455888 495978
rect 455568 495888 455888 495922
rect 466218 490350 466838 507922
rect 466218 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 466838 490350
rect 466218 490226 466838 490294
rect 466218 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 466838 490226
rect 466218 490102 466838 490170
rect 466218 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 466838 490102
rect 466218 489978 466838 490046
rect 466218 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 466838 489978
rect 455568 478350 455888 478384
rect 455568 478294 455638 478350
rect 455694 478294 455762 478350
rect 455818 478294 455888 478350
rect 455568 478226 455888 478294
rect 455568 478170 455638 478226
rect 455694 478170 455762 478226
rect 455818 478170 455888 478226
rect 455568 478102 455888 478170
rect 455568 478046 455638 478102
rect 455694 478046 455762 478102
rect 455818 478046 455888 478102
rect 455568 477978 455888 478046
rect 455568 477922 455638 477978
rect 455694 477922 455762 477978
rect 455818 477922 455888 477978
rect 455568 477888 455888 477922
rect 466218 472350 466838 489922
rect 466218 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 466838 472350
rect 466218 472226 466838 472294
rect 466218 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 466838 472226
rect 466218 472102 466838 472170
rect 466218 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 466838 472102
rect 466218 471978 466838 472046
rect 466218 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 466838 471978
rect 455568 460350 455888 460384
rect 455568 460294 455638 460350
rect 455694 460294 455762 460350
rect 455818 460294 455888 460350
rect 455568 460226 455888 460294
rect 455568 460170 455638 460226
rect 455694 460170 455762 460226
rect 455818 460170 455888 460226
rect 455568 460102 455888 460170
rect 455568 460046 455638 460102
rect 455694 460046 455762 460102
rect 455818 460046 455888 460102
rect 455568 459978 455888 460046
rect 455568 459922 455638 459978
rect 455694 459922 455762 459978
rect 455818 459922 455888 459978
rect 455568 459888 455888 459922
rect 466218 454350 466838 471922
rect 466218 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 466838 454350
rect 466218 454226 466838 454294
rect 466218 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 466838 454226
rect 466218 454102 466838 454170
rect 466218 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 466838 454102
rect 466218 453978 466838 454046
rect 466218 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 466838 453978
rect 455568 442350 455888 442384
rect 455568 442294 455638 442350
rect 455694 442294 455762 442350
rect 455818 442294 455888 442350
rect 455568 442226 455888 442294
rect 455568 442170 455638 442226
rect 455694 442170 455762 442226
rect 455818 442170 455888 442226
rect 455568 442102 455888 442170
rect 455568 442046 455638 442102
rect 455694 442046 455762 442102
rect 455818 442046 455888 442102
rect 455568 441978 455888 442046
rect 455568 441922 455638 441978
rect 455694 441922 455762 441978
rect 455818 441922 455888 441978
rect 455568 441888 455888 441922
rect 466218 436350 466838 453922
rect 466218 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 466838 436350
rect 466218 436226 466838 436294
rect 466218 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 466838 436226
rect 466218 436102 466838 436170
rect 466218 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 466838 436102
rect 466218 435978 466838 436046
rect 466218 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 466838 435978
rect 444332 409378 444388 409388
rect 446012 428518 446068 428528
rect 444892 407876 444948 407886
rect 444892 407278 444948 407820
rect 444892 407212 444948 407222
rect 357756 407138 357812 407148
rect 446012 406420 446068 428462
rect 455568 424350 455888 424384
rect 455568 424294 455638 424350
rect 455694 424294 455762 424350
rect 455818 424294 455888 424350
rect 455568 424226 455888 424294
rect 455568 424170 455638 424226
rect 455694 424170 455762 424226
rect 455818 424170 455888 424226
rect 455568 424102 455888 424170
rect 455568 424046 455638 424102
rect 455694 424046 455762 424102
rect 455818 424046 455888 424102
rect 455568 423978 455888 424046
rect 455568 423922 455638 423978
rect 455694 423922 455762 423978
rect 455818 423922 455888 423978
rect 455568 423888 455888 423922
rect 446012 406354 446068 406364
rect 466218 418350 466838 435922
rect 466218 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 466838 418350
rect 466218 418226 466838 418294
rect 466218 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 466838 418226
rect 466218 418102 466838 418170
rect 466218 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 466838 418102
rect 466218 417978 466838 418046
rect 466218 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 466838 417978
rect 466218 400350 466838 417922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 568350 470558 585922
rect 469938 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 470558 568350
rect 469938 568226 470558 568294
rect 469938 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 470558 568226
rect 469938 568102 470558 568170
rect 469938 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 470558 568102
rect 469938 567978 470558 568046
rect 469938 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 470558 567978
rect 469938 550350 470558 567922
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 470928 562350 471248 562384
rect 470928 562294 470998 562350
rect 471054 562294 471122 562350
rect 471178 562294 471248 562350
rect 470928 562226 471248 562294
rect 470928 562170 470998 562226
rect 471054 562170 471122 562226
rect 471178 562170 471248 562226
rect 470928 562102 471248 562170
rect 470928 562046 470998 562102
rect 471054 562046 471122 562102
rect 471178 562046 471248 562102
rect 470928 561978 471248 562046
rect 470928 561922 470998 561978
rect 471054 561922 471122 561978
rect 471178 561922 471248 561978
rect 470928 561888 471248 561922
rect 496938 562350 497558 579922
rect 496938 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 497558 562350
rect 496938 562226 497558 562294
rect 496938 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 497558 562226
rect 496938 562102 497558 562170
rect 496938 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 497558 562102
rect 496938 561978 497558 562046
rect 496938 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 497558 561978
rect 469938 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 470558 550350
rect 469938 550226 470558 550294
rect 469938 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 470558 550226
rect 469938 550102 470558 550170
rect 469938 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 470558 550102
rect 469938 549978 470558 550046
rect 469938 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 470558 549978
rect 469938 532350 470558 549922
rect 486288 550350 486608 550384
rect 486288 550294 486358 550350
rect 486414 550294 486482 550350
rect 486538 550294 486608 550350
rect 486288 550226 486608 550294
rect 486288 550170 486358 550226
rect 486414 550170 486482 550226
rect 486538 550170 486608 550226
rect 486288 550102 486608 550170
rect 486288 550046 486358 550102
rect 486414 550046 486482 550102
rect 486538 550046 486608 550102
rect 486288 549978 486608 550046
rect 486288 549922 486358 549978
rect 486414 549922 486482 549978
rect 486538 549922 486608 549978
rect 486288 549888 486608 549922
rect 470928 544350 471248 544384
rect 470928 544294 470998 544350
rect 471054 544294 471122 544350
rect 471178 544294 471248 544350
rect 470928 544226 471248 544294
rect 470928 544170 470998 544226
rect 471054 544170 471122 544226
rect 471178 544170 471248 544226
rect 470928 544102 471248 544170
rect 470928 544046 470998 544102
rect 471054 544046 471122 544102
rect 471178 544046 471248 544102
rect 470928 543978 471248 544046
rect 470928 543922 470998 543978
rect 471054 543922 471122 543978
rect 471178 543922 471248 543978
rect 470928 543888 471248 543922
rect 496938 544350 497558 561922
rect 496938 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 497558 544350
rect 496938 544226 497558 544294
rect 496938 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 497558 544226
rect 496938 544102 497558 544170
rect 496938 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 497558 544102
rect 496938 543978 497558 544046
rect 496938 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 497558 543978
rect 469938 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 470558 532350
rect 469938 532226 470558 532294
rect 469938 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 470558 532226
rect 469938 532102 470558 532170
rect 469938 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 470558 532102
rect 469938 531978 470558 532046
rect 469938 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 470558 531978
rect 469938 514350 470558 531922
rect 486288 532350 486608 532384
rect 486288 532294 486358 532350
rect 486414 532294 486482 532350
rect 486538 532294 486608 532350
rect 486288 532226 486608 532294
rect 486288 532170 486358 532226
rect 486414 532170 486482 532226
rect 486538 532170 486608 532226
rect 486288 532102 486608 532170
rect 486288 532046 486358 532102
rect 486414 532046 486482 532102
rect 486538 532046 486608 532102
rect 486288 531978 486608 532046
rect 486288 531922 486358 531978
rect 486414 531922 486482 531978
rect 486538 531922 486608 531978
rect 486288 531888 486608 531922
rect 470928 526350 471248 526384
rect 470928 526294 470998 526350
rect 471054 526294 471122 526350
rect 471178 526294 471248 526350
rect 470928 526226 471248 526294
rect 470928 526170 470998 526226
rect 471054 526170 471122 526226
rect 471178 526170 471248 526226
rect 470928 526102 471248 526170
rect 470928 526046 470998 526102
rect 471054 526046 471122 526102
rect 471178 526046 471248 526102
rect 470928 525978 471248 526046
rect 470928 525922 470998 525978
rect 471054 525922 471122 525978
rect 471178 525922 471248 525978
rect 470928 525888 471248 525922
rect 496938 526350 497558 543922
rect 496938 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 497558 526350
rect 496938 526226 497558 526294
rect 496938 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 497558 526226
rect 496938 526102 497558 526170
rect 496938 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 497558 526102
rect 496938 525978 497558 526046
rect 496938 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 497558 525978
rect 469938 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 470558 514350
rect 469938 514226 470558 514294
rect 469938 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 470558 514226
rect 469938 514102 470558 514170
rect 469938 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 470558 514102
rect 469938 513978 470558 514046
rect 469938 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 470558 513978
rect 469938 496350 470558 513922
rect 486288 514350 486608 514384
rect 486288 514294 486358 514350
rect 486414 514294 486482 514350
rect 486538 514294 486608 514350
rect 486288 514226 486608 514294
rect 486288 514170 486358 514226
rect 486414 514170 486482 514226
rect 486538 514170 486608 514226
rect 486288 514102 486608 514170
rect 486288 514046 486358 514102
rect 486414 514046 486482 514102
rect 486538 514046 486608 514102
rect 486288 513978 486608 514046
rect 486288 513922 486358 513978
rect 486414 513922 486482 513978
rect 486538 513922 486608 513978
rect 486288 513888 486608 513922
rect 470928 508350 471248 508384
rect 470928 508294 470998 508350
rect 471054 508294 471122 508350
rect 471178 508294 471248 508350
rect 470928 508226 471248 508294
rect 470928 508170 470998 508226
rect 471054 508170 471122 508226
rect 471178 508170 471248 508226
rect 470928 508102 471248 508170
rect 470928 508046 470998 508102
rect 471054 508046 471122 508102
rect 471178 508046 471248 508102
rect 470928 507978 471248 508046
rect 470928 507922 470998 507978
rect 471054 507922 471122 507978
rect 471178 507922 471248 507978
rect 470928 507888 471248 507922
rect 496938 508350 497558 525922
rect 496938 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 497558 508350
rect 496938 508226 497558 508294
rect 496938 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 497558 508226
rect 496938 508102 497558 508170
rect 496938 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 497558 508102
rect 496938 507978 497558 508046
rect 496938 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 497558 507978
rect 469938 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 470558 496350
rect 469938 496226 470558 496294
rect 469938 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 470558 496226
rect 469938 496102 470558 496170
rect 469938 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 470558 496102
rect 469938 495978 470558 496046
rect 469938 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 470558 495978
rect 469938 478350 470558 495922
rect 486288 496350 486608 496384
rect 486288 496294 486358 496350
rect 486414 496294 486482 496350
rect 486538 496294 486608 496350
rect 486288 496226 486608 496294
rect 486288 496170 486358 496226
rect 486414 496170 486482 496226
rect 486538 496170 486608 496226
rect 486288 496102 486608 496170
rect 486288 496046 486358 496102
rect 486414 496046 486482 496102
rect 486538 496046 486608 496102
rect 486288 495978 486608 496046
rect 486288 495922 486358 495978
rect 486414 495922 486482 495978
rect 486538 495922 486608 495978
rect 486288 495888 486608 495922
rect 470928 490350 471248 490384
rect 470928 490294 470998 490350
rect 471054 490294 471122 490350
rect 471178 490294 471248 490350
rect 470928 490226 471248 490294
rect 470928 490170 470998 490226
rect 471054 490170 471122 490226
rect 471178 490170 471248 490226
rect 470928 490102 471248 490170
rect 470928 490046 470998 490102
rect 471054 490046 471122 490102
rect 471178 490046 471248 490102
rect 470928 489978 471248 490046
rect 470928 489922 470998 489978
rect 471054 489922 471122 489978
rect 471178 489922 471248 489978
rect 470928 489888 471248 489922
rect 496938 490350 497558 507922
rect 496938 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 497558 490350
rect 496938 490226 497558 490294
rect 496938 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 497558 490226
rect 496938 490102 497558 490170
rect 496938 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 497558 490102
rect 496938 489978 497558 490046
rect 496938 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 497558 489978
rect 469938 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 470558 478350
rect 469938 478226 470558 478294
rect 469938 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 470558 478226
rect 469938 478102 470558 478170
rect 469938 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 470558 478102
rect 469938 477978 470558 478046
rect 469938 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 470558 477978
rect 469938 460350 470558 477922
rect 486288 478350 486608 478384
rect 486288 478294 486358 478350
rect 486414 478294 486482 478350
rect 486538 478294 486608 478350
rect 486288 478226 486608 478294
rect 486288 478170 486358 478226
rect 486414 478170 486482 478226
rect 486538 478170 486608 478226
rect 486288 478102 486608 478170
rect 486288 478046 486358 478102
rect 486414 478046 486482 478102
rect 486538 478046 486608 478102
rect 486288 477978 486608 478046
rect 486288 477922 486358 477978
rect 486414 477922 486482 477978
rect 486538 477922 486608 477978
rect 486288 477888 486608 477922
rect 470928 472350 471248 472384
rect 470928 472294 470998 472350
rect 471054 472294 471122 472350
rect 471178 472294 471248 472350
rect 470928 472226 471248 472294
rect 470928 472170 470998 472226
rect 471054 472170 471122 472226
rect 471178 472170 471248 472226
rect 470928 472102 471248 472170
rect 470928 472046 470998 472102
rect 471054 472046 471122 472102
rect 471178 472046 471248 472102
rect 470928 471978 471248 472046
rect 470928 471922 470998 471978
rect 471054 471922 471122 471978
rect 471178 471922 471248 471978
rect 470928 471888 471248 471922
rect 496938 472350 497558 489922
rect 496938 472294 497034 472350
rect 497090 472294 497158 472350
rect 497214 472294 497282 472350
rect 497338 472294 497406 472350
rect 497462 472294 497558 472350
rect 496938 472226 497558 472294
rect 496938 472170 497034 472226
rect 497090 472170 497158 472226
rect 497214 472170 497282 472226
rect 497338 472170 497406 472226
rect 497462 472170 497558 472226
rect 496938 472102 497558 472170
rect 496938 472046 497034 472102
rect 497090 472046 497158 472102
rect 497214 472046 497282 472102
rect 497338 472046 497406 472102
rect 497462 472046 497558 472102
rect 496938 471978 497558 472046
rect 496938 471922 497034 471978
rect 497090 471922 497158 471978
rect 497214 471922 497282 471978
rect 497338 471922 497406 471978
rect 497462 471922 497558 471978
rect 469938 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 470558 460350
rect 469938 460226 470558 460294
rect 469938 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 470558 460226
rect 469938 460102 470558 460170
rect 469938 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 470558 460102
rect 469938 459978 470558 460046
rect 469938 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 470558 459978
rect 469938 442350 470558 459922
rect 486288 460350 486608 460384
rect 486288 460294 486358 460350
rect 486414 460294 486482 460350
rect 486538 460294 486608 460350
rect 486288 460226 486608 460294
rect 486288 460170 486358 460226
rect 486414 460170 486482 460226
rect 486538 460170 486608 460226
rect 486288 460102 486608 460170
rect 486288 460046 486358 460102
rect 486414 460046 486482 460102
rect 486538 460046 486608 460102
rect 486288 459978 486608 460046
rect 486288 459922 486358 459978
rect 486414 459922 486482 459978
rect 486538 459922 486608 459978
rect 486288 459888 486608 459922
rect 470928 454350 471248 454384
rect 470928 454294 470998 454350
rect 471054 454294 471122 454350
rect 471178 454294 471248 454350
rect 470928 454226 471248 454294
rect 470928 454170 470998 454226
rect 471054 454170 471122 454226
rect 471178 454170 471248 454226
rect 470928 454102 471248 454170
rect 470928 454046 470998 454102
rect 471054 454046 471122 454102
rect 471178 454046 471248 454102
rect 470928 453978 471248 454046
rect 470928 453922 470998 453978
rect 471054 453922 471122 453978
rect 471178 453922 471248 453978
rect 470928 453888 471248 453922
rect 496938 454350 497558 471922
rect 496938 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 497558 454350
rect 496938 454226 497558 454294
rect 496938 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 497558 454226
rect 496938 454102 497558 454170
rect 496938 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 497558 454102
rect 496938 453978 497558 454046
rect 496938 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 497558 453978
rect 469938 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 470558 442350
rect 469938 442226 470558 442294
rect 469938 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 470558 442226
rect 469938 442102 470558 442170
rect 469938 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 470558 442102
rect 469938 441978 470558 442046
rect 469938 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 470558 441978
rect 469938 424350 470558 441922
rect 486288 442350 486608 442384
rect 486288 442294 486358 442350
rect 486414 442294 486482 442350
rect 486538 442294 486608 442350
rect 486288 442226 486608 442294
rect 486288 442170 486358 442226
rect 486414 442170 486482 442226
rect 486538 442170 486608 442226
rect 486288 442102 486608 442170
rect 486288 442046 486358 442102
rect 486414 442046 486482 442102
rect 486538 442046 486608 442102
rect 486288 441978 486608 442046
rect 486288 441922 486358 441978
rect 486414 441922 486482 441978
rect 486538 441922 486608 441978
rect 486288 441888 486608 441922
rect 470928 436350 471248 436384
rect 470928 436294 470998 436350
rect 471054 436294 471122 436350
rect 471178 436294 471248 436350
rect 470928 436226 471248 436294
rect 470928 436170 470998 436226
rect 471054 436170 471122 436226
rect 471178 436170 471248 436226
rect 470928 436102 471248 436170
rect 470928 436046 470998 436102
rect 471054 436046 471122 436102
rect 471178 436046 471248 436102
rect 470928 435978 471248 436046
rect 470928 435922 470998 435978
rect 471054 435922 471122 435978
rect 471178 435922 471248 435978
rect 470928 435888 471248 435922
rect 496938 436350 497558 453922
rect 496938 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 497558 436350
rect 496938 436226 497558 436294
rect 496938 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 497558 436226
rect 496938 436102 497558 436170
rect 496938 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 497558 436102
rect 496938 435978 497558 436046
rect 496938 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 497558 435978
rect 469938 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 470558 424350
rect 469938 424226 470558 424294
rect 469938 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 470558 424226
rect 469938 424102 470558 424170
rect 469938 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 470558 424102
rect 469938 423978 470558 424046
rect 469938 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 470558 423978
rect 466218 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 466838 400350
rect 466218 400226 466838 400294
rect 466218 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 466838 400226
rect 466218 400102 466838 400170
rect 466218 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 466838 400102
rect 466218 399978 466838 400046
rect 466218 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 466838 399978
rect 361228 395220 361284 395230
rect 361228 393876 361284 395164
rect 361228 393810 361284 393820
rect 365148 395108 365204 395118
rect 365148 393876 365204 395052
rect 365148 393810 365204 393820
rect 379820 395108 379876 395118
rect 364476 393316 364532 393326
rect 364476 392698 364532 393260
rect 379820 392868 379876 395052
rect 463036 394660 463092 394670
rect 463036 394100 463092 394604
rect 463036 394034 463092 394044
rect 463708 394660 463764 394670
rect 393148 393316 393204 393326
rect 393148 393092 393204 393260
rect 393148 393026 393204 393036
rect 463708 393092 463764 394604
rect 466218 394566 466838 399922
rect 466956 408548 467012 408558
rect 463708 393026 463764 393036
rect 379820 392802 379876 392812
rect 466956 392868 467012 408492
rect 469938 406350 470558 423922
rect 486288 424350 486608 424384
rect 486288 424294 486358 424350
rect 486414 424294 486482 424350
rect 486538 424294 486608 424350
rect 486288 424226 486608 424294
rect 486288 424170 486358 424226
rect 486414 424170 486482 424226
rect 486538 424170 486608 424226
rect 486288 424102 486608 424170
rect 486288 424046 486358 424102
rect 486414 424046 486482 424102
rect 486538 424046 486608 424102
rect 486288 423978 486608 424046
rect 486288 423922 486358 423978
rect 486414 423922 486482 423978
rect 486538 423922 486608 423978
rect 486288 423888 486608 423922
rect 470928 418350 471248 418384
rect 470928 418294 470998 418350
rect 471054 418294 471122 418350
rect 471178 418294 471248 418350
rect 470928 418226 471248 418294
rect 470928 418170 470998 418226
rect 471054 418170 471122 418226
rect 471178 418170 471248 418226
rect 470928 418102 471248 418170
rect 470928 418046 470998 418102
rect 471054 418046 471122 418102
rect 471178 418046 471248 418102
rect 470928 417978 471248 418046
rect 470928 417922 470998 417978
rect 471054 417922 471122 417978
rect 471178 417922 471248 417978
rect 470928 417888 471248 417922
rect 496938 418350 497558 435922
rect 496938 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 497558 418350
rect 496938 418226 497558 418294
rect 496938 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 497558 418226
rect 496938 418102 497558 418170
rect 496938 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 497558 418102
rect 496938 417978 497558 418046
rect 496938 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 497558 417978
rect 496412 407652 496468 407662
rect 496412 407098 496468 407596
rect 496412 407032 496468 407042
rect 469938 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 470558 406350
rect 469938 406226 470558 406294
rect 469938 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 470558 406226
rect 469938 406102 470558 406170
rect 469938 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 470558 406102
rect 469938 405978 470558 406046
rect 469938 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 470558 405978
rect 469938 394566 470558 405922
rect 490588 406756 490644 406766
rect 490588 395578 490644 406700
rect 490588 395512 490644 395522
rect 496938 400350 497558 417922
rect 496938 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 497558 400350
rect 496938 400226 497558 400294
rect 496938 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 497558 400226
rect 496938 400102 497558 400170
rect 496938 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 497558 400102
rect 496938 399978 497558 400046
rect 496938 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 497558 399978
rect 476924 394772 476980 394782
rect 476924 394212 476980 394716
rect 496938 394566 497558 399922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 568350 501278 585922
rect 500658 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 501278 568350
rect 500658 568226 501278 568294
rect 500658 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 501278 568226
rect 500658 568102 501278 568170
rect 500658 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 501278 568102
rect 500658 567978 501278 568046
rect 500658 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 501278 567978
rect 500658 550350 501278 567922
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 501648 562350 501968 562384
rect 501648 562294 501718 562350
rect 501774 562294 501842 562350
rect 501898 562294 501968 562350
rect 501648 562226 501968 562294
rect 501648 562170 501718 562226
rect 501774 562170 501842 562226
rect 501898 562170 501968 562226
rect 501648 562102 501968 562170
rect 501648 562046 501718 562102
rect 501774 562046 501842 562102
rect 501898 562046 501968 562102
rect 501648 561978 501968 562046
rect 501648 561922 501718 561978
rect 501774 561922 501842 561978
rect 501898 561922 501968 561978
rect 501648 561888 501968 561922
rect 527658 562350 528278 579922
rect 527658 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 528278 562350
rect 527658 562226 528278 562294
rect 527658 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 528278 562226
rect 527658 562102 528278 562170
rect 527658 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 528278 562102
rect 527658 561978 528278 562046
rect 527658 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 528278 561978
rect 500658 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 501278 550350
rect 500658 550226 501278 550294
rect 500658 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 501278 550226
rect 500658 550102 501278 550170
rect 500658 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 501278 550102
rect 500658 549978 501278 550046
rect 500658 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 501278 549978
rect 500658 532350 501278 549922
rect 517008 550350 517328 550384
rect 517008 550294 517078 550350
rect 517134 550294 517202 550350
rect 517258 550294 517328 550350
rect 517008 550226 517328 550294
rect 517008 550170 517078 550226
rect 517134 550170 517202 550226
rect 517258 550170 517328 550226
rect 517008 550102 517328 550170
rect 517008 550046 517078 550102
rect 517134 550046 517202 550102
rect 517258 550046 517328 550102
rect 517008 549978 517328 550046
rect 517008 549922 517078 549978
rect 517134 549922 517202 549978
rect 517258 549922 517328 549978
rect 517008 549888 517328 549922
rect 501648 544350 501968 544384
rect 501648 544294 501718 544350
rect 501774 544294 501842 544350
rect 501898 544294 501968 544350
rect 501648 544226 501968 544294
rect 501648 544170 501718 544226
rect 501774 544170 501842 544226
rect 501898 544170 501968 544226
rect 501648 544102 501968 544170
rect 501648 544046 501718 544102
rect 501774 544046 501842 544102
rect 501898 544046 501968 544102
rect 501648 543978 501968 544046
rect 501648 543922 501718 543978
rect 501774 543922 501842 543978
rect 501898 543922 501968 543978
rect 501648 543888 501968 543922
rect 527658 544350 528278 561922
rect 527658 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 528278 544350
rect 527658 544226 528278 544294
rect 527658 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 528278 544226
rect 527658 544102 528278 544170
rect 527658 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 528278 544102
rect 527658 543978 528278 544046
rect 527658 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 528278 543978
rect 500658 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 501278 532350
rect 500658 532226 501278 532294
rect 500658 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 501278 532226
rect 500658 532102 501278 532170
rect 500658 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 501278 532102
rect 500658 531978 501278 532046
rect 500658 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 501278 531978
rect 500658 514350 501278 531922
rect 517008 532350 517328 532384
rect 517008 532294 517078 532350
rect 517134 532294 517202 532350
rect 517258 532294 517328 532350
rect 517008 532226 517328 532294
rect 517008 532170 517078 532226
rect 517134 532170 517202 532226
rect 517258 532170 517328 532226
rect 517008 532102 517328 532170
rect 517008 532046 517078 532102
rect 517134 532046 517202 532102
rect 517258 532046 517328 532102
rect 517008 531978 517328 532046
rect 517008 531922 517078 531978
rect 517134 531922 517202 531978
rect 517258 531922 517328 531978
rect 517008 531888 517328 531922
rect 501648 526350 501968 526384
rect 501648 526294 501718 526350
rect 501774 526294 501842 526350
rect 501898 526294 501968 526350
rect 501648 526226 501968 526294
rect 501648 526170 501718 526226
rect 501774 526170 501842 526226
rect 501898 526170 501968 526226
rect 501648 526102 501968 526170
rect 501648 526046 501718 526102
rect 501774 526046 501842 526102
rect 501898 526046 501968 526102
rect 501648 525978 501968 526046
rect 501648 525922 501718 525978
rect 501774 525922 501842 525978
rect 501898 525922 501968 525978
rect 501648 525888 501968 525922
rect 527658 526350 528278 543922
rect 527658 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 528278 526350
rect 527658 526226 528278 526294
rect 527658 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 528278 526226
rect 527658 526102 528278 526170
rect 527658 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 528278 526102
rect 527658 525978 528278 526046
rect 527658 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 528278 525978
rect 500658 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 501278 514350
rect 500658 514226 501278 514294
rect 500658 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 501278 514226
rect 500658 514102 501278 514170
rect 500658 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 501278 514102
rect 500658 513978 501278 514046
rect 500658 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 501278 513978
rect 500658 496350 501278 513922
rect 517008 514350 517328 514384
rect 517008 514294 517078 514350
rect 517134 514294 517202 514350
rect 517258 514294 517328 514350
rect 517008 514226 517328 514294
rect 517008 514170 517078 514226
rect 517134 514170 517202 514226
rect 517258 514170 517328 514226
rect 517008 514102 517328 514170
rect 517008 514046 517078 514102
rect 517134 514046 517202 514102
rect 517258 514046 517328 514102
rect 517008 513978 517328 514046
rect 517008 513922 517078 513978
rect 517134 513922 517202 513978
rect 517258 513922 517328 513978
rect 517008 513888 517328 513922
rect 501648 508350 501968 508384
rect 501648 508294 501718 508350
rect 501774 508294 501842 508350
rect 501898 508294 501968 508350
rect 501648 508226 501968 508294
rect 501648 508170 501718 508226
rect 501774 508170 501842 508226
rect 501898 508170 501968 508226
rect 501648 508102 501968 508170
rect 501648 508046 501718 508102
rect 501774 508046 501842 508102
rect 501898 508046 501968 508102
rect 501648 507978 501968 508046
rect 501648 507922 501718 507978
rect 501774 507922 501842 507978
rect 501898 507922 501968 507978
rect 501648 507888 501968 507922
rect 527658 508350 528278 525922
rect 527658 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 528278 508350
rect 527658 508226 528278 508294
rect 527658 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 528278 508226
rect 527658 508102 528278 508170
rect 527658 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 528278 508102
rect 527658 507978 528278 508046
rect 527658 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 528278 507978
rect 500658 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 501278 496350
rect 500658 496226 501278 496294
rect 500658 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 501278 496226
rect 500658 496102 501278 496170
rect 500658 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 501278 496102
rect 500658 495978 501278 496046
rect 500658 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 501278 495978
rect 500658 478350 501278 495922
rect 517008 496350 517328 496384
rect 517008 496294 517078 496350
rect 517134 496294 517202 496350
rect 517258 496294 517328 496350
rect 517008 496226 517328 496294
rect 517008 496170 517078 496226
rect 517134 496170 517202 496226
rect 517258 496170 517328 496226
rect 517008 496102 517328 496170
rect 517008 496046 517078 496102
rect 517134 496046 517202 496102
rect 517258 496046 517328 496102
rect 517008 495978 517328 496046
rect 517008 495922 517078 495978
rect 517134 495922 517202 495978
rect 517258 495922 517328 495978
rect 517008 495888 517328 495922
rect 501648 490350 501968 490384
rect 501648 490294 501718 490350
rect 501774 490294 501842 490350
rect 501898 490294 501968 490350
rect 501648 490226 501968 490294
rect 501648 490170 501718 490226
rect 501774 490170 501842 490226
rect 501898 490170 501968 490226
rect 501648 490102 501968 490170
rect 501648 490046 501718 490102
rect 501774 490046 501842 490102
rect 501898 490046 501968 490102
rect 501648 489978 501968 490046
rect 501648 489922 501718 489978
rect 501774 489922 501842 489978
rect 501898 489922 501968 489978
rect 501648 489888 501968 489922
rect 527658 490350 528278 507922
rect 527658 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 528278 490350
rect 527658 490226 528278 490294
rect 527658 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 528278 490226
rect 527658 490102 528278 490170
rect 527658 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 528278 490102
rect 527658 489978 528278 490046
rect 527658 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 528278 489978
rect 500658 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 501278 478350
rect 500658 478226 501278 478294
rect 500658 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 501278 478226
rect 500658 478102 501278 478170
rect 500658 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 501278 478102
rect 500658 477978 501278 478046
rect 500658 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 501278 477978
rect 500658 460350 501278 477922
rect 517008 478350 517328 478384
rect 517008 478294 517078 478350
rect 517134 478294 517202 478350
rect 517258 478294 517328 478350
rect 517008 478226 517328 478294
rect 517008 478170 517078 478226
rect 517134 478170 517202 478226
rect 517258 478170 517328 478226
rect 517008 478102 517328 478170
rect 517008 478046 517078 478102
rect 517134 478046 517202 478102
rect 517258 478046 517328 478102
rect 517008 477978 517328 478046
rect 517008 477922 517078 477978
rect 517134 477922 517202 477978
rect 517258 477922 517328 477978
rect 517008 477888 517328 477922
rect 501648 472350 501968 472384
rect 501648 472294 501718 472350
rect 501774 472294 501842 472350
rect 501898 472294 501968 472350
rect 501648 472226 501968 472294
rect 501648 472170 501718 472226
rect 501774 472170 501842 472226
rect 501898 472170 501968 472226
rect 501648 472102 501968 472170
rect 501648 472046 501718 472102
rect 501774 472046 501842 472102
rect 501898 472046 501968 472102
rect 501648 471978 501968 472046
rect 501648 471922 501718 471978
rect 501774 471922 501842 471978
rect 501898 471922 501968 471978
rect 501648 471888 501968 471922
rect 527658 472350 528278 489922
rect 527658 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 528278 472350
rect 527658 472226 528278 472294
rect 527658 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 528278 472226
rect 527658 472102 528278 472170
rect 527658 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 528278 472102
rect 527658 471978 528278 472046
rect 527658 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 528278 471978
rect 500658 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 501278 460350
rect 500658 460226 501278 460294
rect 500658 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 501278 460226
rect 500658 460102 501278 460170
rect 500658 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 501278 460102
rect 500658 459978 501278 460046
rect 500658 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 501278 459978
rect 500658 442350 501278 459922
rect 517008 460350 517328 460384
rect 517008 460294 517078 460350
rect 517134 460294 517202 460350
rect 517258 460294 517328 460350
rect 517008 460226 517328 460294
rect 517008 460170 517078 460226
rect 517134 460170 517202 460226
rect 517258 460170 517328 460226
rect 517008 460102 517328 460170
rect 517008 460046 517078 460102
rect 517134 460046 517202 460102
rect 517258 460046 517328 460102
rect 517008 459978 517328 460046
rect 517008 459922 517078 459978
rect 517134 459922 517202 459978
rect 517258 459922 517328 459978
rect 517008 459888 517328 459922
rect 501648 454350 501968 454384
rect 501648 454294 501718 454350
rect 501774 454294 501842 454350
rect 501898 454294 501968 454350
rect 501648 454226 501968 454294
rect 501648 454170 501718 454226
rect 501774 454170 501842 454226
rect 501898 454170 501968 454226
rect 501648 454102 501968 454170
rect 501648 454046 501718 454102
rect 501774 454046 501842 454102
rect 501898 454046 501968 454102
rect 501648 453978 501968 454046
rect 501648 453922 501718 453978
rect 501774 453922 501842 453978
rect 501898 453922 501968 453978
rect 501648 453888 501968 453922
rect 527658 454350 528278 471922
rect 527658 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 528278 454350
rect 527658 454226 528278 454294
rect 527658 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 528278 454226
rect 527658 454102 528278 454170
rect 527658 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 528278 454102
rect 527658 453978 528278 454046
rect 527658 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 528278 453978
rect 500658 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 501278 442350
rect 500658 442226 501278 442294
rect 500658 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 501278 442226
rect 500658 442102 501278 442170
rect 500658 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 501278 442102
rect 500658 441978 501278 442046
rect 500658 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 501278 441978
rect 500658 424350 501278 441922
rect 517008 442350 517328 442384
rect 517008 442294 517078 442350
rect 517134 442294 517202 442350
rect 517258 442294 517328 442350
rect 517008 442226 517328 442294
rect 517008 442170 517078 442226
rect 517134 442170 517202 442226
rect 517258 442170 517328 442226
rect 517008 442102 517328 442170
rect 517008 442046 517078 442102
rect 517134 442046 517202 442102
rect 517258 442046 517328 442102
rect 517008 441978 517328 442046
rect 517008 441922 517078 441978
rect 517134 441922 517202 441978
rect 517258 441922 517328 441978
rect 517008 441888 517328 441922
rect 501648 436350 501968 436384
rect 501648 436294 501718 436350
rect 501774 436294 501842 436350
rect 501898 436294 501968 436350
rect 501648 436226 501968 436294
rect 501648 436170 501718 436226
rect 501774 436170 501842 436226
rect 501898 436170 501968 436226
rect 501648 436102 501968 436170
rect 501648 436046 501718 436102
rect 501774 436046 501842 436102
rect 501898 436046 501968 436102
rect 501648 435978 501968 436046
rect 501648 435922 501718 435978
rect 501774 435922 501842 435978
rect 501898 435922 501968 435978
rect 501648 435888 501968 435922
rect 527658 436350 528278 453922
rect 527658 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 528278 436350
rect 527658 436226 528278 436294
rect 527658 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 528278 436226
rect 527658 436102 528278 436170
rect 527658 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 528278 436102
rect 527658 435978 528278 436046
rect 527658 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 528278 435978
rect 500658 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 501278 424350
rect 500658 424226 501278 424294
rect 500658 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 501278 424226
rect 500658 424102 501278 424170
rect 500658 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 501278 424102
rect 500658 423978 501278 424046
rect 500658 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 501278 423978
rect 500658 406350 501278 423922
rect 517008 424350 517328 424384
rect 517008 424294 517078 424350
rect 517134 424294 517202 424350
rect 517258 424294 517328 424350
rect 517008 424226 517328 424294
rect 517008 424170 517078 424226
rect 517134 424170 517202 424226
rect 517258 424170 517328 424226
rect 517008 424102 517328 424170
rect 517008 424046 517078 424102
rect 517134 424046 517202 424102
rect 517258 424046 517328 424102
rect 517008 423978 517328 424046
rect 517008 423922 517078 423978
rect 517134 423922 517202 423978
rect 517258 423922 517328 423978
rect 517008 423888 517328 423922
rect 501648 418350 501968 418384
rect 501648 418294 501718 418350
rect 501774 418294 501842 418350
rect 501898 418294 501968 418350
rect 501648 418226 501968 418294
rect 501648 418170 501718 418226
rect 501774 418170 501842 418226
rect 501898 418170 501968 418226
rect 501648 418102 501968 418170
rect 501648 418046 501718 418102
rect 501774 418046 501842 418102
rect 501898 418046 501968 418102
rect 501648 417978 501968 418046
rect 501648 417922 501718 417978
rect 501774 417922 501842 417978
rect 501898 417922 501968 417978
rect 501648 417888 501968 417922
rect 527658 418350 528278 435922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 568350 531998 585922
rect 531378 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 531998 568350
rect 531378 568226 531998 568294
rect 531378 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 531998 568226
rect 531378 568102 531998 568170
rect 531378 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 531998 568102
rect 531378 567978 531998 568046
rect 531378 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 531998 567978
rect 531378 550350 531998 567922
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 558378 580350 558998 596784
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 532924 565124 532980 565134
rect 531378 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 531998 550350
rect 531378 550226 531998 550294
rect 531378 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 531998 550226
rect 531378 550102 531998 550170
rect 531378 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 531998 550102
rect 531378 549978 531998 550046
rect 531378 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 531998 549978
rect 531378 532350 531998 549922
rect 531378 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 531998 532350
rect 531378 532226 531998 532294
rect 531378 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 531998 532226
rect 531378 532102 531998 532170
rect 531378 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 531998 532102
rect 531378 531978 531998 532046
rect 531378 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 531998 531978
rect 531378 514350 531998 531922
rect 531378 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 531998 514350
rect 531378 514226 531998 514294
rect 531378 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 531998 514226
rect 531378 514102 531998 514170
rect 531378 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 531998 514102
rect 531378 513978 531998 514046
rect 531378 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 531998 513978
rect 531378 496350 531998 513922
rect 531378 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 531998 496350
rect 531378 496226 531998 496294
rect 531378 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 531998 496226
rect 531378 496102 531998 496170
rect 531378 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 531998 496102
rect 531378 495978 531998 496046
rect 531378 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 531998 495978
rect 531378 478350 531998 495922
rect 531378 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 531998 478350
rect 531378 478226 531998 478294
rect 531378 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 531998 478226
rect 531378 478102 531998 478170
rect 531378 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 531998 478102
rect 531378 477978 531998 478046
rect 531378 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 531998 477978
rect 531378 460350 531998 477922
rect 531378 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 531998 460350
rect 531378 460226 531998 460294
rect 531378 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 531998 460226
rect 531378 460102 531998 460170
rect 531378 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 531998 460102
rect 531378 459978 531998 460046
rect 531378 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 531998 459978
rect 531378 442350 531998 459922
rect 531378 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 531998 442350
rect 531378 442226 531998 442294
rect 531378 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 531998 442226
rect 531378 442102 531998 442170
rect 531378 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 531998 442102
rect 531378 441978 531998 442046
rect 531378 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 531998 441978
rect 529228 428708 529284 428718
rect 529228 428614 529284 428642
rect 527658 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 528278 418350
rect 527658 418226 528278 418294
rect 527658 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 528278 418226
rect 527658 418102 528278 418170
rect 527658 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 528278 418102
rect 527658 417978 528278 418046
rect 527658 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 528278 417978
rect 522172 407540 522228 407550
rect 522172 406918 522228 407484
rect 522172 406852 522228 406862
rect 527324 407540 527380 407550
rect 527324 406738 527380 407484
rect 527324 406672 527380 406682
rect 500658 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 501278 406350
rect 500658 406226 501278 406294
rect 500658 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 501278 406226
rect 500658 406102 501278 406170
rect 500658 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 501278 406102
rect 500658 405978 501278 406046
rect 500658 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 501278 405978
rect 500658 394566 501278 405922
rect 527658 400350 528278 417922
rect 527658 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 528278 400350
rect 527658 400226 528278 400294
rect 527658 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 528278 400226
rect 527658 400102 528278 400170
rect 527658 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 528278 400102
rect 527658 399978 528278 400046
rect 527658 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 528278 399978
rect 525532 395038 525588 395048
rect 525532 394930 525588 394940
rect 511644 394772 511700 394782
rect 511644 394436 511700 394716
rect 527658 394566 528278 399922
rect 531378 424350 531998 441922
rect 531378 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 531998 424350
rect 531378 424226 531998 424294
rect 531378 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 531998 424226
rect 531378 424102 531998 424170
rect 531378 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 531998 424102
rect 531378 423978 531998 424046
rect 531378 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 531998 423978
rect 531378 406350 531998 423922
rect 532700 555716 532756 555726
rect 532700 409438 532756 555660
rect 532700 409372 532756 409382
rect 532812 442820 532868 442830
rect 532812 407458 532868 442764
rect 532812 407392 532868 407402
rect 531378 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 531998 406350
rect 531378 406226 531998 406294
rect 531378 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 531998 406226
rect 531378 406102 531998 406170
rect 531378 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 531998 406102
rect 531378 405978 531998 406046
rect 531378 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 531998 405978
rect 531378 394566 531998 405922
rect 532924 405478 532980 565068
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 535948 560420 536004 560430
rect 532924 405412 532980 405422
rect 534268 475748 534324 475758
rect 534268 398998 534324 475692
rect 535948 405658 536004 560364
rect 537628 551012 537684 551022
rect 537628 409258 537684 550956
rect 558378 544350 558998 561922
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 543452 535780 543508 535790
rect 541772 496132 541828 496142
rect 537628 409192 537684 409202
rect 540092 416836 540148 416846
rect 535948 405592 536004 405602
rect 540092 404218 540148 416780
rect 541772 404398 541828 496076
rect 541772 404332 541828 404342
rect 540092 404152 540148 404162
rect 543452 402778 543508 535724
rect 543452 402712 543508 402722
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 558378 472350 558998 489922
rect 558378 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 558998 472350
rect 558378 472226 558998 472294
rect 558378 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 558998 472226
rect 558378 472102 558998 472170
rect 558378 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 558998 472102
rect 558378 471978 558998 472046
rect 558378 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 558998 471978
rect 558378 454350 558998 471922
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 534268 398932 534324 398942
rect 558378 400350 558998 417922
rect 558378 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 558998 400350
rect 558378 400226 558998 400294
rect 558378 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 558998 400226
rect 558378 400102 558998 400170
rect 558378 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 558998 400102
rect 558378 399978 558998 400046
rect 558378 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 558998 399978
rect 546252 397378 546308 397388
rect 546252 396900 546308 397322
rect 546252 396834 546308 396844
rect 553196 396838 553252 396848
rect 553196 396676 553252 396782
rect 553196 396610 553252 396620
rect 558378 394566 558998 399922
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 562098 550350 562718 567922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 562098 532350 562718 549922
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 562098 478350 562718 495922
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 562098 460350 562718 477922
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 584668 590212 584724 590222
rect 584668 409798 584724 590156
rect 584668 409732 584724 409742
rect 589098 580350 589718 596784
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 589098 562350 589718 579922
rect 590492 588644 590548 588654
rect 590492 573748 590548 588588
rect 590492 573682 590548 573692
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 590604 567924 590660 567934
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 562098 394566 562718 405922
rect 581756 406644 581812 406654
rect 574028 397198 574084 397208
rect 574028 396900 574084 397142
rect 574028 396834 574084 396844
rect 580972 397018 581028 397028
rect 580972 396788 581028 396962
rect 580972 396722 581028 396732
rect 567084 396658 567140 396668
rect 567084 396564 567140 396602
rect 567084 396498 567140 396508
rect 511644 394370 511700 394380
rect 476924 394146 476980 394156
rect 466956 392802 467012 392812
rect 364476 392632 364532 392642
rect 374808 388350 375128 388384
rect 374808 388294 374878 388350
rect 374934 388294 375002 388350
rect 375058 388294 375128 388350
rect 374808 388226 375128 388294
rect 374808 388170 374878 388226
rect 374934 388170 375002 388226
rect 375058 388170 375128 388226
rect 374808 388102 375128 388170
rect 374808 388046 374878 388102
rect 374934 388046 375002 388102
rect 375058 388046 375128 388102
rect 374808 387978 375128 388046
rect 374808 387922 374878 387978
rect 374934 387922 375002 387978
rect 375058 387922 375128 387978
rect 374808 387888 375128 387922
rect 405528 388350 405848 388384
rect 405528 388294 405598 388350
rect 405654 388294 405722 388350
rect 405778 388294 405848 388350
rect 405528 388226 405848 388294
rect 405528 388170 405598 388226
rect 405654 388170 405722 388226
rect 405778 388170 405848 388226
rect 405528 388102 405848 388170
rect 405528 388046 405598 388102
rect 405654 388046 405722 388102
rect 405778 388046 405848 388102
rect 405528 387978 405848 388046
rect 405528 387922 405598 387978
rect 405654 387922 405722 387978
rect 405778 387922 405848 387978
rect 405528 387888 405848 387922
rect 436248 388350 436568 388384
rect 436248 388294 436318 388350
rect 436374 388294 436442 388350
rect 436498 388294 436568 388350
rect 436248 388226 436568 388294
rect 436248 388170 436318 388226
rect 436374 388170 436442 388226
rect 436498 388170 436568 388226
rect 436248 388102 436568 388170
rect 436248 388046 436318 388102
rect 436374 388046 436442 388102
rect 436498 388046 436568 388102
rect 436248 387978 436568 388046
rect 436248 387922 436318 387978
rect 436374 387922 436442 387978
rect 436498 387922 436568 387978
rect 436248 387888 436568 387922
rect 466968 388350 467288 388384
rect 466968 388294 467038 388350
rect 467094 388294 467162 388350
rect 467218 388294 467288 388350
rect 466968 388226 467288 388294
rect 466968 388170 467038 388226
rect 467094 388170 467162 388226
rect 467218 388170 467288 388226
rect 466968 388102 467288 388170
rect 466968 388046 467038 388102
rect 467094 388046 467162 388102
rect 467218 388046 467288 388102
rect 466968 387978 467288 388046
rect 466968 387922 467038 387978
rect 467094 387922 467162 387978
rect 467218 387922 467288 387978
rect 466968 387888 467288 387922
rect 497688 388350 498008 388384
rect 497688 388294 497758 388350
rect 497814 388294 497882 388350
rect 497938 388294 498008 388350
rect 497688 388226 498008 388294
rect 497688 388170 497758 388226
rect 497814 388170 497882 388226
rect 497938 388170 498008 388226
rect 497688 388102 498008 388170
rect 497688 388046 497758 388102
rect 497814 388046 497882 388102
rect 497938 388046 498008 388102
rect 497688 387978 498008 388046
rect 497688 387922 497758 387978
rect 497814 387922 497882 387978
rect 497938 387922 498008 387978
rect 497688 387888 498008 387922
rect 528408 388350 528728 388384
rect 528408 388294 528478 388350
rect 528534 388294 528602 388350
rect 528658 388294 528728 388350
rect 528408 388226 528728 388294
rect 528408 388170 528478 388226
rect 528534 388170 528602 388226
rect 528658 388170 528728 388226
rect 528408 388102 528728 388170
rect 528408 388046 528478 388102
rect 528534 388046 528602 388102
rect 528658 388046 528728 388102
rect 528408 387978 528728 388046
rect 528408 387922 528478 387978
rect 528534 387922 528602 387978
rect 528658 387922 528728 387978
rect 528408 387888 528728 387922
rect 559128 388350 559448 388384
rect 559128 388294 559198 388350
rect 559254 388294 559322 388350
rect 559378 388294 559448 388350
rect 559128 388226 559448 388294
rect 559128 388170 559198 388226
rect 559254 388170 559322 388226
rect 559378 388170 559448 388226
rect 559128 388102 559448 388170
rect 559128 388046 559198 388102
rect 559254 388046 559322 388102
rect 559378 388046 559448 388102
rect 559128 387978 559448 388046
rect 559128 387922 559198 387978
rect 559254 387922 559322 387978
rect 559378 387922 559448 387978
rect 559128 387888 559448 387922
rect 359448 382350 359768 382384
rect 359448 382294 359518 382350
rect 359574 382294 359642 382350
rect 359698 382294 359768 382350
rect 359448 382226 359768 382294
rect 359448 382170 359518 382226
rect 359574 382170 359642 382226
rect 359698 382170 359768 382226
rect 359448 382102 359768 382170
rect 359448 382046 359518 382102
rect 359574 382046 359642 382102
rect 359698 382046 359768 382102
rect 359448 381978 359768 382046
rect 359448 381922 359518 381978
rect 359574 381922 359642 381978
rect 359698 381922 359768 381978
rect 359448 381888 359768 381922
rect 390168 382350 390488 382384
rect 390168 382294 390238 382350
rect 390294 382294 390362 382350
rect 390418 382294 390488 382350
rect 390168 382226 390488 382294
rect 390168 382170 390238 382226
rect 390294 382170 390362 382226
rect 390418 382170 390488 382226
rect 390168 382102 390488 382170
rect 390168 382046 390238 382102
rect 390294 382046 390362 382102
rect 390418 382046 390488 382102
rect 390168 381978 390488 382046
rect 390168 381922 390238 381978
rect 390294 381922 390362 381978
rect 390418 381922 390488 381978
rect 390168 381888 390488 381922
rect 420888 382350 421208 382384
rect 420888 382294 420958 382350
rect 421014 382294 421082 382350
rect 421138 382294 421208 382350
rect 420888 382226 421208 382294
rect 420888 382170 420958 382226
rect 421014 382170 421082 382226
rect 421138 382170 421208 382226
rect 420888 382102 421208 382170
rect 420888 382046 420958 382102
rect 421014 382046 421082 382102
rect 421138 382046 421208 382102
rect 420888 381978 421208 382046
rect 420888 381922 420958 381978
rect 421014 381922 421082 381978
rect 421138 381922 421208 381978
rect 420888 381888 421208 381922
rect 451608 382350 451928 382384
rect 451608 382294 451678 382350
rect 451734 382294 451802 382350
rect 451858 382294 451928 382350
rect 451608 382226 451928 382294
rect 451608 382170 451678 382226
rect 451734 382170 451802 382226
rect 451858 382170 451928 382226
rect 451608 382102 451928 382170
rect 451608 382046 451678 382102
rect 451734 382046 451802 382102
rect 451858 382046 451928 382102
rect 451608 381978 451928 382046
rect 451608 381922 451678 381978
rect 451734 381922 451802 381978
rect 451858 381922 451928 381978
rect 451608 381888 451928 381922
rect 482328 382350 482648 382384
rect 482328 382294 482398 382350
rect 482454 382294 482522 382350
rect 482578 382294 482648 382350
rect 482328 382226 482648 382294
rect 482328 382170 482398 382226
rect 482454 382170 482522 382226
rect 482578 382170 482648 382226
rect 482328 382102 482648 382170
rect 482328 382046 482398 382102
rect 482454 382046 482522 382102
rect 482578 382046 482648 382102
rect 482328 381978 482648 382046
rect 482328 381922 482398 381978
rect 482454 381922 482522 381978
rect 482578 381922 482648 381978
rect 482328 381888 482648 381922
rect 513048 382350 513368 382384
rect 513048 382294 513118 382350
rect 513174 382294 513242 382350
rect 513298 382294 513368 382350
rect 513048 382226 513368 382294
rect 513048 382170 513118 382226
rect 513174 382170 513242 382226
rect 513298 382170 513368 382226
rect 513048 382102 513368 382170
rect 513048 382046 513118 382102
rect 513174 382046 513242 382102
rect 513298 382046 513368 382102
rect 513048 381978 513368 382046
rect 513048 381922 513118 381978
rect 513174 381922 513242 381978
rect 513298 381922 513368 381978
rect 513048 381888 513368 381922
rect 543768 382350 544088 382384
rect 543768 382294 543838 382350
rect 543894 382294 543962 382350
rect 544018 382294 544088 382350
rect 543768 382226 544088 382294
rect 543768 382170 543838 382226
rect 543894 382170 543962 382226
rect 544018 382170 544088 382226
rect 543768 382102 544088 382170
rect 543768 382046 543838 382102
rect 543894 382046 543962 382102
rect 544018 382046 544088 382102
rect 543768 381978 544088 382046
rect 543768 381922 543838 381978
rect 543894 381922 543962 381978
rect 544018 381922 544088 381978
rect 543768 381888 544088 381922
rect 574488 382350 574808 382384
rect 574488 382294 574558 382350
rect 574614 382294 574682 382350
rect 574738 382294 574808 382350
rect 574488 382226 574808 382294
rect 574488 382170 574558 382226
rect 574614 382170 574682 382226
rect 574738 382170 574808 382226
rect 574488 382102 574808 382170
rect 574488 382046 574558 382102
rect 574614 382046 574682 382102
rect 574738 382046 574808 382102
rect 574488 381978 574808 382046
rect 574488 381922 574558 381978
rect 574614 381922 574682 381978
rect 574738 381922 574808 381978
rect 574488 381888 574808 381922
rect 374808 370350 375128 370384
rect 374808 370294 374878 370350
rect 374934 370294 375002 370350
rect 375058 370294 375128 370350
rect 374808 370226 375128 370294
rect 374808 370170 374878 370226
rect 374934 370170 375002 370226
rect 375058 370170 375128 370226
rect 374808 370102 375128 370170
rect 374808 370046 374878 370102
rect 374934 370046 375002 370102
rect 375058 370046 375128 370102
rect 374808 369978 375128 370046
rect 374808 369922 374878 369978
rect 374934 369922 375002 369978
rect 375058 369922 375128 369978
rect 374808 369888 375128 369922
rect 405528 370350 405848 370384
rect 405528 370294 405598 370350
rect 405654 370294 405722 370350
rect 405778 370294 405848 370350
rect 405528 370226 405848 370294
rect 405528 370170 405598 370226
rect 405654 370170 405722 370226
rect 405778 370170 405848 370226
rect 405528 370102 405848 370170
rect 405528 370046 405598 370102
rect 405654 370046 405722 370102
rect 405778 370046 405848 370102
rect 405528 369978 405848 370046
rect 405528 369922 405598 369978
rect 405654 369922 405722 369978
rect 405778 369922 405848 369978
rect 405528 369888 405848 369922
rect 436248 370350 436568 370384
rect 436248 370294 436318 370350
rect 436374 370294 436442 370350
rect 436498 370294 436568 370350
rect 436248 370226 436568 370294
rect 436248 370170 436318 370226
rect 436374 370170 436442 370226
rect 436498 370170 436568 370226
rect 436248 370102 436568 370170
rect 436248 370046 436318 370102
rect 436374 370046 436442 370102
rect 436498 370046 436568 370102
rect 436248 369978 436568 370046
rect 436248 369922 436318 369978
rect 436374 369922 436442 369978
rect 436498 369922 436568 369978
rect 436248 369888 436568 369922
rect 466968 370350 467288 370384
rect 466968 370294 467038 370350
rect 467094 370294 467162 370350
rect 467218 370294 467288 370350
rect 466968 370226 467288 370294
rect 466968 370170 467038 370226
rect 467094 370170 467162 370226
rect 467218 370170 467288 370226
rect 466968 370102 467288 370170
rect 466968 370046 467038 370102
rect 467094 370046 467162 370102
rect 467218 370046 467288 370102
rect 466968 369978 467288 370046
rect 466968 369922 467038 369978
rect 467094 369922 467162 369978
rect 467218 369922 467288 369978
rect 466968 369888 467288 369922
rect 497688 370350 498008 370384
rect 497688 370294 497758 370350
rect 497814 370294 497882 370350
rect 497938 370294 498008 370350
rect 497688 370226 498008 370294
rect 497688 370170 497758 370226
rect 497814 370170 497882 370226
rect 497938 370170 498008 370226
rect 497688 370102 498008 370170
rect 497688 370046 497758 370102
rect 497814 370046 497882 370102
rect 497938 370046 498008 370102
rect 497688 369978 498008 370046
rect 497688 369922 497758 369978
rect 497814 369922 497882 369978
rect 497938 369922 498008 369978
rect 497688 369888 498008 369922
rect 528408 370350 528728 370384
rect 528408 370294 528478 370350
rect 528534 370294 528602 370350
rect 528658 370294 528728 370350
rect 528408 370226 528728 370294
rect 528408 370170 528478 370226
rect 528534 370170 528602 370226
rect 528658 370170 528728 370226
rect 528408 370102 528728 370170
rect 528408 370046 528478 370102
rect 528534 370046 528602 370102
rect 528658 370046 528728 370102
rect 528408 369978 528728 370046
rect 528408 369922 528478 369978
rect 528534 369922 528602 369978
rect 528658 369922 528728 369978
rect 528408 369888 528728 369922
rect 559128 370350 559448 370384
rect 559128 370294 559198 370350
rect 559254 370294 559322 370350
rect 559378 370294 559448 370350
rect 559128 370226 559448 370294
rect 559128 370170 559198 370226
rect 559254 370170 559322 370226
rect 559378 370170 559448 370226
rect 559128 370102 559448 370170
rect 559128 370046 559198 370102
rect 559254 370046 559322 370102
rect 559378 370046 559448 370102
rect 559128 369978 559448 370046
rect 559128 369922 559198 369978
rect 559254 369922 559322 369978
rect 559378 369922 559448 369978
rect 559128 369888 559448 369922
rect 359448 364350 359768 364384
rect 359448 364294 359518 364350
rect 359574 364294 359642 364350
rect 359698 364294 359768 364350
rect 359448 364226 359768 364294
rect 359448 364170 359518 364226
rect 359574 364170 359642 364226
rect 359698 364170 359768 364226
rect 359448 364102 359768 364170
rect 359448 364046 359518 364102
rect 359574 364046 359642 364102
rect 359698 364046 359768 364102
rect 359448 363978 359768 364046
rect 359448 363922 359518 363978
rect 359574 363922 359642 363978
rect 359698 363922 359768 363978
rect 359448 363888 359768 363922
rect 390168 364350 390488 364384
rect 390168 364294 390238 364350
rect 390294 364294 390362 364350
rect 390418 364294 390488 364350
rect 390168 364226 390488 364294
rect 390168 364170 390238 364226
rect 390294 364170 390362 364226
rect 390418 364170 390488 364226
rect 390168 364102 390488 364170
rect 390168 364046 390238 364102
rect 390294 364046 390362 364102
rect 390418 364046 390488 364102
rect 390168 363978 390488 364046
rect 390168 363922 390238 363978
rect 390294 363922 390362 363978
rect 390418 363922 390488 363978
rect 390168 363888 390488 363922
rect 420888 364350 421208 364384
rect 420888 364294 420958 364350
rect 421014 364294 421082 364350
rect 421138 364294 421208 364350
rect 420888 364226 421208 364294
rect 420888 364170 420958 364226
rect 421014 364170 421082 364226
rect 421138 364170 421208 364226
rect 420888 364102 421208 364170
rect 420888 364046 420958 364102
rect 421014 364046 421082 364102
rect 421138 364046 421208 364102
rect 420888 363978 421208 364046
rect 420888 363922 420958 363978
rect 421014 363922 421082 363978
rect 421138 363922 421208 363978
rect 420888 363888 421208 363922
rect 451608 364350 451928 364384
rect 451608 364294 451678 364350
rect 451734 364294 451802 364350
rect 451858 364294 451928 364350
rect 451608 364226 451928 364294
rect 451608 364170 451678 364226
rect 451734 364170 451802 364226
rect 451858 364170 451928 364226
rect 451608 364102 451928 364170
rect 451608 364046 451678 364102
rect 451734 364046 451802 364102
rect 451858 364046 451928 364102
rect 451608 363978 451928 364046
rect 451608 363922 451678 363978
rect 451734 363922 451802 363978
rect 451858 363922 451928 363978
rect 451608 363888 451928 363922
rect 482328 364350 482648 364384
rect 482328 364294 482398 364350
rect 482454 364294 482522 364350
rect 482578 364294 482648 364350
rect 482328 364226 482648 364294
rect 482328 364170 482398 364226
rect 482454 364170 482522 364226
rect 482578 364170 482648 364226
rect 482328 364102 482648 364170
rect 482328 364046 482398 364102
rect 482454 364046 482522 364102
rect 482578 364046 482648 364102
rect 482328 363978 482648 364046
rect 482328 363922 482398 363978
rect 482454 363922 482522 363978
rect 482578 363922 482648 363978
rect 482328 363888 482648 363922
rect 513048 364350 513368 364384
rect 513048 364294 513118 364350
rect 513174 364294 513242 364350
rect 513298 364294 513368 364350
rect 513048 364226 513368 364294
rect 513048 364170 513118 364226
rect 513174 364170 513242 364226
rect 513298 364170 513368 364226
rect 513048 364102 513368 364170
rect 513048 364046 513118 364102
rect 513174 364046 513242 364102
rect 513298 364046 513368 364102
rect 513048 363978 513368 364046
rect 513048 363922 513118 363978
rect 513174 363922 513242 363978
rect 513298 363922 513368 363978
rect 513048 363888 513368 363922
rect 543768 364350 544088 364384
rect 543768 364294 543838 364350
rect 543894 364294 543962 364350
rect 544018 364294 544088 364350
rect 543768 364226 544088 364294
rect 543768 364170 543838 364226
rect 543894 364170 543962 364226
rect 544018 364170 544088 364226
rect 543768 364102 544088 364170
rect 543768 364046 543838 364102
rect 543894 364046 543962 364102
rect 544018 364046 544088 364102
rect 543768 363978 544088 364046
rect 543768 363922 543838 363978
rect 543894 363922 543962 363978
rect 544018 363922 544088 363978
rect 543768 363888 544088 363922
rect 574488 364350 574808 364384
rect 574488 364294 574558 364350
rect 574614 364294 574682 364350
rect 574738 364294 574808 364350
rect 574488 364226 574808 364294
rect 574488 364170 574558 364226
rect 574614 364170 574682 364226
rect 574738 364170 574808 364226
rect 574488 364102 574808 364170
rect 574488 364046 574558 364102
rect 574614 364046 574682 364102
rect 574738 364046 574808 364102
rect 574488 363978 574808 364046
rect 574488 363922 574558 363978
rect 574614 363922 574682 363978
rect 574738 363922 574808 363978
rect 574488 363888 574808 363922
rect 374808 352350 375128 352384
rect 374808 352294 374878 352350
rect 374934 352294 375002 352350
rect 375058 352294 375128 352350
rect 374808 352226 375128 352294
rect 374808 352170 374878 352226
rect 374934 352170 375002 352226
rect 375058 352170 375128 352226
rect 374808 352102 375128 352170
rect 374808 352046 374878 352102
rect 374934 352046 375002 352102
rect 375058 352046 375128 352102
rect 374808 351978 375128 352046
rect 374808 351922 374878 351978
rect 374934 351922 375002 351978
rect 375058 351922 375128 351978
rect 374808 351888 375128 351922
rect 405528 352350 405848 352384
rect 405528 352294 405598 352350
rect 405654 352294 405722 352350
rect 405778 352294 405848 352350
rect 405528 352226 405848 352294
rect 405528 352170 405598 352226
rect 405654 352170 405722 352226
rect 405778 352170 405848 352226
rect 405528 352102 405848 352170
rect 405528 352046 405598 352102
rect 405654 352046 405722 352102
rect 405778 352046 405848 352102
rect 405528 351978 405848 352046
rect 405528 351922 405598 351978
rect 405654 351922 405722 351978
rect 405778 351922 405848 351978
rect 405528 351888 405848 351922
rect 436248 352350 436568 352384
rect 436248 352294 436318 352350
rect 436374 352294 436442 352350
rect 436498 352294 436568 352350
rect 436248 352226 436568 352294
rect 436248 352170 436318 352226
rect 436374 352170 436442 352226
rect 436498 352170 436568 352226
rect 436248 352102 436568 352170
rect 436248 352046 436318 352102
rect 436374 352046 436442 352102
rect 436498 352046 436568 352102
rect 436248 351978 436568 352046
rect 436248 351922 436318 351978
rect 436374 351922 436442 351978
rect 436498 351922 436568 351978
rect 436248 351888 436568 351922
rect 466968 352350 467288 352384
rect 466968 352294 467038 352350
rect 467094 352294 467162 352350
rect 467218 352294 467288 352350
rect 466968 352226 467288 352294
rect 466968 352170 467038 352226
rect 467094 352170 467162 352226
rect 467218 352170 467288 352226
rect 466968 352102 467288 352170
rect 466968 352046 467038 352102
rect 467094 352046 467162 352102
rect 467218 352046 467288 352102
rect 466968 351978 467288 352046
rect 466968 351922 467038 351978
rect 467094 351922 467162 351978
rect 467218 351922 467288 351978
rect 466968 351888 467288 351922
rect 497688 352350 498008 352384
rect 497688 352294 497758 352350
rect 497814 352294 497882 352350
rect 497938 352294 498008 352350
rect 497688 352226 498008 352294
rect 497688 352170 497758 352226
rect 497814 352170 497882 352226
rect 497938 352170 498008 352226
rect 497688 352102 498008 352170
rect 497688 352046 497758 352102
rect 497814 352046 497882 352102
rect 497938 352046 498008 352102
rect 497688 351978 498008 352046
rect 497688 351922 497758 351978
rect 497814 351922 497882 351978
rect 497938 351922 498008 351978
rect 497688 351888 498008 351922
rect 528408 352350 528728 352384
rect 528408 352294 528478 352350
rect 528534 352294 528602 352350
rect 528658 352294 528728 352350
rect 528408 352226 528728 352294
rect 528408 352170 528478 352226
rect 528534 352170 528602 352226
rect 528658 352170 528728 352226
rect 528408 352102 528728 352170
rect 528408 352046 528478 352102
rect 528534 352046 528602 352102
rect 528658 352046 528728 352102
rect 528408 351978 528728 352046
rect 528408 351922 528478 351978
rect 528534 351922 528602 351978
rect 528658 351922 528728 351978
rect 528408 351888 528728 351922
rect 559128 352350 559448 352384
rect 559128 352294 559198 352350
rect 559254 352294 559322 352350
rect 559378 352294 559448 352350
rect 559128 352226 559448 352294
rect 559128 352170 559198 352226
rect 559254 352170 559322 352226
rect 559378 352170 559448 352226
rect 559128 352102 559448 352170
rect 559128 352046 559198 352102
rect 559254 352046 559322 352102
rect 559378 352046 559448 352102
rect 559128 351978 559448 352046
rect 559128 351922 559198 351978
rect 559254 351922 559322 351978
rect 559378 351922 559448 351978
rect 559128 351888 559448 351922
rect 359448 346350 359768 346384
rect 359448 346294 359518 346350
rect 359574 346294 359642 346350
rect 359698 346294 359768 346350
rect 359448 346226 359768 346294
rect 359448 346170 359518 346226
rect 359574 346170 359642 346226
rect 359698 346170 359768 346226
rect 359448 346102 359768 346170
rect 359448 346046 359518 346102
rect 359574 346046 359642 346102
rect 359698 346046 359768 346102
rect 359448 345978 359768 346046
rect 359448 345922 359518 345978
rect 359574 345922 359642 345978
rect 359698 345922 359768 345978
rect 359448 345888 359768 345922
rect 390168 346350 390488 346384
rect 390168 346294 390238 346350
rect 390294 346294 390362 346350
rect 390418 346294 390488 346350
rect 390168 346226 390488 346294
rect 390168 346170 390238 346226
rect 390294 346170 390362 346226
rect 390418 346170 390488 346226
rect 390168 346102 390488 346170
rect 390168 346046 390238 346102
rect 390294 346046 390362 346102
rect 390418 346046 390488 346102
rect 390168 345978 390488 346046
rect 390168 345922 390238 345978
rect 390294 345922 390362 345978
rect 390418 345922 390488 345978
rect 390168 345888 390488 345922
rect 420888 346350 421208 346384
rect 420888 346294 420958 346350
rect 421014 346294 421082 346350
rect 421138 346294 421208 346350
rect 420888 346226 421208 346294
rect 420888 346170 420958 346226
rect 421014 346170 421082 346226
rect 421138 346170 421208 346226
rect 420888 346102 421208 346170
rect 420888 346046 420958 346102
rect 421014 346046 421082 346102
rect 421138 346046 421208 346102
rect 420888 345978 421208 346046
rect 420888 345922 420958 345978
rect 421014 345922 421082 345978
rect 421138 345922 421208 345978
rect 420888 345888 421208 345922
rect 451608 346350 451928 346384
rect 451608 346294 451678 346350
rect 451734 346294 451802 346350
rect 451858 346294 451928 346350
rect 451608 346226 451928 346294
rect 451608 346170 451678 346226
rect 451734 346170 451802 346226
rect 451858 346170 451928 346226
rect 451608 346102 451928 346170
rect 451608 346046 451678 346102
rect 451734 346046 451802 346102
rect 451858 346046 451928 346102
rect 451608 345978 451928 346046
rect 451608 345922 451678 345978
rect 451734 345922 451802 345978
rect 451858 345922 451928 345978
rect 451608 345888 451928 345922
rect 482328 346350 482648 346384
rect 482328 346294 482398 346350
rect 482454 346294 482522 346350
rect 482578 346294 482648 346350
rect 482328 346226 482648 346294
rect 482328 346170 482398 346226
rect 482454 346170 482522 346226
rect 482578 346170 482648 346226
rect 482328 346102 482648 346170
rect 482328 346046 482398 346102
rect 482454 346046 482522 346102
rect 482578 346046 482648 346102
rect 482328 345978 482648 346046
rect 482328 345922 482398 345978
rect 482454 345922 482522 345978
rect 482578 345922 482648 345978
rect 482328 345888 482648 345922
rect 513048 346350 513368 346384
rect 513048 346294 513118 346350
rect 513174 346294 513242 346350
rect 513298 346294 513368 346350
rect 513048 346226 513368 346294
rect 513048 346170 513118 346226
rect 513174 346170 513242 346226
rect 513298 346170 513368 346226
rect 513048 346102 513368 346170
rect 513048 346046 513118 346102
rect 513174 346046 513242 346102
rect 513298 346046 513368 346102
rect 513048 345978 513368 346046
rect 513048 345922 513118 345978
rect 513174 345922 513242 345978
rect 513298 345922 513368 345978
rect 513048 345888 513368 345922
rect 543768 346350 544088 346384
rect 543768 346294 543838 346350
rect 543894 346294 543962 346350
rect 544018 346294 544088 346350
rect 543768 346226 544088 346294
rect 543768 346170 543838 346226
rect 543894 346170 543962 346226
rect 544018 346170 544088 346226
rect 543768 346102 544088 346170
rect 543768 346046 543838 346102
rect 543894 346046 543962 346102
rect 544018 346046 544088 346102
rect 543768 345978 544088 346046
rect 543768 345922 543838 345978
rect 543894 345922 543962 345978
rect 544018 345922 544088 345978
rect 543768 345888 544088 345922
rect 574488 346350 574808 346384
rect 574488 346294 574558 346350
rect 574614 346294 574682 346350
rect 574738 346294 574808 346350
rect 574488 346226 574808 346294
rect 574488 346170 574558 346226
rect 574614 346170 574682 346226
rect 574738 346170 574808 346226
rect 574488 346102 574808 346170
rect 574488 346046 574558 346102
rect 574614 346046 574682 346102
rect 574738 346046 574808 346102
rect 574488 345978 574808 346046
rect 574488 345922 574558 345978
rect 574614 345922 574682 345978
rect 574738 345922 574808 345978
rect 574488 345888 574808 345922
rect 374808 334350 375128 334384
rect 374808 334294 374878 334350
rect 374934 334294 375002 334350
rect 375058 334294 375128 334350
rect 374808 334226 375128 334294
rect 374808 334170 374878 334226
rect 374934 334170 375002 334226
rect 375058 334170 375128 334226
rect 374808 334102 375128 334170
rect 374808 334046 374878 334102
rect 374934 334046 375002 334102
rect 375058 334046 375128 334102
rect 374808 333978 375128 334046
rect 374808 333922 374878 333978
rect 374934 333922 375002 333978
rect 375058 333922 375128 333978
rect 374808 333888 375128 333922
rect 405528 334350 405848 334384
rect 405528 334294 405598 334350
rect 405654 334294 405722 334350
rect 405778 334294 405848 334350
rect 405528 334226 405848 334294
rect 405528 334170 405598 334226
rect 405654 334170 405722 334226
rect 405778 334170 405848 334226
rect 405528 334102 405848 334170
rect 405528 334046 405598 334102
rect 405654 334046 405722 334102
rect 405778 334046 405848 334102
rect 405528 333978 405848 334046
rect 405528 333922 405598 333978
rect 405654 333922 405722 333978
rect 405778 333922 405848 333978
rect 405528 333888 405848 333922
rect 436248 334350 436568 334384
rect 436248 334294 436318 334350
rect 436374 334294 436442 334350
rect 436498 334294 436568 334350
rect 436248 334226 436568 334294
rect 436248 334170 436318 334226
rect 436374 334170 436442 334226
rect 436498 334170 436568 334226
rect 436248 334102 436568 334170
rect 436248 334046 436318 334102
rect 436374 334046 436442 334102
rect 436498 334046 436568 334102
rect 436248 333978 436568 334046
rect 436248 333922 436318 333978
rect 436374 333922 436442 333978
rect 436498 333922 436568 333978
rect 436248 333888 436568 333922
rect 466968 334350 467288 334384
rect 466968 334294 467038 334350
rect 467094 334294 467162 334350
rect 467218 334294 467288 334350
rect 466968 334226 467288 334294
rect 466968 334170 467038 334226
rect 467094 334170 467162 334226
rect 467218 334170 467288 334226
rect 466968 334102 467288 334170
rect 466968 334046 467038 334102
rect 467094 334046 467162 334102
rect 467218 334046 467288 334102
rect 466968 333978 467288 334046
rect 466968 333922 467038 333978
rect 467094 333922 467162 333978
rect 467218 333922 467288 333978
rect 466968 333888 467288 333922
rect 497688 334350 498008 334384
rect 497688 334294 497758 334350
rect 497814 334294 497882 334350
rect 497938 334294 498008 334350
rect 497688 334226 498008 334294
rect 497688 334170 497758 334226
rect 497814 334170 497882 334226
rect 497938 334170 498008 334226
rect 497688 334102 498008 334170
rect 497688 334046 497758 334102
rect 497814 334046 497882 334102
rect 497938 334046 498008 334102
rect 497688 333978 498008 334046
rect 497688 333922 497758 333978
rect 497814 333922 497882 333978
rect 497938 333922 498008 333978
rect 497688 333888 498008 333922
rect 528408 334350 528728 334384
rect 528408 334294 528478 334350
rect 528534 334294 528602 334350
rect 528658 334294 528728 334350
rect 528408 334226 528728 334294
rect 528408 334170 528478 334226
rect 528534 334170 528602 334226
rect 528658 334170 528728 334226
rect 528408 334102 528728 334170
rect 528408 334046 528478 334102
rect 528534 334046 528602 334102
rect 528658 334046 528728 334102
rect 528408 333978 528728 334046
rect 528408 333922 528478 333978
rect 528534 333922 528602 333978
rect 528658 333922 528728 333978
rect 528408 333888 528728 333922
rect 559128 334350 559448 334384
rect 559128 334294 559198 334350
rect 559254 334294 559322 334350
rect 559378 334294 559448 334350
rect 559128 334226 559448 334294
rect 559128 334170 559198 334226
rect 559254 334170 559322 334226
rect 559378 334170 559448 334226
rect 559128 334102 559448 334170
rect 559128 334046 559198 334102
rect 559254 334046 559322 334102
rect 559378 334046 559448 334102
rect 559128 333978 559448 334046
rect 559128 333922 559198 333978
rect 559254 333922 559322 333978
rect 559378 333922 559448 333978
rect 559128 333888 559448 333922
rect 359448 328350 359768 328384
rect 359448 328294 359518 328350
rect 359574 328294 359642 328350
rect 359698 328294 359768 328350
rect 359448 328226 359768 328294
rect 359448 328170 359518 328226
rect 359574 328170 359642 328226
rect 359698 328170 359768 328226
rect 359448 328102 359768 328170
rect 359448 328046 359518 328102
rect 359574 328046 359642 328102
rect 359698 328046 359768 328102
rect 359448 327978 359768 328046
rect 359448 327922 359518 327978
rect 359574 327922 359642 327978
rect 359698 327922 359768 327978
rect 359448 327888 359768 327922
rect 390168 328350 390488 328384
rect 390168 328294 390238 328350
rect 390294 328294 390362 328350
rect 390418 328294 390488 328350
rect 390168 328226 390488 328294
rect 390168 328170 390238 328226
rect 390294 328170 390362 328226
rect 390418 328170 390488 328226
rect 390168 328102 390488 328170
rect 390168 328046 390238 328102
rect 390294 328046 390362 328102
rect 390418 328046 390488 328102
rect 390168 327978 390488 328046
rect 390168 327922 390238 327978
rect 390294 327922 390362 327978
rect 390418 327922 390488 327978
rect 390168 327888 390488 327922
rect 420888 328350 421208 328384
rect 420888 328294 420958 328350
rect 421014 328294 421082 328350
rect 421138 328294 421208 328350
rect 420888 328226 421208 328294
rect 420888 328170 420958 328226
rect 421014 328170 421082 328226
rect 421138 328170 421208 328226
rect 420888 328102 421208 328170
rect 420888 328046 420958 328102
rect 421014 328046 421082 328102
rect 421138 328046 421208 328102
rect 420888 327978 421208 328046
rect 420888 327922 420958 327978
rect 421014 327922 421082 327978
rect 421138 327922 421208 327978
rect 420888 327888 421208 327922
rect 451608 328350 451928 328384
rect 451608 328294 451678 328350
rect 451734 328294 451802 328350
rect 451858 328294 451928 328350
rect 451608 328226 451928 328294
rect 451608 328170 451678 328226
rect 451734 328170 451802 328226
rect 451858 328170 451928 328226
rect 451608 328102 451928 328170
rect 451608 328046 451678 328102
rect 451734 328046 451802 328102
rect 451858 328046 451928 328102
rect 451608 327978 451928 328046
rect 451608 327922 451678 327978
rect 451734 327922 451802 327978
rect 451858 327922 451928 327978
rect 451608 327888 451928 327922
rect 482328 328350 482648 328384
rect 482328 328294 482398 328350
rect 482454 328294 482522 328350
rect 482578 328294 482648 328350
rect 482328 328226 482648 328294
rect 482328 328170 482398 328226
rect 482454 328170 482522 328226
rect 482578 328170 482648 328226
rect 482328 328102 482648 328170
rect 482328 328046 482398 328102
rect 482454 328046 482522 328102
rect 482578 328046 482648 328102
rect 482328 327978 482648 328046
rect 482328 327922 482398 327978
rect 482454 327922 482522 327978
rect 482578 327922 482648 327978
rect 482328 327888 482648 327922
rect 513048 328350 513368 328384
rect 513048 328294 513118 328350
rect 513174 328294 513242 328350
rect 513298 328294 513368 328350
rect 513048 328226 513368 328294
rect 513048 328170 513118 328226
rect 513174 328170 513242 328226
rect 513298 328170 513368 328226
rect 513048 328102 513368 328170
rect 513048 328046 513118 328102
rect 513174 328046 513242 328102
rect 513298 328046 513368 328102
rect 513048 327978 513368 328046
rect 513048 327922 513118 327978
rect 513174 327922 513242 327978
rect 513298 327922 513368 327978
rect 513048 327888 513368 327922
rect 543768 328350 544088 328384
rect 543768 328294 543838 328350
rect 543894 328294 543962 328350
rect 544018 328294 544088 328350
rect 543768 328226 544088 328294
rect 543768 328170 543838 328226
rect 543894 328170 543962 328226
rect 544018 328170 544088 328226
rect 543768 328102 544088 328170
rect 543768 328046 543838 328102
rect 543894 328046 543962 328102
rect 544018 328046 544088 328102
rect 543768 327978 544088 328046
rect 543768 327922 543838 327978
rect 543894 327922 543962 327978
rect 544018 327922 544088 327978
rect 543768 327888 544088 327922
rect 574488 328350 574808 328384
rect 574488 328294 574558 328350
rect 574614 328294 574682 328350
rect 574738 328294 574808 328350
rect 574488 328226 574808 328294
rect 574488 328170 574558 328226
rect 574614 328170 574682 328226
rect 574738 328170 574808 328226
rect 574488 328102 574808 328170
rect 574488 328046 574558 328102
rect 574614 328046 574682 328102
rect 574738 328046 574808 328102
rect 574488 327978 574808 328046
rect 574488 327922 574558 327978
rect 574614 327922 574682 327978
rect 574738 327922 574808 327978
rect 574488 327888 574808 327922
rect 374808 316350 375128 316384
rect 374808 316294 374878 316350
rect 374934 316294 375002 316350
rect 375058 316294 375128 316350
rect 374808 316226 375128 316294
rect 374808 316170 374878 316226
rect 374934 316170 375002 316226
rect 375058 316170 375128 316226
rect 374808 316102 375128 316170
rect 374808 316046 374878 316102
rect 374934 316046 375002 316102
rect 375058 316046 375128 316102
rect 374808 315978 375128 316046
rect 374808 315922 374878 315978
rect 374934 315922 375002 315978
rect 375058 315922 375128 315978
rect 374808 315888 375128 315922
rect 405528 316350 405848 316384
rect 405528 316294 405598 316350
rect 405654 316294 405722 316350
rect 405778 316294 405848 316350
rect 405528 316226 405848 316294
rect 405528 316170 405598 316226
rect 405654 316170 405722 316226
rect 405778 316170 405848 316226
rect 405528 316102 405848 316170
rect 405528 316046 405598 316102
rect 405654 316046 405722 316102
rect 405778 316046 405848 316102
rect 405528 315978 405848 316046
rect 405528 315922 405598 315978
rect 405654 315922 405722 315978
rect 405778 315922 405848 315978
rect 405528 315888 405848 315922
rect 436248 316350 436568 316384
rect 436248 316294 436318 316350
rect 436374 316294 436442 316350
rect 436498 316294 436568 316350
rect 436248 316226 436568 316294
rect 436248 316170 436318 316226
rect 436374 316170 436442 316226
rect 436498 316170 436568 316226
rect 436248 316102 436568 316170
rect 436248 316046 436318 316102
rect 436374 316046 436442 316102
rect 436498 316046 436568 316102
rect 436248 315978 436568 316046
rect 436248 315922 436318 315978
rect 436374 315922 436442 315978
rect 436498 315922 436568 315978
rect 436248 315888 436568 315922
rect 466968 316350 467288 316384
rect 466968 316294 467038 316350
rect 467094 316294 467162 316350
rect 467218 316294 467288 316350
rect 466968 316226 467288 316294
rect 466968 316170 467038 316226
rect 467094 316170 467162 316226
rect 467218 316170 467288 316226
rect 466968 316102 467288 316170
rect 466968 316046 467038 316102
rect 467094 316046 467162 316102
rect 467218 316046 467288 316102
rect 466968 315978 467288 316046
rect 466968 315922 467038 315978
rect 467094 315922 467162 315978
rect 467218 315922 467288 315978
rect 466968 315888 467288 315922
rect 497688 316350 498008 316384
rect 497688 316294 497758 316350
rect 497814 316294 497882 316350
rect 497938 316294 498008 316350
rect 497688 316226 498008 316294
rect 497688 316170 497758 316226
rect 497814 316170 497882 316226
rect 497938 316170 498008 316226
rect 497688 316102 498008 316170
rect 497688 316046 497758 316102
rect 497814 316046 497882 316102
rect 497938 316046 498008 316102
rect 497688 315978 498008 316046
rect 497688 315922 497758 315978
rect 497814 315922 497882 315978
rect 497938 315922 498008 315978
rect 497688 315888 498008 315922
rect 528408 316350 528728 316384
rect 528408 316294 528478 316350
rect 528534 316294 528602 316350
rect 528658 316294 528728 316350
rect 528408 316226 528728 316294
rect 528408 316170 528478 316226
rect 528534 316170 528602 316226
rect 528658 316170 528728 316226
rect 528408 316102 528728 316170
rect 528408 316046 528478 316102
rect 528534 316046 528602 316102
rect 528658 316046 528728 316102
rect 528408 315978 528728 316046
rect 528408 315922 528478 315978
rect 528534 315922 528602 315978
rect 528658 315922 528728 315978
rect 528408 315888 528728 315922
rect 559128 316350 559448 316384
rect 559128 316294 559198 316350
rect 559254 316294 559322 316350
rect 559378 316294 559448 316350
rect 559128 316226 559448 316294
rect 559128 316170 559198 316226
rect 559254 316170 559322 316226
rect 559378 316170 559448 316226
rect 559128 316102 559448 316170
rect 559128 316046 559198 316102
rect 559254 316046 559322 316102
rect 559378 316046 559448 316102
rect 559128 315978 559448 316046
rect 559128 315922 559198 315978
rect 559254 315922 559322 315978
rect 559378 315922 559448 315978
rect 559128 315888 559448 315922
rect 359448 310350 359768 310384
rect 359448 310294 359518 310350
rect 359574 310294 359642 310350
rect 359698 310294 359768 310350
rect 359448 310226 359768 310294
rect 359448 310170 359518 310226
rect 359574 310170 359642 310226
rect 359698 310170 359768 310226
rect 359448 310102 359768 310170
rect 359448 310046 359518 310102
rect 359574 310046 359642 310102
rect 359698 310046 359768 310102
rect 359448 309978 359768 310046
rect 359448 309922 359518 309978
rect 359574 309922 359642 309978
rect 359698 309922 359768 309978
rect 359448 309888 359768 309922
rect 390168 310350 390488 310384
rect 390168 310294 390238 310350
rect 390294 310294 390362 310350
rect 390418 310294 390488 310350
rect 390168 310226 390488 310294
rect 390168 310170 390238 310226
rect 390294 310170 390362 310226
rect 390418 310170 390488 310226
rect 390168 310102 390488 310170
rect 390168 310046 390238 310102
rect 390294 310046 390362 310102
rect 390418 310046 390488 310102
rect 390168 309978 390488 310046
rect 390168 309922 390238 309978
rect 390294 309922 390362 309978
rect 390418 309922 390488 309978
rect 390168 309888 390488 309922
rect 420888 310350 421208 310384
rect 420888 310294 420958 310350
rect 421014 310294 421082 310350
rect 421138 310294 421208 310350
rect 420888 310226 421208 310294
rect 420888 310170 420958 310226
rect 421014 310170 421082 310226
rect 421138 310170 421208 310226
rect 420888 310102 421208 310170
rect 420888 310046 420958 310102
rect 421014 310046 421082 310102
rect 421138 310046 421208 310102
rect 420888 309978 421208 310046
rect 420888 309922 420958 309978
rect 421014 309922 421082 309978
rect 421138 309922 421208 309978
rect 420888 309888 421208 309922
rect 451608 310350 451928 310384
rect 451608 310294 451678 310350
rect 451734 310294 451802 310350
rect 451858 310294 451928 310350
rect 451608 310226 451928 310294
rect 451608 310170 451678 310226
rect 451734 310170 451802 310226
rect 451858 310170 451928 310226
rect 451608 310102 451928 310170
rect 451608 310046 451678 310102
rect 451734 310046 451802 310102
rect 451858 310046 451928 310102
rect 451608 309978 451928 310046
rect 451608 309922 451678 309978
rect 451734 309922 451802 309978
rect 451858 309922 451928 309978
rect 451608 309888 451928 309922
rect 482328 310350 482648 310384
rect 482328 310294 482398 310350
rect 482454 310294 482522 310350
rect 482578 310294 482648 310350
rect 482328 310226 482648 310294
rect 482328 310170 482398 310226
rect 482454 310170 482522 310226
rect 482578 310170 482648 310226
rect 482328 310102 482648 310170
rect 482328 310046 482398 310102
rect 482454 310046 482522 310102
rect 482578 310046 482648 310102
rect 482328 309978 482648 310046
rect 482328 309922 482398 309978
rect 482454 309922 482522 309978
rect 482578 309922 482648 309978
rect 482328 309888 482648 309922
rect 513048 310350 513368 310384
rect 513048 310294 513118 310350
rect 513174 310294 513242 310350
rect 513298 310294 513368 310350
rect 513048 310226 513368 310294
rect 513048 310170 513118 310226
rect 513174 310170 513242 310226
rect 513298 310170 513368 310226
rect 513048 310102 513368 310170
rect 513048 310046 513118 310102
rect 513174 310046 513242 310102
rect 513298 310046 513368 310102
rect 513048 309978 513368 310046
rect 513048 309922 513118 309978
rect 513174 309922 513242 309978
rect 513298 309922 513368 309978
rect 513048 309888 513368 309922
rect 543768 310350 544088 310384
rect 543768 310294 543838 310350
rect 543894 310294 543962 310350
rect 544018 310294 544088 310350
rect 543768 310226 544088 310294
rect 543768 310170 543838 310226
rect 543894 310170 543962 310226
rect 544018 310170 544088 310226
rect 543768 310102 544088 310170
rect 543768 310046 543838 310102
rect 543894 310046 543962 310102
rect 544018 310046 544088 310102
rect 543768 309978 544088 310046
rect 543768 309922 543838 309978
rect 543894 309922 543962 309978
rect 544018 309922 544088 309978
rect 543768 309888 544088 309922
rect 574488 310350 574808 310384
rect 574488 310294 574558 310350
rect 574614 310294 574682 310350
rect 574738 310294 574808 310350
rect 574488 310226 574808 310294
rect 574488 310170 574558 310226
rect 574614 310170 574682 310226
rect 574738 310170 574808 310226
rect 574488 310102 574808 310170
rect 574488 310046 574558 310102
rect 574614 310046 574682 310102
rect 574738 310046 574808 310102
rect 574488 309978 574808 310046
rect 574488 309922 574558 309978
rect 574614 309922 574682 309978
rect 574738 309922 574808 309978
rect 574488 309888 574808 309922
rect 374808 298350 375128 298384
rect 374808 298294 374878 298350
rect 374934 298294 375002 298350
rect 375058 298294 375128 298350
rect 374808 298226 375128 298294
rect 374808 298170 374878 298226
rect 374934 298170 375002 298226
rect 375058 298170 375128 298226
rect 374808 298102 375128 298170
rect 374808 298046 374878 298102
rect 374934 298046 375002 298102
rect 375058 298046 375128 298102
rect 374808 297978 375128 298046
rect 374808 297922 374878 297978
rect 374934 297922 375002 297978
rect 375058 297922 375128 297978
rect 374808 297888 375128 297922
rect 405528 298350 405848 298384
rect 405528 298294 405598 298350
rect 405654 298294 405722 298350
rect 405778 298294 405848 298350
rect 405528 298226 405848 298294
rect 405528 298170 405598 298226
rect 405654 298170 405722 298226
rect 405778 298170 405848 298226
rect 405528 298102 405848 298170
rect 405528 298046 405598 298102
rect 405654 298046 405722 298102
rect 405778 298046 405848 298102
rect 405528 297978 405848 298046
rect 405528 297922 405598 297978
rect 405654 297922 405722 297978
rect 405778 297922 405848 297978
rect 405528 297888 405848 297922
rect 436248 298350 436568 298384
rect 436248 298294 436318 298350
rect 436374 298294 436442 298350
rect 436498 298294 436568 298350
rect 436248 298226 436568 298294
rect 436248 298170 436318 298226
rect 436374 298170 436442 298226
rect 436498 298170 436568 298226
rect 436248 298102 436568 298170
rect 436248 298046 436318 298102
rect 436374 298046 436442 298102
rect 436498 298046 436568 298102
rect 436248 297978 436568 298046
rect 436248 297922 436318 297978
rect 436374 297922 436442 297978
rect 436498 297922 436568 297978
rect 436248 297888 436568 297922
rect 466968 298350 467288 298384
rect 466968 298294 467038 298350
rect 467094 298294 467162 298350
rect 467218 298294 467288 298350
rect 466968 298226 467288 298294
rect 466968 298170 467038 298226
rect 467094 298170 467162 298226
rect 467218 298170 467288 298226
rect 466968 298102 467288 298170
rect 466968 298046 467038 298102
rect 467094 298046 467162 298102
rect 467218 298046 467288 298102
rect 466968 297978 467288 298046
rect 466968 297922 467038 297978
rect 467094 297922 467162 297978
rect 467218 297922 467288 297978
rect 466968 297888 467288 297922
rect 497688 298350 498008 298384
rect 497688 298294 497758 298350
rect 497814 298294 497882 298350
rect 497938 298294 498008 298350
rect 497688 298226 498008 298294
rect 497688 298170 497758 298226
rect 497814 298170 497882 298226
rect 497938 298170 498008 298226
rect 497688 298102 498008 298170
rect 497688 298046 497758 298102
rect 497814 298046 497882 298102
rect 497938 298046 498008 298102
rect 497688 297978 498008 298046
rect 497688 297922 497758 297978
rect 497814 297922 497882 297978
rect 497938 297922 498008 297978
rect 497688 297888 498008 297922
rect 528408 298350 528728 298384
rect 528408 298294 528478 298350
rect 528534 298294 528602 298350
rect 528658 298294 528728 298350
rect 528408 298226 528728 298294
rect 528408 298170 528478 298226
rect 528534 298170 528602 298226
rect 528658 298170 528728 298226
rect 528408 298102 528728 298170
rect 528408 298046 528478 298102
rect 528534 298046 528602 298102
rect 528658 298046 528728 298102
rect 528408 297978 528728 298046
rect 528408 297922 528478 297978
rect 528534 297922 528602 297978
rect 528658 297922 528728 297978
rect 528408 297888 528728 297922
rect 559128 298350 559448 298384
rect 559128 298294 559198 298350
rect 559254 298294 559322 298350
rect 559378 298294 559448 298350
rect 559128 298226 559448 298294
rect 559128 298170 559198 298226
rect 559254 298170 559322 298226
rect 559378 298170 559448 298226
rect 559128 298102 559448 298170
rect 559128 298046 559198 298102
rect 559254 298046 559322 298102
rect 559378 298046 559448 298102
rect 559128 297978 559448 298046
rect 559128 297922 559198 297978
rect 559254 297922 559322 297978
rect 559378 297922 559448 297978
rect 559128 297888 559448 297922
rect 359448 292350 359768 292384
rect 359448 292294 359518 292350
rect 359574 292294 359642 292350
rect 359698 292294 359768 292350
rect 359448 292226 359768 292294
rect 359448 292170 359518 292226
rect 359574 292170 359642 292226
rect 359698 292170 359768 292226
rect 359448 292102 359768 292170
rect 359448 292046 359518 292102
rect 359574 292046 359642 292102
rect 359698 292046 359768 292102
rect 359448 291978 359768 292046
rect 359448 291922 359518 291978
rect 359574 291922 359642 291978
rect 359698 291922 359768 291978
rect 359448 291888 359768 291922
rect 390168 292350 390488 292384
rect 390168 292294 390238 292350
rect 390294 292294 390362 292350
rect 390418 292294 390488 292350
rect 390168 292226 390488 292294
rect 390168 292170 390238 292226
rect 390294 292170 390362 292226
rect 390418 292170 390488 292226
rect 390168 292102 390488 292170
rect 390168 292046 390238 292102
rect 390294 292046 390362 292102
rect 390418 292046 390488 292102
rect 390168 291978 390488 292046
rect 390168 291922 390238 291978
rect 390294 291922 390362 291978
rect 390418 291922 390488 291978
rect 390168 291888 390488 291922
rect 420888 292350 421208 292384
rect 420888 292294 420958 292350
rect 421014 292294 421082 292350
rect 421138 292294 421208 292350
rect 420888 292226 421208 292294
rect 420888 292170 420958 292226
rect 421014 292170 421082 292226
rect 421138 292170 421208 292226
rect 420888 292102 421208 292170
rect 420888 292046 420958 292102
rect 421014 292046 421082 292102
rect 421138 292046 421208 292102
rect 420888 291978 421208 292046
rect 420888 291922 420958 291978
rect 421014 291922 421082 291978
rect 421138 291922 421208 291978
rect 420888 291888 421208 291922
rect 451608 292350 451928 292384
rect 451608 292294 451678 292350
rect 451734 292294 451802 292350
rect 451858 292294 451928 292350
rect 451608 292226 451928 292294
rect 451608 292170 451678 292226
rect 451734 292170 451802 292226
rect 451858 292170 451928 292226
rect 451608 292102 451928 292170
rect 451608 292046 451678 292102
rect 451734 292046 451802 292102
rect 451858 292046 451928 292102
rect 451608 291978 451928 292046
rect 451608 291922 451678 291978
rect 451734 291922 451802 291978
rect 451858 291922 451928 291978
rect 451608 291888 451928 291922
rect 482328 292350 482648 292384
rect 482328 292294 482398 292350
rect 482454 292294 482522 292350
rect 482578 292294 482648 292350
rect 482328 292226 482648 292294
rect 482328 292170 482398 292226
rect 482454 292170 482522 292226
rect 482578 292170 482648 292226
rect 482328 292102 482648 292170
rect 482328 292046 482398 292102
rect 482454 292046 482522 292102
rect 482578 292046 482648 292102
rect 482328 291978 482648 292046
rect 482328 291922 482398 291978
rect 482454 291922 482522 291978
rect 482578 291922 482648 291978
rect 482328 291888 482648 291922
rect 513048 292350 513368 292384
rect 513048 292294 513118 292350
rect 513174 292294 513242 292350
rect 513298 292294 513368 292350
rect 513048 292226 513368 292294
rect 513048 292170 513118 292226
rect 513174 292170 513242 292226
rect 513298 292170 513368 292226
rect 513048 292102 513368 292170
rect 513048 292046 513118 292102
rect 513174 292046 513242 292102
rect 513298 292046 513368 292102
rect 513048 291978 513368 292046
rect 513048 291922 513118 291978
rect 513174 291922 513242 291978
rect 513298 291922 513368 291978
rect 513048 291888 513368 291922
rect 543768 292350 544088 292384
rect 543768 292294 543838 292350
rect 543894 292294 543962 292350
rect 544018 292294 544088 292350
rect 543768 292226 544088 292294
rect 543768 292170 543838 292226
rect 543894 292170 543962 292226
rect 544018 292170 544088 292226
rect 543768 292102 544088 292170
rect 543768 292046 543838 292102
rect 543894 292046 543962 292102
rect 544018 292046 544088 292102
rect 543768 291978 544088 292046
rect 543768 291922 543838 291978
rect 543894 291922 543962 291978
rect 544018 291922 544088 291978
rect 543768 291888 544088 291922
rect 574488 292350 574808 292384
rect 574488 292294 574558 292350
rect 574614 292294 574682 292350
rect 574738 292294 574808 292350
rect 574488 292226 574808 292294
rect 574488 292170 574558 292226
rect 574614 292170 574682 292226
rect 574738 292170 574808 292226
rect 574488 292102 574808 292170
rect 574488 292046 574558 292102
rect 574614 292046 574682 292102
rect 574738 292046 574808 292102
rect 574488 291978 574808 292046
rect 574488 291922 574558 291978
rect 574614 291922 574682 291978
rect 574738 291922 574808 291978
rect 574488 291888 574808 291922
rect 374808 280350 375128 280384
rect 374808 280294 374878 280350
rect 374934 280294 375002 280350
rect 375058 280294 375128 280350
rect 374808 280226 375128 280294
rect 374808 280170 374878 280226
rect 374934 280170 375002 280226
rect 375058 280170 375128 280226
rect 374808 280102 375128 280170
rect 374808 280046 374878 280102
rect 374934 280046 375002 280102
rect 375058 280046 375128 280102
rect 374808 279978 375128 280046
rect 374808 279922 374878 279978
rect 374934 279922 375002 279978
rect 375058 279922 375128 279978
rect 374808 279888 375128 279922
rect 405528 280350 405848 280384
rect 405528 280294 405598 280350
rect 405654 280294 405722 280350
rect 405778 280294 405848 280350
rect 405528 280226 405848 280294
rect 405528 280170 405598 280226
rect 405654 280170 405722 280226
rect 405778 280170 405848 280226
rect 405528 280102 405848 280170
rect 405528 280046 405598 280102
rect 405654 280046 405722 280102
rect 405778 280046 405848 280102
rect 405528 279978 405848 280046
rect 405528 279922 405598 279978
rect 405654 279922 405722 279978
rect 405778 279922 405848 279978
rect 405528 279888 405848 279922
rect 436248 280350 436568 280384
rect 436248 280294 436318 280350
rect 436374 280294 436442 280350
rect 436498 280294 436568 280350
rect 436248 280226 436568 280294
rect 436248 280170 436318 280226
rect 436374 280170 436442 280226
rect 436498 280170 436568 280226
rect 436248 280102 436568 280170
rect 436248 280046 436318 280102
rect 436374 280046 436442 280102
rect 436498 280046 436568 280102
rect 436248 279978 436568 280046
rect 436248 279922 436318 279978
rect 436374 279922 436442 279978
rect 436498 279922 436568 279978
rect 436248 279888 436568 279922
rect 466968 280350 467288 280384
rect 466968 280294 467038 280350
rect 467094 280294 467162 280350
rect 467218 280294 467288 280350
rect 466968 280226 467288 280294
rect 466968 280170 467038 280226
rect 467094 280170 467162 280226
rect 467218 280170 467288 280226
rect 466968 280102 467288 280170
rect 466968 280046 467038 280102
rect 467094 280046 467162 280102
rect 467218 280046 467288 280102
rect 466968 279978 467288 280046
rect 466968 279922 467038 279978
rect 467094 279922 467162 279978
rect 467218 279922 467288 279978
rect 466968 279888 467288 279922
rect 497688 280350 498008 280384
rect 497688 280294 497758 280350
rect 497814 280294 497882 280350
rect 497938 280294 498008 280350
rect 497688 280226 498008 280294
rect 497688 280170 497758 280226
rect 497814 280170 497882 280226
rect 497938 280170 498008 280226
rect 497688 280102 498008 280170
rect 497688 280046 497758 280102
rect 497814 280046 497882 280102
rect 497938 280046 498008 280102
rect 497688 279978 498008 280046
rect 497688 279922 497758 279978
rect 497814 279922 497882 279978
rect 497938 279922 498008 279978
rect 497688 279888 498008 279922
rect 528408 280350 528728 280384
rect 528408 280294 528478 280350
rect 528534 280294 528602 280350
rect 528658 280294 528728 280350
rect 528408 280226 528728 280294
rect 528408 280170 528478 280226
rect 528534 280170 528602 280226
rect 528658 280170 528728 280226
rect 528408 280102 528728 280170
rect 528408 280046 528478 280102
rect 528534 280046 528602 280102
rect 528658 280046 528728 280102
rect 528408 279978 528728 280046
rect 528408 279922 528478 279978
rect 528534 279922 528602 279978
rect 528658 279922 528728 279978
rect 528408 279888 528728 279922
rect 559128 280350 559448 280384
rect 559128 280294 559198 280350
rect 559254 280294 559322 280350
rect 559378 280294 559448 280350
rect 559128 280226 559448 280294
rect 559128 280170 559198 280226
rect 559254 280170 559322 280226
rect 559378 280170 559448 280226
rect 559128 280102 559448 280170
rect 559128 280046 559198 280102
rect 559254 280046 559322 280102
rect 559378 280046 559448 280102
rect 559128 279978 559448 280046
rect 559128 279922 559198 279978
rect 559254 279922 559322 279978
rect 559378 279922 559448 279978
rect 559128 279888 559448 279922
rect 359448 274350 359768 274384
rect 359448 274294 359518 274350
rect 359574 274294 359642 274350
rect 359698 274294 359768 274350
rect 359448 274226 359768 274294
rect 359448 274170 359518 274226
rect 359574 274170 359642 274226
rect 359698 274170 359768 274226
rect 359448 274102 359768 274170
rect 359448 274046 359518 274102
rect 359574 274046 359642 274102
rect 359698 274046 359768 274102
rect 359448 273978 359768 274046
rect 359448 273922 359518 273978
rect 359574 273922 359642 273978
rect 359698 273922 359768 273978
rect 359448 273888 359768 273922
rect 390168 274350 390488 274384
rect 390168 274294 390238 274350
rect 390294 274294 390362 274350
rect 390418 274294 390488 274350
rect 390168 274226 390488 274294
rect 390168 274170 390238 274226
rect 390294 274170 390362 274226
rect 390418 274170 390488 274226
rect 390168 274102 390488 274170
rect 390168 274046 390238 274102
rect 390294 274046 390362 274102
rect 390418 274046 390488 274102
rect 390168 273978 390488 274046
rect 390168 273922 390238 273978
rect 390294 273922 390362 273978
rect 390418 273922 390488 273978
rect 390168 273888 390488 273922
rect 420888 274350 421208 274384
rect 420888 274294 420958 274350
rect 421014 274294 421082 274350
rect 421138 274294 421208 274350
rect 420888 274226 421208 274294
rect 420888 274170 420958 274226
rect 421014 274170 421082 274226
rect 421138 274170 421208 274226
rect 420888 274102 421208 274170
rect 420888 274046 420958 274102
rect 421014 274046 421082 274102
rect 421138 274046 421208 274102
rect 420888 273978 421208 274046
rect 420888 273922 420958 273978
rect 421014 273922 421082 273978
rect 421138 273922 421208 273978
rect 420888 273888 421208 273922
rect 451608 274350 451928 274384
rect 451608 274294 451678 274350
rect 451734 274294 451802 274350
rect 451858 274294 451928 274350
rect 451608 274226 451928 274294
rect 451608 274170 451678 274226
rect 451734 274170 451802 274226
rect 451858 274170 451928 274226
rect 451608 274102 451928 274170
rect 451608 274046 451678 274102
rect 451734 274046 451802 274102
rect 451858 274046 451928 274102
rect 451608 273978 451928 274046
rect 451608 273922 451678 273978
rect 451734 273922 451802 273978
rect 451858 273922 451928 273978
rect 451608 273888 451928 273922
rect 482328 274350 482648 274384
rect 482328 274294 482398 274350
rect 482454 274294 482522 274350
rect 482578 274294 482648 274350
rect 482328 274226 482648 274294
rect 482328 274170 482398 274226
rect 482454 274170 482522 274226
rect 482578 274170 482648 274226
rect 482328 274102 482648 274170
rect 482328 274046 482398 274102
rect 482454 274046 482522 274102
rect 482578 274046 482648 274102
rect 482328 273978 482648 274046
rect 482328 273922 482398 273978
rect 482454 273922 482522 273978
rect 482578 273922 482648 273978
rect 482328 273888 482648 273922
rect 513048 274350 513368 274384
rect 513048 274294 513118 274350
rect 513174 274294 513242 274350
rect 513298 274294 513368 274350
rect 513048 274226 513368 274294
rect 513048 274170 513118 274226
rect 513174 274170 513242 274226
rect 513298 274170 513368 274226
rect 513048 274102 513368 274170
rect 513048 274046 513118 274102
rect 513174 274046 513242 274102
rect 513298 274046 513368 274102
rect 513048 273978 513368 274046
rect 513048 273922 513118 273978
rect 513174 273922 513242 273978
rect 513298 273922 513368 273978
rect 513048 273888 513368 273922
rect 543768 274350 544088 274384
rect 543768 274294 543838 274350
rect 543894 274294 543962 274350
rect 544018 274294 544088 274350
rect 543768 274226 544088 274294
rect 543768 274170 543838 274226
rect 543894 274170 543962 274226
rect 544018 274170 544088 274226
rect 543768 274102 544088 274170
rect 543768 274046 543838 274102
rect 543894 274046 543962 274102
rect 544018 274046 544088 274102
rect 543768 273978 544088 274046
rect 543768 273922 543838 273978
rect 543894 273922 543962 273978
rect 544018 273922 544088 273978
rect 543768 273888 544088 273922
rect 574488 274350 574808 274384
rect 574488 274294 574558 274350
rect 574614 274294 574682 274350
rect 574738 274294 574808 274350
rect 574488 274226 574808 274294
rect 574488 274170 574558 274226
rect 574614 274170 574682 274226
rect 574738 274170 574808 274226
rect 574488 274102 574808 274170
rect 574488 274046 574558 274102
rect 574614 274046 574682 274102
rect 574738 274046 574808 274102
rect 574488 273978 574808 274046
rect 574488 273922 574558 273978
rect 574614 273922 574682 273978
rect 574738 273922 574808 273978
rect 574488 273888 574808 273922
rect 374808 262350 375128 262384
rect 374808 262294 374878 262350
rect 374934 262294 375002 262350
rect 375058 262294 375128 262350
rect 374808 262226 375128 262294
rect 374808 262170 374878 262226
rect 374934 262170 375002 262226
rect 375058 262170 375128 262226
rect 374808 262102 375128 262170
rect 374808 262046 374878 262102
rect 374934 262046 375002 262102
rect 375058 262046 375128 262102
rect 374808 261978 375128 262046
rect 374808 261922 374878 261978
rect 374934 261922 375002 261978
rect 375058 261922 375128 261978
rect 374808 261888 375128 261922
rect 405528 262350 405848 262384
rect 405528 262294 405598 262350
rect 405654 262294 405722 262350
rect 405778 262294 405848 262350
rect 405528 262226 405848 262294
rect 405528 262170 405598 262226
rect 405654 262170 405722 262226
rect 405778 262170 405848 262226
rect 405528 262102 405848 262170
rect 405528 262046 405598 262102
rect 405654 262046 405722 262102
rect 405778 262046 405848 262102
rect 405528 261978 405848 262046
rect 405528 261922 405598 261978
rect 405654 261922 405722 261978
rect 405778 261922 405848 261978
rect 405528 261888 405848 261922
rect 436248 262350 436568 262384
rect 436248 262294 436318 262350
rect 436374 262294 436442 262350
rect 436498 262294 436568 262350
rect 436248 262226 436568 262294
rect 436248 262170 436318 262226
rect 436374 262170 436442 262226
rect 436498 262170 436568 262226
rect 436248 262102 436568 262170
rect 436248 262046 436318 262102
rect 436374 262046 436442 262102
rect 436498 262046 436568 262102
rect 436248 261978 436568 262046
rect 436248 261922 436318 261978
rect 436374 261922 436442 261978
rect 436498 261922 436568 261978
rect 436248 261888 436568 261922
rect 466968 262350 467288 262384
rect 466968 262294 467038 262350
rect 467094 262294 467162 262350
rect 467218 262294 467288 262350
rect 466968 262226 467288 262294
rect 466968 262170 467038 262226
rect 467094 262170 467162 262226
rect 467218 262170 467288 262226
rect 466968 262102 467288 262170
rect 466968 262046 467038 262102
rect 467094 262046 467162 262102
rect 467218 262046 467288 262102
rect 466968 261978 467288 262046
rect 466968 261922 467038 261978
rect 467094 261922 467162 261978
rect 467218 261922 467288 261978
rect 466968 261888 467288 261922
rect 497688 262350 498008 262384
rect 497688 262294 497758 262350
rect 497814 262294 497882 262350
rect 497938 262294 498008 262350
rect 497688 262226 498008 262294
rect 497688 262170 497758 262226
rect 497814 262170 497882 262226
rect 497938 262170 498008 262226
rect 497688 262102 498008 262170
rect 497688 262046 497758 262102
rect 497814 262046 497882 262102
rect 497938 262046 498008 262102
rect 497688 261978 498008 262046
rect 497688 261922 497758 261978
rect 497814 261922 497882 261978
rect 497938 261922 498008 261978
rect 497688 261888 498008 261922
rect 528408 262350 528728 262384
rect 528408 262294 528478 262350
rect 528534 262294 528602 262350
rect 528658 262294 528728 262350
rect 528408 262226 528728 262294
rect 528408 262170 528478 262226
rect 528534 262170 528602 262226
rect 528658 262170 528728 262226
rect 528408 262102 528728 262170
rect 528408 262046 528478 262102
rect 528534 262046 528602 262102
rect 528658 262046 528728 262102
rect 528408 261978 528728 262046
rect 528408 261922 528478 261978
rect 528534 261922 528602 261978
rect 528658 261922 528728 261978
rect 528408 261888 528728 261922
rect 559128 262350 559448 262384
rect 559128 262294 559198 262350
rect 559254 262294 559322 262350
rect 559378 262294 559448 262350
rect 559128 262226 559448 262294
rect 559128 262170 559198 262226
rect 559254 262170 559322 262226
rect 559378 262170 559448 262226
rect 559128 262102 559448 262170
rect 559128 262046 559198 262102
rect 559254 262046 559322 262102
rect 559378 262046 559448 262102
rect 559128 261978 559448 262046
rect 559128 261922 559198 261978
rect 559254 261922 559322 261978
rect 559378 261922 559448 261978
rect 559128 261888 559448 261922
rect 359448 256350 359768 256384
rect 359448 256294 359518 256350
rect 359574 256294 359642 256350
rect 359698 256294 359768 256350
rect 359448 256226 359768 256294
rect 359448 256170 359518 256226
rect 359574 256170 359642 256226
rect 359698 256170 359768 256226
rect 359448 256102 359768 256170
rect 359448 256046 359518 256102
rect 359574 256046 359642 256102
rect 359698 256046 359768 256102
rect 359448 255978 359768 256046
rect 359448 255922 359518 255978
rect 359574 255922 359642 255978
rect 359698 255922 359768 255978
rect 359448 255888 359768 255922
rect 390168 256350 390488 256384
rect 390168 256294 390238 256350
rect 390294 256294 390362 256350
rect 390418 256294 390488 256350
rect 390168 256226 390488 256294
rect 390168 256170 390238 256226
rect 390294 256170 390362 256226
rect 390418 256170 390488 256226
rect 390168 256102 390488 256170
rect 390168 256046 390238 256102
rect 390294 256046 390362 256102
rect 390418 256046 390488 256102
rect 390168 255978 390488 256046
rect 390168 255922 390238 255978
rect 390294 255922 390362 255978
rect 390418 255922 390488 255978
rect 390168 255888 390488 255922
rect 420888 256350 421208 256384
rect 420888 256294 420958 256350
rect 421014 256294 421082 256350
rect 421138 256294 421208 256350
rect 420888 256226 421208 256294
rect 420888 256170 420958 256226
rect 421014 256170 421082 256226
rect 421138 256170 421208 256226
rect 420888 256102 421208 256170
rect 420888 256046 420958 256102
rect 421014 256046 421082 256102
rect 421138 256046 421208 256102
rect 420888 255978 421208 256046
rect 420888 255922 420958 255978
rect 421014 255922 421082 255978
rect 421138 255922 421208 255978
rect 420888 255888 421208 255922
rect 451608 256350 451928 256384
rect 451608 256294 451678 256350
rect 451734 256294 451802 256350
rect 451858 256294 451928 256350
rect 451608 256226 451928 256294
rect 451608 256170 451678 256226
rect 451734 256170 451802 256226
rect 451858 256170 451928 256226
rect 451608 256102 451928 256170
rect 451608 256046 451678 256102
rect 451734 256046 451802 256102
rect 451858 256046 451928 256102
rect 451608 255978 451928 256046
rect 451608 255922 451678 255978
rect 451734 255922 451802 255978
rect 451858 255922 451928 255978
rect 451608 255888 451928 255922
rect 482328 256350 482648 256384
rect 482328 256294 482398 256350
rect 482454 256294 482522 256350
rect 482578 256294 482648 256350
rect 482328 256226 482648 256294
rect 482328 256170 482398 256226
rect 482454 256170 482522 256226
rect 482578 256170 482648 256226
rect 482328 256102 482648 256170
rect 482328 256046 482398 256102
rect 482454 256046 482522 256102
rect 482578 256046 482648 256102
rect 482328 255978 482648 256046
rect 482328 255922 482398 255978
rect 482454 255922 482522 255978
rect 482578 255922 482648 255978
rect 482328 255888 482648 255922
rect 513048 256350 513368 256384
rect 513048 256294 513118 256350
rect 513174 256294 513242 256350
rect 513298 256294 513368 256350
rect 513048 256226 513368 256294
rect 513048 256170 513118 256226
rect 513174 256170 513242 256226
rect 513298 256170 513368 256226
rect 513048 256102 513368 256170
rect 513048 256046 513118 256102
rect 513174 256046 513242 256102
rect 513298 256046 513368 256102
rect 513048 255978 513368 256046
rect 513048 255922 513118 255978
rect 513174 255922 513242 255978
rect 513298 255922 513368 255978
rect 513048 255888 513368 255922
rect 543768 256350 544088 256384
rect 543768 256294 543838 256350
rect 543894 256294 543962 256350
rect 544018 256294 544088 256350
rect 543768 256226 544088 256294
rect 543768 256170 543838 256226
rect 543894 256170 543962 256226
rect 544018 256170 544088 256226
rect 543768 256102 544088 256170
rect 543768 256046 543838 256102
rect 543894 256046 543962 256102
rect 544018 256046 544088 256102
rect 543768 255978 544088 256046
rect 543768 255922 543838 255978
rect 543894 255922 543962 255978
rect 544018 255922 544088 255978
rect 543768 255888 544088 255922
rect 574488 256350 574808 256384
rect 574488 256294 574558 256350
rect 574614 256294 574682 256350
rect 574738 256294 574808 256350
rect 574488 256226 574808 256294
rect 574488 256170 574558 256226
rect 574614 256170 574682 256226
rect 574738 256170 574808 256226
rect 574488 256102 574808 256170
rect 574488 256046 574558 256102
rect 574614 256046 574682 256102
rect 574738 256046 574808 256102
rect 574488 255978 574808 256046
rect 574488 255922 574558 255978
rect 574614 255922 574682 255978
rect 574738 255922 574808 255978
rect 574488 255888 574808 255922
rect 374808 244350 375128 244384
rect 374808 244294 374878 244350
rect 374934 244294 375002 244350
rect 375058 244294 375128 244350
rect 374808 244226 375128 244294
rect 374808 244170 374878 244226
rect 374934 244170 375002 244226
rect 375058 244170 375128 244226
rect 374808 244102 375128 244170
rect 374808 244046 374878 244102
rect 374934 244046 375002 244102
rect 375058 244046 375128 244102
rect 374808 243978 375128 244046
rect 374808 243922 374878 243978
rect 374934 243922 375002 243978
rect 375058 243922 375128 243978
rect 374808 243888 375128 243922
rect 405528 244350 405848 244384
rect 405528 244294 405598 244350
rect 405654 244294 405722 244350
rect 405778 244294 405848 244350
rect 405528 244226 405848 244294
rect 405528 244170 405598 244226
rect 405654 244170 405722 244226
rect 405778 244170 405848 244226
rect 405528 244102 405848 244170
rect 405528 244046 405598 244102
rect 405654 244046 405722 244102
rect 405778 244046 405848 244102
rect 405528 243978 405848 244046
rect 405528 243922 405598 243978
rect 405654 243922 405722 243978
rect 405778 243922 405848 243978
rect 405528 243888 405848 243922
rect 436248 244350 436568 244384
rect 436248 244294 436318 244350
rect 436374 244294 436442 244350
rect 436498 244294 436568 244350
rect 436248 244226 436568 244294
rect 436248 244170 436318 244226
rect 436374 244170 436442 244226
rect 436498 244170 436568 244226
rect 436248 244102 436568 244170
rect 436248 244046 436318 244102
rect 436374 244046 436442 244102
rect 436498 244046 436568 244102
rect 436248 243978 436568 244046
rect 436248 243922 436318 243978
rect 436374 243922 436442 243978
rect 436498 243922 436568 243978
rect 436248 243888 436568 243922
rect 466968 244350 467288 244384
rect 466968 244294 467038 244350
rect 467094 244294 467162 244350
rect 467218 244294 467288 244350
rect 466968 244226 467288 244294
rect 466968 244170 467038 244226
rect 467094 244170 467162 244226
rect 467218 244170 467288 244226
rect 466968 244102 467288 244170
rect 466968 244046 467038 244102
rect 467094 244046 467162 244102
rect 467218 244046 467288 244102
rect 466968 243978 467288 244046
rect 466968 243922 467038 243978
rect 467094 243922 467162 243978
rect 467218 243922 467288 243978
rect 466968 243888 467288 243922
rect 497688 244350 498008 244384
rect 497688 244294 497758 244350
rect 497814 244294 497882 244350
rect 497938 244294 498008 244350
rect 497688 244226 498008 244294
rect 497688 244170 497758 244226
rect 497814 244170 497882 244226
rect 497938 244170 498008 244226
rect 497688 244102 498008 244170
rect 497688 244046 497758 244102
rect 497814 244046 497882 244102
rect 497938 244046 498008 244102
rect 497688 243978 498008 244046
rect 497688 243922 497758 243978
rect 497814 243922 497882 243978
rect 497938 243922 498008 243978
rect 497688 243888 498008 243922
rect 528408 244350 528728 244384
rect 528408 244294 528478 244350
rect 528534 244294 528602 244350
rect 528658 244294 528728 244350
rect 528408 244226 528728 244294
rect 528408 244170 528478 244226
rect 528534 244170 528602 244226
rect 528658 244170 528728 244226
rect 528408 244102 528728 244170
rect 528408 244046 528478 244102
rect 528534 244046 528602 244102
rect 528658 244046 528728 244102
rect 528408 243978 528728 244046
rect 528408 243922 528478 243978
rect 528534 243922 528602 243978
rect 528658 243922 528728 243978
rect 528408 243888 528728 243922
rect 559128 244350 559448 244384
rect 559128 244294 559198 244350
rect 559254 244294 559322 244350
rect 559378 244294 559448 244350
rect 559128 244226 559448 244294
rect 559128 244170 559198 244226
rect 559254 244170 559322 244226
rect 559378 244170 559448 244226
rect 559128 244102 559448 244170
rect 559128 244046 559198 244102
rect 559254 244046 559322 244102
rect 559378 244046 559448 244102
rect 559128 243978 559448 244046
rect 559128 243922 559198 243978
rect 559254 243922 559322 243978
rect 559378 243922 559448 243978
rect 559128 243888 559448 243922
rect 359448 238350 359768 238384
rect 359448 238294 359518 238350
rect 359574 238294 359642 238350
rect 359698 238294 359768 238350
rect 359448 238226 359768 238294
rect 359448 238170 359518 238226
rect 359574 238170 359642 238226
rect 359698 238170 359768 238226
rect 359448 238102 359768 238170
rect 359448 238046 359518 238102
rect 359574 238046 359642 238102
rect 359698 238046 359768 238102
rect 359448 237978 359768 238046
rect 359448 237922 359518 237978
rect 359574 237922 359642 237978
rect 359698 237922 359768 237978
rect 359448 237888 359768 237922
rect 390168 238350 390488 238384
rect 390168 238294 390238 238350
rect 390294 238294 390362 238350
rect 390418 238294 390488 238350
rect 390168 238226 390488 238294
rect 390168 238170 390238 238226
rect 390294 238170 390362 238226
rect 390418 238170 390488 238226
rect 390168 238102 390488 238170
rect 390168 238046 390238 238102
rect 390294 238046 390362 238102
rect 390418 238046 390488 238102
rect 390168 237978 390488 238046
rect 390168 237922 390238 237978
rect 390294 237922 390362 237978
rect 390418 237922 390488 237978
rect 390168 237888 390488 237922
rect 420888 238350 421208 238384
rect 420888 238294 420958 238350
rect 421014 238294 421082 238350
rect 421138 238294 421208 238350
rect 420888 238226 421208 238294
rect 420888 238170 420958 238226
rect 421014 238170 421082 238226
rect 421138 238170 421208 238226
rect 420888 238102 421208 238170
rect 420888 238046 420958 238102
rect 421014 238046 421082 238102
rect 421138 238046 421208 238102
rect 420888 237978 421208 238046
rect 420888 237922 420958 237978
rect 421014 237922 421082 237978
rect 421138 237922 421208 237978
rect 420888 237888 421208 237922
rect 451608 238350 451928 238384
rect 451608 238294 451678 238350
rect 451734 238294 451802 238350
rect 451858 238294 451928 238350
rect 451608 238226 451928 238294
rect 451608 238170 451678 238226
rect 451734 238170 451802 238226
rect 451858 238170 451928 238226
rect 451608 238102 451928 238170
rect 451608 238046 451678 238102
rect 451734 238046 451802 238102
rect 451858 238046 451928 238102
rect 451608 237978 451928 238046
rect 451608 237922 451678 237978
rect 451734 237922 451802 237978
rect 451858 237922 451928 237978
rect 451608 237888 451928 237922
rect 482328 238350 482648 238384
rect 482328 238294 482398 238350
rect 482454 238294 482522 238350
rect 482578 238294 482648 238350
rect 482328 238226 482648 238294
rect 482328 238170 482398 238226
rect 482454 238170 482522 238226
rect 482578 238170 482648 238226
rect 482328 238102 482648 238170
rect 482328 238046 482398 238102
rect 482454 238046 482522 238102
rect 482578 238046 482648 238102
rect 482328 237978 482648 238046
rect 482328 237922 482398 237978
rect 482454 237922 482522 237978
rect 482578 237922 482648 237978
rect 482328 237888 482648 237922
rect 513048 238350 513368 238384
rect 513048 238294 513118 238350
rect 513174 238294 513242 238350
rect 513298 238294 513368 238350
rect 513048 238226 513368 238294
rect 513048 238170 513118 238226
rect 513174 238170 513242 238226
rect 513298 238170 513368 238226
rect 513048 238102 513368 238170
rect 513048 238046 513118 238102
rect 513174 238046 513242 238102
rect 513298 238046 513368 238102
rect 513048 237978 513368 238046
rect 513048 237922 513118 237978
rect 513174 237922 513242 237978
rect 513298 237922 513368 237978
rect 513048 237888 513368 237922
rect 543768 238350 544088 238384
rect 543768 238294 543838 238350
rect 543894 238294 543962 238350
rect 544018 238294 544088 238350
rect 543768 238226 544088 238294
rect 543768 238170 543838 238226
rect 543894 238170 543962 238226
rect 544018 238170 544088 238226
rect 543768 238102 544088 238170
rect 543768 238046 543838 238102
rect 543894 238046 543962 238102
rect 544018 238046 544088 238102
rect 543768 237978 544088 238046
rect 543768 237922 543838 237978
rect 543894 237922 543962 237978
rect 544018 237922 544088 237978
rect 543768 237888 544088 237922
rect 574488 238350 574808 238384
rect 574488 238294 574558 238350
rect 574614 238294 574682 238350
rect 574738 238294 574808 238350
rect 574488 238226 574808 238294
rect 574488 238170 574558 238226
rect 574614 238170 574682 238226
rect 574738 238170 574808 238226
rect 574488 238102 574808 238170
rect 574488 238046 574558 238102
rect 574614 238046 574682 238102
rect 574738 238046 574808 238102
rect 574488 237978 574808 238046
rect 574488 237922 574558 237978
rect 574614 237922 574682 237978
rect 574738 237922 574808 237978
rect 574488 237888 574808 237922
rect 374808 226350 375128 226384
rect 374808 226294 374878 226350
rect 374934 226294 375002 226350
rect 375058 226294 375128 226350
rect 374808 226226 375128 226294
rect 374808 226170 374878 226226
rect 374934 226170 375002 226226
rect 375058 226170 375128 226226
rect 374808 226102 375128 226170
rect 374808 226046 374878 226102
rect 374934 226046 375002 226102
rect 375058 226046 375128 226102
rect 374808 225978 375128 226046
rect 374808 225922 374878 225978
rect 374934 225922 375002 225978
rect 375058 225922 375128 225978
rect 374808 225888 375128 225922
rect 405528 226350 405848 226384
rect 405528 226294 405598 226350
rect 405654 226294 405722 226350
rect 405778 226294 405848 226350
rect 405528 226226 405848 226294
rect 405528 226170 405598 226226
rect 405654 226170 405722 226226
rect 405778 226170 405848 226226
rect 405528 226102 405848 226170
rect 405528 226046 405598 226102
rect 405654 226046 405722 226102
rect 405778 226046 405848 226102
rect 405528 225978 405848 226046
rect 405528 225922 405598 225978
rect 405654 225922 405722 225978
rect 405778 225922 405848 225978
rect 405528 225888 405848 225922
rect 436248 226350 436568 226384
rect 436248 226294 436318 226350
rect 436374 226294 436442 226350
rect 436498 226294 436568 226350
rect 436248 226226 436568 226294
rect 436248 226170 436318 226226
rect 436374 226170 436442 226226
rect 436498 226170 436568 226226
rect 436248 226102 436568 226170
rect 436248 226046 436318 226102
rect 436374 226046 436442 226102
rect 436498 226046 436568 226102
rect 436248 225978 436568 226046
rect 436248 225922 436318 225978
rect 436374 225922 436442 225978
rect 436498 225922 436568 225978
rect 436248 225888 436568 225922
rect 466968 226350 467288 226384
rect 466968 226294 467038 226350
rect 467094 226294 467162 226350
rect 467218 226294 467288 226350
rect 466968 226226 467288 226294
rect 466968 226170 467038 226226
rect 467094 226170 467162 226226
rect 467218 226170 467288 226226
rect 466968 226102 467288 226170
rect 466968 226046 467038 226102
rect 467094 226046 467162 226102
rect 467218 226046 467288 226102
rect 466968 225978 467288 226046
rect 466968 225922 467038 225978
rect 467094 225922 467162 225978
rect 467218 225922 467288 225978
rect 466968 225888 467288 225922
rect 497688 226350 498008 226384
rect 497688 226294 497758 226350
rect 497814 226294 497882 226350
rect 497938 226294 498008 226350
rect 497688 226226 498008 226294
rect 497688 226170 497758 226226
rect 497814 226170 497882 226226
rect 497938 226170 498008 226226
rect 497688 226102 498008 226170
rect 497688 226046 497758 226102
rect 497814 226046 497882 226102
rect 497938 226046 498008 226102
rect 497688 225978 498008 226046
rect 497688 225922 497758 225978
rect 497814 225922 497882 225978
rect 497938 225922 498008 225978
rect 497688 225888 498008 225922
rect 528408 226350 528728 226384
rect 528408 226294 528478 226350
rect 528534 226294 528602 226350
rect 528658 226294 528728 226350
rect 528408 226226 528728 226294
rect 528408 226170 528478 226226
rect 528534 226170 528602 226226
rect 528658 226170 528728 226226
rect 528408 226102 528728 226170
rect 528408 226046 528478 226102
rect 528534 226046 528602 226102
rect 528658 226046 528728 226102
rect 528408 225978 528728 226046
rect 528408 225922 528478 225978
rect 528534 225922 528602 225978
rect 528658 225922 528728 225978
rect 528408 225888 528728 225922
rect 559128 226350 559448 226384
rect 559128 226294 559198 226350
rect 559254 226294 559322 226350
rect 559378 226294 559448 226350
rect 559128 226226 559448 226294
rect 559128 226170 559198 226226
rect 559254 226170 559322 226226
rect 559378 226170 559448 226226
rect 559128 226102 559448 226170
rect 559128 226046 559198 226102
rect 559254 226046 559322 226102
rect 559378 226046 559448 226102
rect 559128 225978 559448 226046
rect 559128 225922 559198 225978
rect 559254 225922 559322 225978
rect 559378 225922 559448 225978
rect 559128 225888 559448 225922
rect 359448 220350 359768 220384
rect 359448 220294 359518 220350
rect 359574 220294 359642 220350
rect 359698 220294 359768 220350
rect 359448 220226 359768 220294
rect 359448 220170 359518 220226
rect 359574 220170 359642 220226
rect 359698 220170 359768 220226
rect 359448 220102 359768 220170
rect 359448 220046 359518 220102
rect 359574 220046 359642 220102
rect 359698 220046 359768 220102
rect 359448 219978 359768 220046
rect 359448 219922 359518 219978
rect 359574 219922 359642 219978
rect 359698 219922 359768 219978
rect 359448 219888 359768 219922
rect 390168 220350 390488 220384
rect 390168 220294 390238 220350
rect 390294 220294 390362 220350
rect 390418 220294 390488 220350
rect 390168 220226 390488 220294
rect 390168 220170 390238 220226
rect 390294 220170 390362 220226
rect 390418 220170 390488 220226
rect 390168 220102 390488 220170
rect 390168 220046 390238 220102
rect 390294 220046 390362 220102
rect 390418 220046 390488 220102
rect 390168 219978 390488 220046
rect 390168 219922 390238 219978
rect 390294 219922 390362 219978
rect 390418 219922 390488 219978
rect 390168 219888 390488 219922
rect 420888 220350 421208 220384
rect 420888 220294 420958 220350
rect 421014 220294 421082 220350
rect 421138 220294 421208 220350
rect 420888 220226 421208 220294
rect 420888 220170 420958 220226
rect 421014 220170 421082 220226
rect 421138 220170 421208 220226
rect 420888 220102 421208 220170
rect 420888 220046 420958 220102
rect 421014 220046 421082 220102
rect 421138 220046 421208 220102
rect 420888 219978 421208 220046
rect 420888 219922 420958 219978
rect 421014 219922 421082 219978
rect 421138 219922 421208 219978
rect 420888 219888 421208 219922
rect 451608 220350 451928 220384
rect 451608 220294 451678 220350
rect 451734 220294 451802 220350
rect 451858 220294 451928 220350
rect 451608 220226 451928 220294
rect 451608 220170 451678 220226
rect 451734 220170 451802 220226
rect 451858 220170 451928 220226
rect 451608 220102 451928 220170
rect 451608 220046 451678 220102
rect 451734 220046 451802 220102
rect 451858 220046 451928 220102
rect 451608 219978 451928 220046
rect 451608 219922 451678 219978
rect 451734 219922 451802 219978
rect 451858 219922 451928 219978
rect 451608 219888 451928 219922
rect 482328 220350 482648 220384
rect 482328 220294 482398 220350
rect 482454 220294 482522 220350
rect 482578 220294 482648 220350
rect 482328 220226 482648 220294
rect 482328 220170 482398 220226
rect 482454 220170 482522 220226
rect 482578 220170 482648 220226
rect 482328 220102 482648 220170
rect 482328 220046 482398 220102
rect 482454 220046 482522 220102
rect 482578 220046 482648 220102
rect 482328 219978 482648 220046
rect 482328 219922 482398 219978
rect 482454 219922 482522 219978
rect 482578 219922 482648 219978
rect 482328 219888 482648 219922
rect 513048 220350 513368 220384
rect 513048 220294 513118 220350
rect 513174 220294 513242 220350
rect 513298 220294 513368 220350
rect 513048 220226 513368 220294
rect 513048 220170 513118 220226
rect 513174 220170 513242 220226
rect 513298 220170 513368 220226
rect 513048 220102 513368 220170
rect 513048 220046 513118 220102
rect 513174 220046 513242 220102
rect 513298 220046 513368 220102
rect 513048 219978 513368 220046
rect 513048 219922 513118 219978
rect 513174 219922 513242 219978
rect 513298 219922 513368 219978
rect 513048 219888 513368 219922
rect 543768 220350 544088 220384
rect 543768 220294 543838 220350
rect 543894 220294 543962 220350
rect 544018 220294 544088 220350
rect 543768 220226 544088 220294
rect 543768 220170 543838 220226
rect 543894 220170 543962 220226
rect 544018 220170 544088 220226
rect 543768 220102 544088 220170
rect 543768 220046 543838 220102
rect 543894 220046 543962 220102
rect 544018 220046 544088 220102
rect 543768 219978 544088 220046
rect 543768 219922 543838 219978
rect 543894 219922 543962 219978
rect 544018 219922 544088 219978
rect 543768 219888 544088 219922
rect 574488 220350 574808 220384
rect 574488 220294 574558 220350
rect 574614 220294 574682 220350
rect 574738 220294 574808 220350
rect 574488 220226 574808 220294
rect 574488 220170 574558 220226
rect 574614 220170 574682 220226
rect 574738 220170 574808 220226
rect 574488 220102 574808 220170
rect 574488 220046 574558 220102
rect 574614 220046 574682 220102
rect 574738 220046 574808 220102
rect 574488 219978 574808 220046
rect 574488 219922 574558 219978
rect 574614 219922 574682 219978
rect 574738 219922 574808 219978
rect 574488 219888 574808 219922
rect 356748 164948 356804 213542
rect 374808 208350 375128 208384
rect 374808 208294 374878 208350
rect 374934 208294 375002 208350
rect 375058 208294 375128 208350
rect 374808 208226 375128 208294
rect 374808 208170 374878 208226
rect 374934 208170 375002 208226
rect 375058 208170 375128 208226
rect 374808 208102 375128 208170
rect 374808 208046 374878 208102
rect 374934 208046 375002 208102
rect 375058 208046 375128 208102
rect 374808 207978 375128 208046
rect 374808 207922 374878 207978
rect 374934 207922 375002 207978
rect 375058 207922 375128 207978
rect 374808 207888 375128 207922
rect 405528 208350 405848 208384
rect 405528 208294 405598 208350
rect 405654 208294 405722 208350
rect 405778 208294 405848 208350
rect 405528 208226 405848 208294
rect 405528 208170 405598 208226
rect 405654 208170 405722 208226
rect 405778 208170 405848 208226
rect 405528 208102 405848 208170
rect 405528 208046 405598 208102
rect 405654 208046 405722 208102
rect 405778 208046 405848 208102
rect 405528 207978 405848 208046
rect 405528 207922 405598 207978
rect 405654 207922 405722 207978
rect 405778 207922 405848 207978
rect 405528 207888 405848 207922
rect 436248 208350 436568 208384
rect 436248 208294 436318 208350
rect 436374 208294 436442 208350
rect 436498 208294 436568 208350
rect 436248 208226 436568 208294
rect 436248 208170 436318 208226
rect 436374 208170 436442 208226
rect 436498 208170 436568 208226
rect 436248 208102 436568 208170
rect 436248 208046 436318 208102
rect 436374 208046 436442 208102
rect 436498 208046 436568 208102
rect 436248 207978 436568 208046
rect 436248 207922 436318 207978
rect 436374 207922 436442 207978
rect 436498 207922 436568 207978
rect 436248 207888 436568 207922
rect 466968 208350 467288 208384
rect 466968 208294 467038 208350
rect 467094 208294 467162 208350
rect 467218 208294 467288 208350
rect 466968 208226 467288 208294
rect 466968 208170 467038 208226
rect 467094 208170 467162 208226
rect 467218 208170 467288 208226
rect 466968 208102 467288 208170
rect 466968 208046 467038 208102
rect 467094 208046 467162 208102
rect 467218 208046 467288 208102
rect 466968 207978 467288 208046
rect 466968 207922 467038 207978
rect 467094 207922 467162 207978
rect 467218 207922 467288 207978
rect 466968 207888 467288 207922
rect 497688 208350 498008 208384
rect 497688 208294 497758 208350
rect 497814 208294 497882 208350
rect 497938 208294 498008 208350
rect 497688 208226 498008 208294
rect 497688 208170 497758 208226
rect 497814 208170 497882 208226
rect 497938 208170 498008 208226
rect 497688 208102 498008 208170
rect 497688 208046 497758 208102
rect 497814 208046 497882 208102
rect 497938 208046 498008 208102
rect 497688 207978 498008 208046
rect 497688 207922 497758 207978
rect 497814 207922 497882 207978
rect 497938 207922 498008 207978
rect 497688 207888 498008 207922
rect 528408 208350 528728 208384
rect 528408 208294 528478 208350
rect 528534 208294 528602 208350
rect 528658 208294 528728 208350
rect 528408 208226 528728 208294
rect 528408 208170 528478 208226
rect 528534 208170 528602 208226
rect 528658 208170 528728 208226
rect 528408 208102 528728 208170
rect 528408 208046 528478 208102
rect 528534 208046 528602 208102
rect 528658 208046 528728 208102
rect 528408 207978 528728 208046
rect 528408 207922 528478 207978
rect 528534 207922 528602 207978
rect 528658 207922 528728 207978
rect 528408 207888 528728 207922
rect 559128 208350 559448 208384
rect 559128 208294 559198 208350
rect 559254 208294 559322 208350
rect 559378 208294 559448 208350
rect 559128 208226 559448 208294
rect 559128 208170 559198 208226
rect 559254 208170 559322 208226
rect 559378 208170 559448 208226
rect 559128 208102 559448 208170
rect 559128 208046 559198 208102
rect 559254 208046 559322 208102
rect 559378 208046 559448 208102
rect 559128 207978 559448 208046
rect 559128 207922 559198 207978
rect 559254 207922 559322 207978
rect 559378 207922 559448 207978
rect 559128 207888 559448 207922
rect 359448 202350 359768 202384
rect 359448 202294 359518 202350
rect 359574 202294 359642 202350
rect 359698 202294 359768 202350
rect 359448 202226 359768 202294
rect 359448 202170 359518 202226
rect 359574 202170 359642 202226
rect 359698 202170 359768 202226
rect 359448 202102 359768 202170
rect 359448 202046 359518 202102
rect 359574 202046 359642 202102
rect 359698 202046 359768 202102
rect 359448 201978 359768 202046
rect 359448 201922 359518 201978
rect 359574 201922 359642 201978
rect 359698 201922 359768 201978
rect 359448 201888 359768 201922
rect 390168 202350 390488 202384
rect 390168 202294 390238 202350
rect 390294 202294 390362 202350
rect 390418 202294 390488 202350
rect 390168 202226 390488 202294
rect 390168 202170 390238 202226
rect 390294 202170 390362 202226
rect 390418 202170 390488 202226
rect 390168 202102 390488 202170
rect 390168 202046 390238 202102
rect 390294 202046 390362 202102
rect 390418 202046 390488 202102
rect 390168 201978 390488 202046
rect 390168 201922 390238 201978
rect 390294 201922 390362 201978
rect 390418 201922 390488 201978
rect 390168 201888 390488 201922
rect 420888 202350 421208 202384
rect 420888 202294 420958 202350
rect 421014 202294 421082 202350
rect 421138 202294 421208 202350
rect 420888 202226 421208 202294
rect 420888 202170 420958 202226
rect 421014 202170 421082 202226
rect 421138 202170 421208 202226
rect 420888 202102 421208 202170
rect 420888 202046 420958 202102
rect 421014 202046 421082 202102
rect 421138 202046 421208 202102
rect 420888 201978 421208 202046
rect 420888 201922 420958 201978
rect 421014 201922 421082 201978
rect 421138 201922 421208 201978
rect 420888 201888 421208 201922
rect 451608 202350 451928 202384
rect 451608 202294 451678 202350
rect 451734 202294 451802 202350
rect 451858 202294 451928 202350
rect 451608 202226 451928 202294
rect 451608 202170 451678 202226
rect 451734 202170 451802 202226
rect 451858 202170 451928 202226
rect 451608 202102 451928 202170
rect 451608 202046 451678 202102
rect 451734 202046 451802 202102
rect 451858 202046 451928 202102
rect 451608 201978 451928 202046
rect 451608 201922 451678 201978
rect 451734 201922 451802 201978
rect 451858 201922 451928 201978
rect 451608 201888 451928 201922
rect 482328 202350 482648 202384
rect 482328 202294 482398 202350
rect 482454 202294 482522 202350
rect 482578 202294 482648 202350
rect 482328 202226 482648 202294
rect 482328 202170 482398 202226
rect 482454 202170 482522 202226
rect 482578 202170 482648 202226
rect 482328 202102 482648 202170
rect 482328 202046 482398 202102
rect 482454 202046 482522 202102
rect 482578 202046 482648 202102
rect 482328 201978 482648 202046
rect 482328 201922 482398 201978
rect 482454 201922 482522 201978
rect 482578 201922 482648 201978
rect 482328 201888 482648 201922
rect 513048 202350 513368 202384
rect 513048 202294 513118 202350
rect 513174 202294 513242 202350
rect 513298 202294 513368 202350
rect 513048 202226 513368 202294
rect 513048 202170 513118 202226
rect 513174 202170 513242 202226
rect 513298 202170 513368 202226
rect 513048 202102 513368 202170
rect 513048 202046 513118 202102
rect 513174 202046 513242 202102
rect 513298 202046 513368 202102
rect 513048 201978 513368 202046
rect 513048 201922 513118 201978
rect 513174 201922 513242 201978
rect 513298 201922 513368 201978
rect 513048 201888 513368 201922
rect 543768 202350 544088 202384
rect 543768 202294 543838 202350
rect 543894 202294 543962 202350
rect 544018 202294 544088 202350
rect 543768 202226 544088 202294
rect 543768 202170 543838 202226
rect 543894 202170 543962 202226
rect 544018 202170 544088 202226
rect 543768 202102 544088 202170
rect 543768 202046 543838 202102
rect 543894 202046 543962 202102
rect 544018 202046 544088 202102
rect 543768 201978 544088 202046
rect 543768 201922 543838 201978
rect 543894 201922 543962 201978
rect 544018 201922 544088 201978
rect 543768 201888 544088 201922
rect 574488 202350 574808 202384
rect 574488 202294 574558 202350
rect 574614 202294 574682 202350
rect 574738 202294 574808 202350
rect 574488 202226 574808 202294
rect 574488 202170 574558 202226
rect 574614 202170 574682 202226
rect 574738 202170 574808 202226
rect 574488 202102 574808 202170
rect 574488 202046 574558 202102
rect 574614 202046 574682 202102
rect 574738 202046 574808 202102
rect 574488 201978 574808 202046
rect 574488 201922 574558 201978
rect 574614 201922 574682 201978
rect 574738 201922 574808 201978
rect 574488 201888 574808 201922
rect 374808 190350 375128 190384
rect 374808 190294 374878 190350
rect 374934 190294 375002 190350
rect 375058 190294 375128 190350
rect 374808 190226 375128 190294
rect 374808 190170 374878 190226
rect 374934 190170 375002 190226
rect 375058 190170 375128 190226
rect 374808 190102 375128 190170
rect 374808 190046 374878 190102
rect 374934 190046 375002 190102
rect 375058 190046 375128 190102
rect 374808 189978 375128 190046
rect 374808 189922 374878 189978
rect 374934 189922 375002 189978
rect 375058 189922 375128 189978
rect 374808 189888 375128 189922
rect 405528 190350 405848 190384
rect 405528 190294 405598 190350
rect 405654 190294 405722 190350
rect 405778 190294 405848 190350
rect 405528 190226 405848 190294
rect 405528 190170 405598 190226
rect 405654 190170 405722 190226
rect 405778 190170 405848 190226
rect 405528 190102 405848 190170
rect 405528 190046 405598 190102
rect 405654 190046 405722 190102
rect 405778 190046 405848 190102
rect 405528 189978 405848 190046
rect 405528 189922 405598 189978
rect 405654 189922 405722 189978
rect 405778 189922 405848 189978
rect 405528 189888 405848 189922
rect 436248 190350 436568 190384
rect 436248 190294 436318 190350
rect 436374 190294 436442 190350
rect 436498 190294 436568 190350
rect 436248 190226 436568 190294
rect 436248 190170 436318 190226
rect 436374 190170 436442 190226
rect 436498 190170 436568 190226
rect 436248 190102 436568 190170
rect 436248 190046 436318 190102
rect 436374 190046 436442 190102
rect 436498 190046 436568 190102
rect 436248 189978 436568 190046
rect 436248 189922 436318 189978
rect 436374 189922 436442 189978
rect 436498 189922 436568 189978
rect 436248 189888 436568 189922
rect 466968 190350 467288 190384
rect 466968 190294 467038 190350
rect 467094 190294 467162 190350
rect 467218 190294 467288 190350
rect 466968 190226 467288 190294
rect 466968 190170 467038 190226
rect 467094 190170 467162 190226
rect 467218 190170 467288 190226
rect 466968 190102 467288 190170
rect 466968 190046 467038 190102
rect 467094 190046 467162 190102
rect 467218 190046 467288 190102
rect 466968 189978 467288 190046
rect 466968 189922 467038 189978
rect 467094 189922 467162 189978
rect 467218 189922 467288 189978
rect 466968 189888 467288 189922
rect 497688 190350 498008 190384
rect 497688 190294 497758 190350
rect 497814 190294 497882 190350
rect 497938 190294 498008 190350
rect 497688 190226 498008 190294
rect 497688 190170 497758 190226
rect 497814 190170 497882 190226
rect 497938 190170 498008 190226
rect 497688 190102 498008 190170
rect 497688 190046 497758 190102
rect 497814 190046 497882 190102
rect 497938 190046 498008 190102
rect 497688 189978 498008 190046
rect 497688 189922 497758 189978
rect 497814 189922 497882 189978
rect 497938 189922 498008 189978
rect 497688 189888 498008 189922
rect 528408 190350 528728 190384
rect 528408 190294 528478 190350
rect 528534 190294 528602 190350
rect 528658 190294 528728 190350
rect 528408 190226 528728 190294
rect 528408 190170 528478 190226
rect 528534 190170 528602 190226
rect 528658 190170 528728 190226
rect 528408 190102 528728 190170
rect 528408 190046 528478 190102
rect 528534 190046 528602 190102
rect 528658 190046 528728 190102
rect 528408 189978 528728 190046
rect 528408 189922 528478 189978
rect 528534 189922 528602 189978
rect 528658 189922 528728 189978
rect 528408 189888 528728 189922
rect 559128 190350 559448 190384
rect 559128 190294 559198 190350
rect 559254 190294 559322 190350
rect 559378 190294 559448 190350
rect 559128 190226 559448 190294
rect 559128 190170 559198 190226
rect 559254 190170 559322 190226
rect 559378 190170 559448 190226
rect 559128 190102 559448 190170
rect 559128 190046 559198 190102
rect 559254 190046 559322 190102
rect 559378 190046 559448 190102
rect 559128 189978 559448 190046
rect 559128 189922 559198 189978
rect 559254 189922 559322 189978
rect 559378 189922 559448 189978
rect 559128 189888 559448 189922
rect 359448 184350 359768 184384
rect 359448 184294 359518 184350
rect 359574 184294 359642 184350
rect 359698 184294 359768 184350
rect 359448 184226 359768 184294
rect 359448 184170 359518 184226
rect 359574 184170 359642 184226
rect 359698 184170 359768 184226
rect 359448 184102 359768 184170
rect 359448 184046 359518 184102
rect 359574 184046 359642 184102
rect 359698 184046 359768 184102
rect 359448 183978 359768 184046
rect 359448 183922 359518 183978
rect 359574 183922 359642 183978
rect 359698 183922 359768 183978
rect 359448 183888 359768 183922
rect 390168 184350 390488 184384
rect 390168 184294 390238 184350
rect 390294 184294 390362 184350
rect 390418 184294 390488 184350
rect 390168 184226 390488 184294
rect 390168 184170 390238 184226
rect 390294 184170 390362 184226
rect 390418 184170 390488 184226
rect 390168 184102 390488 184170
rect 390168 184046 390238 184102
rect 390294 184046 390362 184102
rect 390418 184046 390488 184102
rect 390168 183978 390488 184046
rect 390168 183922 390238 183978
rect 390294 183922 390362 183978
rect 390418 183922 390488 183978
rect 390168 183888 390488 183922
rect 420888 184350 421208 184384
rect 420888 184294 420958 184350
rect 421014 184294 421082 184350
rect 421138 184294 421208 184350
rect 420888 184226 421208 184294
rect 420888 184170 420958 184226
rect 421014 184170 421082 184226
rect 421138 184170 421208 184226
rect 420888 184102 421208 184170
rect 420888 184046 420958 184102
rect 421014 184046 421082 184102
rect 421138 184046 421208 184102
rect 420888 183978 421208 184046
rect 420888 183922 420958 183978
rect 421014 183922 421082 183978
rect 421138 183922 421208 183978
rect 420888 183888 421208 183922
rect 451608 184350 451928 184384
rect 451608 184294 451678 184350
rect 451734 184294 451802 184350
rect 451858 184294 451928 184350
rect 451608 184226 451928 184294
rect 451608 184170 451678 184226
rect 451734 184170 451802 184226
rect 451858 184170 451928 184226
rect 451608 184102 451928 184170
rect 451608 184046 451678 184102
rect 451734 184046 451802 184102
rect 451858 184046 451928 184102
rect 451608 183978 451928 184046
rect 451608 183922 451678 183978
rect 451734 183922 451802 183978
rect 451858 183922 451928 183978
rect 451608 183888 451928 183922
rect 482328 184350 482648 184384
rect 482328 184294 482398 184350
rect 482454 184294 482522 184350
rect 482578 184294 482648 184350
rect 482328 184226 482648 184294
rect 482328 184170 482398 184226
rect 482454 184170 482522 184226
rect 482578 184170 482648 184226
rect 482328 184102 482648 184170
rect 482328 184046 482398 184102
rect 482454 184046 482522 184102
rect 482578 184046 482648 184102
rect 482328 183978 482648 184046
rect 482328 183922 482398 183978
rect 482454 183922 482522 183978
rect 482578 183922 482648 183978
rect 482328 183888 482648 183922
rect 513048 184350 513368 184384
rect 513048 184294 513118 184350
rect 513174 184294 513242 184350
rect 513298 184294 513368 184350
rect 513048 184226 513368 184294
rect 513048 184170 513118 184226
rect 513174 184170 513242 184226
rect 513298 184170 513368 184226
rect 513048 184102 513368 184170
rect 513048 184046 513118 184102
rect 513174 184046 513242 184102
rect 513298 184046 513368 184102
rect 513048 183978 513368 184046
rect 513048 183922 513118 183978
rect 513174 183922 513242 183978
rect 513298 183922 513368 183978
rect 513048 183888 513368 183922
rect 543768 184350 544088 184384
rect 543768 184294 543838 184350
rect 543894 184294 543962 184350
rect 544018 184294 544088 184350
rect 543768 184226 544088 184294
rect 543768 184170 543838 184226
rect 543894 184170 543962 184226
rect 544018 184170 544088 184226
rect 543768 184102 544088 184170
rect 543768 184046 543838 184102
rect 543894 184046 543962 184102
rect 544018 184046 544088 184102
rect 543768 183978 544088 184046
rect 543768 183922 543838 183978
rect 543894 183922 543962 183978
rect 544018 183922 544088 183978
rect 543768 183888 544088 183922
rect 574488 184350 574808 184384
rect 574488 184294 574558 184350
rect 574614 184294 574682 184350
rect 574738 184294 574808 184350
rect 574488 184226 574808 184294
rect 574488 184170 574558 184226
rect 574614 184170 574682 184226
rect 574738 184170 574808 184226
rect 574488 184102 574808 184170
rect 574488 184046 574558 184102
rect 574614 184046 574682 184102
rect 574738 184046 574808 184102
rect 574488 183978 574808 184046
rect 574488 183922 574558 183978
rect 574614 183922 574682 183978
rect 574738 183922 574808 183978
rect 574488 183888 574808 183922
rect 374808 172350 375128 172384
rect 374808 172294 374878 172350
rect 374934 172294 375002 172350
rect 375058 172294 375128 172350
rect 374808 172226 375128 172294
rect 374808 172170 374878 172226
rect 374934 172170 375002 172226
rect 375058 172170 375128 172226
rect 374808 172102 375128 172170
rect 374808 172046 374878 172102
rect 374934 172046 375002 172102
rect 375058 172046 375128 172102
rect 374808 171978 375128 172046
rect 374808 171922 374878 171978
rect 374934 171922 375002 171978
rect 375058 171922 375128 171978
rect 374808 171888 375128 171922
rect 405528 172350 405848 172384
rect 405528 172294 405598 172350
rect 405654 172294 405722 172350
rect 405778 172294 405848 172350
rect 405528 172226 405848 172294
rect 405528 172170 405598 172226
rect 405654 172170 405722 172226
rect 405778 172170 405848 172226
rect 405528 172102 405848 172170
rect 405528 172046 405598 172102
rect 405654 172046 405722 172102
rect 405778 172046 405848 172102
rect 405528 171978 405848 172046
rect 405528 171922 405598 171978
rect 405654 171922 405722 171978
rect 405778 171922 405848 171978
rect 405528 171888 405848 171922
rect 436248 172350 436568 172384
rect 436248 172294 436318 172350
rect 436374 172294 436442 172350
rect 436498 172294 436568 172350
rect 436248 172226 436568 172294
rect 436248 172170 436318 172226
rect 436374 172170 436442 172226
rect 436498 172170 436568 172226
rect 436248 172102 436568 172170
rect 436248 172046 436318 172102
rect 436374 172046 436442 172102
rect 436498 172046 436568 172102
rect 436248 171978 436568 172046
rect 436248 171922 436318 171978
rect 436374 171922 436442 171978
rect 436498 171922 436568 171978
rect 436248 171888 436568 171922
rect 466968 172350 467288 172384
rect 466968 172294 467038 172350
rect 467094 172294 467162 172350
rect 467218 172294 467288 172350
rect 466968 172226 467288 172294
rect 466968 172170 467038 172226
rect 467094 172170 467162 172226
rect 467218 172170 467288 172226
rect 466968 172102 467288 172170
rect 466968 172046 467038 172102
rect 467094 172046 467162 172102
rect 467218 172046 467288 172102
rect 466968 171978 467288 172046
rect 466968 171922 467038 171978
rect 467094 171922 467162 171978
rect 467218 171922 467288 171978
rect 466968 171888 467288 171922
rect 497688 172350 498008 172384
rect 497688 172294 497758 172350
rect 497814 172294 497882 172350
rect 497938 172294 498008 172350
rect 497688 172226 498008 172294
rect 497688 172170 497758 172226
rect 497814 172170 497882 172226
rect 497938 172170 498008 172226
rect 497688 172102 498008 172170
rect 497688 172046 497758 172102
rect 497814 172046 497882 172102
rect 497938 172046 498008 172102
rect 497688 171978 498008 172046
rect 497688 171922 497758 171978
rect 497814 171922 497882 171978
rect 497938 171922 498008 171978
rect 497688 171888 498008 171922
rect 528408 172350 528728 172384
rect 528408 172294 528478 172350
rect 528534 172294 528602 172350
rect 528658 172294 528728 172350
rect 528408 172226 528728 172294
rect 528408 172170 528478 172226
rect 528534 172170 528602 172226
rect 528658 172170 528728 172226
rect 528408 172102 528728 172170
rect 528408 172046 528478 172102
rect 528534 172046 528602 172102
rect 528658 172046 528728 172102
rect 528408 171978 528728 172046
rect 528408 171922 528478 171978
rect 528534 171922 528602 171978
rect 528658 171922 528728 171978
rect 528408 171888 528728 171922
rect 559128 172350 559448 172384
rect 559128 172294 559198 172350
rect 559254 172294 559322 172350
rect 559378 172294 559448 172350
rect 559128 172226 559448 172294
rect 559128 172170 559198 172226
rect 559254 172170 559322 172226
rect 559378 172170 559448 172226
rect 559128 172102 559448 172170
rect 559128 172046 559198 172102
rect 559254 172046 559322 172102
rect 559378 172046 559448 172102
rect 559128 171978 559448 172046
rect 559128 171922 559198 171978
rect 559254 171922 559322 171978
rect 559378 171922 559448 171978
rect 559128 171888 559448 171922
rect 356748 164882 356804 164892
rect 488908 165538 488964 165548
rect 457884 164836 457940 164846
rect 374058 148350 374678 164250
rect 374058 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 374678 148350
rect 374058 148226 374678 148294
rect 374058 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 374678 148226
rect 374058 148102 374678 148170
rect 374058 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 374678 148102
rect 374058 147978 374678 148046
rect 374058 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 374678 147978
rect 366268 145918 366324 145946
rect 366268 145842 366324 145852
rect 374058 130350 374678 147922
rect 374058 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 374678 130350
rect 374058 130226 374678 130294
rect 374058 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 374678 130226
rect 374058 130102 374678 130170
rect 374058 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 374678 130102
rect 374058 129978 374678 130046
rect 374058 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 374678 129978
rect 374058 112350 374678 129922
rect 374058 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 374678 112350
rect 374058 112226 374678 112294
rect 374058 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 374678 112226
rect 374058 112102 374678 112170
rect 374058 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 374678 112102
rect 374058 111978 374678 112046
rect 374058 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 374678 111978
rect 374058 98428 374678 111922
rect 377778 154350 378398 164250
rect 377778 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 378398 154350
rect 377778 154226 378398 154294
rect 377778 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 378398 154226
rect 377778 154102 378398 154170
rect 377778 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 378398 154102
rect 377778 153978 378398 154046
rect 377778 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 378398 153978
rect 377778 136350 378398 153922
rect 377778 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 378398 136350
rect 377778 136226 378398 136294
rect 377778 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 378398 136226
rect 377778 136102 378398 136170
rect 377778 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 378398 136102
rect 377778 135978 378398 136046
rect 377778 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 378398 135978
rect 377778 118350 378398 135922
rect 377778 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 378398 118350
rect 377778 118226 378398 118294
rect 377778 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 378398 118226
rect 377778 118102 378398 118170
rect 377778 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 378398 118102
rect 377778 117978 378398 118046
rect 377778 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 378398 117978
rect 377778 100350 378398 117922
rect 404778 148350 405398 164250
rect 404778 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 405398 148350
rect 404778 148226 405398 148294
rect 404778 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 405398 148226
rect 404778 148102 405398 148170
rect 404778 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 405398 148102
rect 404778 147978 405398 148046
rect 404778 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 405398 147978
rect 404778 130350 405398 147922
rect 404778 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 405398 130350
rect 404778 130226 405398 130294
rect 404778 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 405398 130226
rect 404778 130102 405398 130170
rect 404778 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 405398 130102
rect 404778 129978 405398 130046
rect 404778 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 405398 129978
rect 404778 112350 405398 129922
rect 404778 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 405398 112350
rect 404778 112226 405398 112294
rect 404778 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 405398 112226
rect 404778 112102 405398 112170
rect 404778 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 405398 112102
rect 404778 111978 405398 112046
rect 404778 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 405398 111978
rect 398188 110098 398244 110108
rect 396508 106678 396564 106688
rect 392364 104158 392420 104168
rect 389228 103978 389284 103988
rect 389228 103236 389284 103922
rect 392364 103348 392420 104102
rect 396508 104132 396564 106622
rect 396508 104066 396564 104076
rect 398188 104132 398244 110042
rect 398188 104066 398244 104076
rect 392364 103282 392420 103292
rect 389228 103170 389284 103180
rect 377778 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 378398 100350
rect 377778 100226 378398 100294
rect 377778 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 378398 100226
rect 377778 100102 378398 100170
rect 377778 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 378398 100102
rect 377778 99978 378398 100046
rect 377778 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 378398 99978
rect 356636 97234 356692 97244
rect 377778 96334 378398 99922
rect 404778 98428 405398 111922
rect 408498 154350 409118 164250
rect 422492 159572 422548 159582
rect 421596 156358 421652 156368
rect 421596 154532 421652 156302
rect 421596 154466 421652 154476
rect 408498 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 409118 154350
rect 408498 154226 409118 154294
rect 408498 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 409118 154226
rect 408498 154102 409118 154170
rect 408498 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 409118 154102
rect 408498 153978 409118 154046
rect 408498 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 409118 153978
rect 408498 136350 409118 153922
rect 421708 145738 421764 145748
rect 421708 144564 421764 145682
rect 422492 145558 422548 159516
rect 422492 144676 422548 145502
rect 422492 144610 422548 144620
rect 435498 148350 436118 164250
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 421708 144498 421764 144508
rect 408498 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 409118 136350
rect 408498 136226 409118 136294
rect 408498 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 409118 136226
rect 408498 136102 409118 136170
rect 408498 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 409118 136102
rect 408498 135978 409118 136046
rect 408498 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 409118 135978
rect 408498 118350 409118 135922
rect 435498 130350 436118 147922
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 423276 122724 423332 122734
rect 423276 122518 423332 122668
rect 423276 122452 423332 122462
rect 408498 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 409118 118350
rect 408498 118226 409118 118294
rect 408498 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 409118 118226
rect 408498 118102 409118 118170
rect 408498 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 409118 118102
rect 408498 117978 409118 118046
rect 408498 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 409118 117978
rect 408498 100350 409118 117922
rect 408498 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 409118 100350
rect 408498 100226 409118 100294
rect 408498 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 409118 100226
rect 408498 100102 409118 100170
rect 408498 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 409118 100102
rect 408498 99978 409118 100046
rect 408498 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 409118 99978
rect 408498 96334 409118 99922
rect 435498 112350 436118 129922
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 419356 99092 419412 99102
rect 419356 97076 419412 99036
rect 419356 97010 419412 97020
rect 421708 98196 421764 98206
rect 374448 94350 374768 94384
rect 374448 94294 374518 94350
rect 374574 94294 374642 94350
rect 374698 94294 374768 94350
rect 374448 94226 374768 94294
rect 374448 94170 374518 94226
rect 374574 94170 374642 94226
rect 374698 94170 374768 94226
rect 374448 94102 374768 94170
rect 374448 94046 374518 94102
rect 374574 94046 374642 94102
rect 374698 94046 374768 94102
rect 374448 93978 374768 94046
rect 374448 93922 374518 93978
rect 374574 93922 374642 93978
rect 374698 93922 374768 93978
rect 374448 93888 374768 93922
rect 405168 94350 405488 94384
rect 405168 94294 405238 94350
rect 405294 94294 405362 94350
rect 405418 94294 405488 94350
rect 405168 94226 405488 94294
rect 405168 94170 405238 94226
rect 405294 94170 405362 94226
rect 405418 94170 405488 94226
rect 405168 94102 405488 94170
rect 405168 94046 405238 94102
rect 405294 94046 405362 94102
rect 405418 94046 405488 94102
rect 405168 93978 405488 94046
rect 405168 93922 405238 93978
rect 405294 93922 405362 93978
rect 405418 93922 405488 93978
rect 405168 93888 405488 93922
rect 351932 91522 351988 91532
rect 421708 91588 421764 98140
rect 425852 96628 425908 96638
rect 421708 91522 421764 91532
rect 424172 91588 424228 91598
rect 347058 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 347678 82350
rect 347058 82226 347678 82294
rect 347058 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 347678 82226
rect 347058 82102 347678 82170
rect 347058 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 347678 82102
rect 347058 81978 347678 82046
rect 347058 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 347678 81978
rect 347058 64350 347678 81922
rect 389808 82350 390128 82384
rect 389808 82294 389878 82350
rect 389934 82294 390002 82350
rect 390058 82294 390128 82350
rect 389808 82226 390128 82294
rect 389808 82170 389878 82226
rect 389934 82170 390002 82226
rect 390058 82170 390128 82226
rect 389808 82102 390128 82170
rect 389808 82046 389878 82102
rect 389934 82046 390002 82102
rect 390058 82046 390128 82102
rect 389808 81978 390128 82046
rect 389808 81922 389878 81978
rect 389934 81922 390002 81978
rect 390058 81922 390128 81978
rect 389808 81888 390128 81922
rect 374448 76350 374768 76384
rect 374448 76294 374518 76350
rect 374574 76294 374642 76350
rect 374698 76294 374768 76350
rect 374448 76226 374768 76294
rect 374448 76170 374518 76226
rect 374574 76170 374642 76226
rect 374698 76170 374768 76226
rect 374448 76102 374768 76170
rect 374448 76046 374518 76102
rect 374574 76046 374642 76102
rect 374698 76046 374768 76102
rect 374448 75978 374768 76046
rect 374448 75922 374518 75978
rect 374574 75922 374642 75978
rect 374698 75922 374768 75978
rect 374448 75888 374768 75922
rect 405168 76350 405488 76384
rect 405168 76294 405238 76350
rect 405294 76294 405362 76350
rect 405418 76294 405488 76350
rect 405168 76226 405488 76294
rect 405168 76170 405238 76226
rect 405294 76170 405362 76226
rect 405418 76170 405488 76226
rect 405168 76102 405488 76170
rect 405168 76046 405238 76102
rect 405294 76046 405362 76102
rect 405418 76046 405488 76102
rect 405168 75978 405488 76046
rect 405168 75922 405238 75978
rect 405294 75922 405362 75978
rect 405418 75922 405488 75978
rect 405168 75888 405488 75922
rect 347058 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 347678 64350
rect 347058 64226 347678 64294
rect 347058 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 347678 64226
rect 347058 64102 347678 64170
rect 347058 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 347678 64102
rect 347058 63978 347678 64046
rect 347058 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 347678 63978
rect 343338 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 343958 40350
rect 343338 40226 343958 40294
rect 343338 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 343958 40226
rect 343338 40102 343958 40170
rect 343338 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 343958 40102
rect 343338 39978 343958 40046
rect 343338 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 343958 39978
rect 316338 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 316958 28350
rect 316338 28226 316958 28294
rect 316338 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 316958 28226
rect 316338 28102 316958 28170
rect 316338 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 316958 28102
rect 316338 27978 316958 28046
rect 316338 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 316958 27978
rect 316338 10350 316958 27922
rect 316338 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 316958 10350
rect 316338 10226 316958 10294
rect 316338 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 316958 10226
rect 316338 10102 316958 10170
rect 316338 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 316958 10102
rect 316338 9978 316958 10046
rect 316338 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 316958 9978
rect 316338 -1120 316958 9922
rect 316338 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 316958 -1120
rect 316338 -1244 316958 -1176
rect 316338 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 316958 -1244
rect 316338 -1368 316958 -1300
rect 316338 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 316958 -1368
rect 316338 -1492 316958 -1424
rect 316338 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 316958 -1492
rect 316338 -1644 316958 -1548
rect 343338 22350 343958 39922
rect 343338 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 343958 22350
rect 343338 22226 343958 22294
rect 343338 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 343958 22226
rect 343338 22102 343958 22170
rect 343338 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 343958 22102
rect 343338 21978 343958 22046
rect 343338 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 343958 21978
rect 343338 4350 343958 21922
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 347058 46350 347678 63922
rect 389808 64350 390128 64384
rect 389808 64294 389878 64350
rect 389934 64294 390002 64350
rect 390058 64294 390128 64350
rect 389808 64226 390128 64294
rect 389808 64170 389878 64226
rect 389934 64170 390002 64226
rect 390058 64170 390128 64226
rect 389808 64102 390128 64170
rect 389808 64046 389878 64102
rect 389934 64046 390002 64102
rect 390058 64046 390128 64102
rect 389808 63978 390128 64046
rect 389808 63922 389878 63978
rect 389934 63922 390002 63978
rect 390058 63922 390128 63978
rect 389808 63888 390128 63922
rect 424172 61348 424228 91532
rect 425852 66388 425908 96572
rect 425852 66322 425908 66332
rect 435498 94350 436118 111922
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 435498 76350 436118 93922
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 424172 61282 424228 61292
rect 374448 58350 374768 58384
rect 374448 58294 374518 58350
rect 374574 58294 374642 58350
rect 374698 58294 374768 58350
rect 374448 58226 374768 58294
rect 374448 58170 374518 58226
rect 374574 58170 374642 58226
rect 374698 58170 374768 58226
rect 374448 58102 374768 58170
rect 374448 58046 374518 58102
rect 374574 58046 374642 58102
rect 374698 58046 374768 58102
rect 374448 57978 374768 58046
rect 374448 57922 374518 57978
rect 374574 57922 374642 57978
rect 374698 57922 374768 57978
rect 374448 57888 374768 57922
rect 405168 58350 405488 58384
rect 405168 58294 405238 58350
rect 405294 58294 405362 58350
rect 405418 58294 405488 58350
rect 405168 58226 405488 58294
rect 405168 58170 405238 58226
rect 405294 58170 405362 58226
rect 405418 58170 405488 58226
rect 405168 58102 405488 58170
rect 405168 58046 405238 58102
rect 405294 58046 405362 58102
rect 405418 58046 405488 58102
rect 405168 57978 405488 58046
rect 405168 57922 405238 57978
rect 405294 57922 405362 57978
rect 405418 57922 405488 57978
rect 405168 57888 405488 57922
rect 435498 58350 436118 75922
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 347058 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 347678 46350
rect 347058 46226 347678 46294
rect 347058 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 347678 46226
rect 347058 46102 347678 46170
rect 347058 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 347678 46102
rect 347058 45978 347678 46046
rect 347058 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 347678 45978
rect 347058 28350 347678 45922
rect 347058 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 347678 28350
rect 347058 28226 347678 28294
rect 347058 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 347678 28226
rect 347058 28102 347678 28170
rect 347058 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 347678 28102
rect 347058 27978 347678 28046
rect 347058 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 347678 27978
rect 347058 10350 347678 27922
rect 347058 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 347678 10350
rect 347058 10226 347678 10294
rect 347058 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 347678 10226
rect 347058 10102 347678 10170
rect 347058 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 347678 10102
rect 347058 9978 347678 10046
rect 347058 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 347678 9978
rect 347058 -1120 347678 9922
rect 347058 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 347678 -1120
rect 347058 -1244 347678 -1176
rect 347058 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 347678 -1244
rect 347058 -1368 347678 -1300
rect 347058 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 347678 -1368
rect 347058 -1492 347678 -1424
rect 347058 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 347678 -1492
rect 347058 -1644 347678 -1548
rect 374058 40350 374678 49026
rect 374058 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 374678 40350
rect 374058 40226 374678 40294
rect 374058 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 374678 40226
rect 374058 40102 374678 40170
rect 374058 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 374678 40102
rect 374058 39978 374678 40046
rect 374058 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 374678 39978
rect 374058 22350 374678 39922
rect 374058 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 374678 22350
rect 374058 22226 374678 22294
rect 374058 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 374678 22226
rect 374058 22102 374678 22170
rect 374058 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 374678 22102
rect 374058 21978 374678 22046
rect 374058 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 374678 21978
rect 374058 4350 374678 21922
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 377778 46350 378398 49026
rect 377778 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 378398 46350
rect 377778 46226 378398 46294
rect 377778 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 378398 46226
rect 377778 46102 378398 46170
rect 377778 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 378398 46102
rect 377778 45978 378398 46046
rect 377778 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 378398 45978
rect 377778 28350 378398 45922
rect 377778 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 378398 28350
rect 377778 28226 378398 28294
rect 377778 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 378398 28226
rect 377778 28102 378398 28170
rect 377778 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 378398 28102
rect 377778 27978 378398 28046
rect 377778 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 378398 27978
rect 377778 10350 378398 27922
rect 377778 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 378398 10350
rect 377778 10226 378398 10294
rect 377778 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 378398 10226
rect 377778 10102 378398 10170
rect 377778 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 378398 10102
rect 377778 9978 378398 10046
rect 377778 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 378398 9978
rect 377778 -1120 378398 9922
rect 377778 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 378398 -1120
rect 377778 -1244 378398 -1176
rect 377778 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 378398 -1244
rect 377778 -1368 378398 -1300
rect 377778 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 378398 -1368
rect 377778 -1492 378398 -1424
rect 377778 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 378398 -1492
rect 377778 -1644 378398 -1548
rect 404778 40350 405398 49026
rect 404778 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 405398 40350
rect 404778 40226 405398 40294
rect 404778 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 405398 40226
rect 404778 40102 405398 40170
rect 404778 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 405398 40102
rect 404778 39978 405398 40046
rect 404778 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 405398 39978
rect 404778 22350 405398 39922
rect 404778 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 405398 22350
rect 404778 22226 405398 22294
rect 404778 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 405398 22226
rect 404778 22102 405398 22170
rect 404778 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 405398 22102
rect 404778 21978 405398 22046
rect 404778 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 405398 21978
rect 404778 4350 405398 21922
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 408498 46350 409118 49026
rect 408498 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 409118 46350
rect 408498 46226 409118 46294
rect 408498 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 409118 46226
rect 408498 46102 409118 46170
rect 408498 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 409118 46102
rect 408498 45978 409118 46046
rect 408498 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 409118 45978
rect 408498 28350 409118 45922
rect 408498 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 409118 28350
rect 408498 28226 409118 28294
rect 408498 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 409118 28226
rect 408498 28102 409118 28170
rect 408498 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 409118 28102
rect 408498 27978 409118 28046
rect 408498 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 409118 27978
rect 408498 10350 409118 27922
rect 408498 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 409118 10350
rect 408498 10226 409118 10294
rect 408498 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 409118 10226
rect 408498 10102 409118 10170
rect 408498 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 409118 10102
rect 408498 9978 409118 10046
rect 408498 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 409118 9978
rect 408498 -1120 409118 9922
rect 408498 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 409118 -1120
rect 408498 -1244 409118 -1176
rect 408498 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 409118 -1244
rect 408498 -1368 409118 -1300
rect 408498 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 409118 -1368
rect 408498 -1492 409118 -1424
rect 408498 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 409118 -1492
rect 408498 -1644 409118 -1548
rect 435498 40350 436118 57922
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 435498 4350 436118 21922
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 435498 4102 436118 4170
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 154350 439838 164250
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 457772 163044 457828 163054
rect 457212 151318 457268 151328
rect 456988 150058 457044 150068
rect 456988 147812 457044 150002
rect 456988 147746 457044 147756
rect 457212 142772 457268 151262
rect 457660 147924 457716 147934
rect 457660 147364 457716 147868
rect 457660 147298 457716 147308
rect 457212 142706 457268 142716
rect 457772 140980 457828 162988
rect 457884 149380 457940 164780
rect 487788 164098 487844 164108
rect 462812 163268 462868 163278
rect 460012 163156 460068 163166
rect 460012 156100 460068 163100
rect 460124 161588 460180 161598
rect 460124 156178 460180 161532
rect 460236 161476 460292 161486
rect 460236 157438 460292 161420
rect 460236 157372 460292 157382
rect 460460 158116 460516 158126
rect 460124 156112 460180 156122
rect 460012 156034 460068 156044
rect 460348 154918 460404 154928
rect 457884 149314 457940 149324
rect 458444 154738 458500 154748
rect 458444 147476 458500 154682
rect 458444 147410 458500 147420
rect 460348 144478 460404 154862
rect 460460 145918 460516 158060
rect 461244 156538 461300 156548
rect 460460 145852 460516 145862
rect 460572 156324 460628 156334
rect 460348 144412 460404 144422
rect 460572 144298 460628 156268
rect 460572 144232 460628 144242
rect 460684 154756 460740 154766
rect 457772 140914 457828 140924
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 439218 118350 439838 135922
rect 460684 122518 460740 154700
rect 461132 149878 461188 149888
rect 461132 140878 461188 149822
rect 461244 147718 461300 156482
rect 461244 147652 461300 147662
rect 461580 151396 461636 151406
rect 461580 145558 461636 151340
rect 461916 150500 461972 150510
rect 461692 149716 461748 149726
rect 461692 145738 461748 149660
rect 461916 148820 461972 150444
rect 461916 148754 461972 148764
rect 461692 145672 461748 145682
rect 461580 145492 461636 145502
rect 462812 141058 462868 163212
rect 477036 162932 477092 162942
rect 462924 161700 462980 161710
rect 462924 142678 462980 161644
rect 468636 157892 468692 157902
rect 468636 154532 468692 157836
rect 477036 157618 477092 162876
rect 483756 162478 483812 162488
rect 480396 160858 480452 160868
rect 480396 159796 480452 160802
rect 480396 159730 480452 159740
rect 477036 157552 477092 157562
rect 468636 154466 468692 154476
rect 475692 154918 475748 154928
rect 463708 153188 463764 153198
rect 463708 152578 463764 153132
rect 475692 152964 475748 154862
rect 483756 154532 483812 162422
rect 483756 154466 483812 154476
rect 485100 155638 485156 155648
rect 475692 152898 475748 152908
rect 485100 152964 485156 155582
rect 487788 154532 487844 164042
rect 487788 154466 487844 154476
rect 488908 154532 488964 165482
rect 557900 164836 557956 164846
rect 488908 154466 488964 154476
rect 489244 164818 489300 164828
rect 489244 154532 489300 164762
rect 493164 163918 493220 163928
rect 489244 154466 489300 154476
rect 491820 162298 491876 162308
rect 491820 154532 491876 162242
rect 491820 154466 491876 154476
rect 493164 154532 493220 163862
rect 553644 163828 553700 163838
rect 497868 162932 497924 162942
rect 497868 157798 497924 162876
rect 532364 162932 532420 162942
rect 532364 159598 532420 162876
rect 539308 162932 539364 162942
rect 539308 162838 539364 162876
rect 539308 162772 539364 162782
rect 546476 162932 546532 162942
rect 546476 161218 546532 162876
rect 546476 161152 546532 161162
rect 532364 159532 532420 159542
rect 497868 157732 497924 157742
rect 493164 154466 493220 154476
rect 494508 156538 494564 156548
rect 485100 152898 485156 152908
rect 494508 152964 494564 156482
rect 494508 152898 494564 152908
rect 497308 154308 497364 154318
rect 497308 152938 497364 154252
rect 499884 153658 499940 153668
rect 498540 153478 498596 153488
rect 498540 152964 498596 153422
rect 498540 152898 498596 152908
rect 499884 152964 499940 153602
rect 499884 152898 499940 152908
rect 497308 152872 497364 152882
rect 463708 152512 463764 152522
rect 463596 151284 463652 151294
rect 462924 142612 462980 142622
rect 463036 149828 463092 149838
rect 462812 140992 462868 141002
rect 461132 140812 461188 140822
rect 463036 139438 463092 149772
rect 463596 146098 463652 151228
rect 477036 149940 477092 149950
rect 477036 149878 477092 149884
rect 477036 149812 477092 149822
rect 494732 149716 494788 149726
rect 494508 149380 494564 149390
rect 494508 149156 494564 149324
rect 494508 149090 494564 149100
rect 494732 149156 494788 149660
rect 500108 149716 500164 149726
rect 500108 149380 500164 149660
rect 500108 149314 500164 149324
rect 494732 149090 494788 149100
rect 463596 146032 463652 146042
rect 463036 139372 463092 139382
rect 479808 136350 480128 136384
rect 479808 136294 479878 136350
rect 479934 136294 480002 136350
rect 480058 136294 480128 136350
rect 479808 136226 480128 136294
rect 479808 136170 479878 136226
rect 479934 136170 480002 136226
rect 480058 136170 480128 136226
rect 479808 136102 480128 136170
rect 479808 136046 479878 136102
rect 479934 136046 480002 136102
rect 480058 136046 480128 136102
rect 479808 135978 480128 136046
rect 479808 135922 479878 135978
rect 479934 135922 480002 135978
rect 480058 135922 480128 135978
rect 479808 135888 480128 135922
rect 510528 136350 510848 136384
rect 510528 136294 510598 136350
rect 510654 136294 510722 136350
rect 510778 136294 510848 136350
rect 510528 136226 510848 136294
rect 510528 136170 510598 136226
rect 510654 136170 510722 136226
rect 510778 136170 510848 136226
rect 510528 136102 510848 136170
rect 510528 136046 510598 136102
rect 510654 136046 510722 136102
rect 510778 136046 510848 136102
rect 510528 135978 510848 136046
rect 510528 135922 510598 135978
rect 510654 135922 510722 135978
rect 510778 135922 510848 135978
rect 510528 135888 510848 135922
rect 541248 136350 541568 136384
rect 541248 136294 541318 136350
rect 541374 136294 541442 136350
rect 541498 136294 541568 136350
rect 541248 136226 541568 136294
rect 541248 136170 541318 136226
rect 541374 136170 541442 136226
rect 541498 136170 541568 136226
rect 541248 136102 541568 136170
rect 541248 136046 541318 136102
rect 541374 136046 541442 136102
rect 541498 136046 541568 136102
rect 541248 135978 541568 136046
rect 541248 135922 541318 135978
rect 541374 135922 541442 135978
rect 541498 135922 541568 135978
rect 541248 135888 541568 135922
rect 464448 130350 464768 130384
rect 464448 130294 464518 130350
rect 464574 130294 464642 130350
rect 464698 130294 464768 130350
rect 464448 130226 464768 130294
rect 464448 130170 464518 130226
rect 464574 130170 464642 130226
rect 464698 130170 464768 130226
rect 464448 130102 464768 130170
rect 464448 130046 464518 130102
rect 464574 130046 464642 130102
rect 464698 130046 464768 130102
rect 464448 129978 464768 130046
rect 464448 129922 464518 129978
rect 464574 129922 464642 129978
rect 464698 129922 464768 129978
rect 464448 129888 464768 129922
rect 495168 130350 495488 130384
rect 495168 130294 495238 130350
rect 495294 130294 495362 130350
rect 495418 130294 495488 130350
rect 495168 130226 495488 130294
rect 495168 130170 495238 130226
rect 495294 130170 495362 130226
rect 495418 130170 495488 130226
rect 495168 130102 495488 130170
rect 495168 130046 495238 130102
rect 495294 130046 495362 130102
rect 495418 130046 495488 130102
rect 495168 129978 495488 130046
rect 495168 129922 495238 129978
rect 495294 129922 495362 129978
rect 495418 129922 495488 129978
rect 495168 129888 495488 129922
rect 525888 130350 526208 130384
rect 525888 130294 525958 130350
rect 526014 130294 526082 130350
rect 526138 130294 526208 130350
rect 525888 130226 526208 130294
rect 525888 130170 525958 130226
rect 526014 130170 526082 130226
rect 526138 130170 526208 130226
rect 525888 130102 526208 130170
rect 525888 130046 525958 130102
rect 526014 130046 526082 130102
rect 526138 130046 526208 130102
rect 525888 129978 526208 130046
rect 525888 129922 525958 129978
rect 526014 129922 526082 129978
rect 526138 129922 526208 129978
rect 525888 129888 526208 129922
rect 460684 122452 460740 122462
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 439218 100350 439838 117922
rect 479808 118350 480128 118384
rect 479808 118294 479878 118350
rect 479934 118294 480002 118350
rect 480058 118294 480128 118350
rect 479808 118226 480128 118294
rect 479808 118170 479878 118226
rect 479934 118170 480002 118226
rect 480058 118170 480128 118226
rect 479808 118102 480128 118170
rect 479808 118046 479878 118102
rect 479934 118046 480002 118102
rect 480058 118046 480128 118102
rect 479808 117978 480128 118046
rect 479808 117922 479878 117978
rect 479934 117922 480002 117978
rect 480058 117922 480128 117978
rect 479808 117888 480128 117922
rect 510528 118350 510848 118384
rect 510528 118294 510598 118350
rect 510654 118294 510722 118350
rect 510778 118294 510848 118350
rect 510528 118226 510848 118294
rect 510528 118170 510598 118226
rect 510654 118170 510722 118226
rect 510778 118170 510848 118226
rect 510528 118102 510848 118170
rect 510528 118046 510598 118102
rect 510654 118046 510722 118102
rect 510778 118046 510848 118102
rect 510528 117978 510848 118046
rect 510528 117922 510598 117978
rect 510654 117922 510722 117978
rect 510778 117922 510848 117978
rect 510528 117888 510848 117922
rect 541248 118350 541568 118384
rect 541248 118294 541318 118350
rect 541374 118294 541442 118350
rect 541498 118294 541568 118350
rect 541248 118226 541568 118294
rect 541248 118170 541318 118226
rect 541374 118170 541442 118226
rect 541498 118170 541568 118226
rect 541248 118102 541568 118170
rect 541248 118046 541318 118102
rect 541374 118046 541442 118102
rect 541498 118046 541568 118102
rect 541248 117978 541568 118046
rect 541248 117922 541318 117978
rect 541374 117922 541442 117978
rect 541498 117922 541568 117978
rect 541248 117888 541568 117922
rect 553644 116938 553700 163772
rect 554316 163738 554372 163748
rect 553980 163156 554036 163166
rect 553868 157978 553924 157988
rect 553644 116872 553700 116882
rect 553756 150058 553812 150068
rect 464448 112350 464768 112384
rect 464448 112294 464518 112350
rect 464574 112294 464642 112350
rect 464698 112294 464768 112350
rect 464448 112226 464768 112294
rect 464448 112170 464518 112226
rect 464574 112170 464642 112226
rect 464698 112170 464768 112226
rect 464448 112102 464768 112170
rect 464448 112046 464518 112102
rect 464574 112046 464642 112102
rect 464698 112046 464768 112102
rect 464448 111978 464768 112046
rect 464448 111922 464518 111978
rect 464574 111922 464642 111978
rect 464698 111922 464768 111978
rect 464448 111888 464768 111922
rect 495168 112350 495488 112384
rect 495168 112294 495238 112350
rect 495294 112294 495362 112350
rect 495418 112294 495488 112350
rect 495168 112226 495488 112294
rect 495168 112170 495238 112226
rect 495294 112170 495362 112226
rect 495418 112170 495488 112226
rect 495168 112102 495488 112170
rect 495168 112046 495238 112102
rect 495294 112046 495362 112102
rect 495418 112046 495488 112102
rect 495168 111978 495488 112046
rect 495168 111922 495238 111978
rect 495294 111922 495362 111978
rect 495418 111922 495488 111978
rect 495168 111888 495488 111922
rect 525888 112350 526208 112384
rect 525888 112294 525958 112350
rect 526014 112294 526082 112350
rect 526138 112294 526208 112350
rect 525888 112226 526208 112294
rect 525888 112170 525958 112226
rect 526014 112170 526082 112226
rect 526138 112170 526208 112226
rect 525888 112102 526208 112170
rect 525888 112046 525958 112102
rect 526014 112046 526082 112102
rect 526138 112046 526208 112102
rect 525888 111978 526208 112046
rect 525888 111922 525958 111978
rect 526014 111922 526082 111978
rect 526138 111922 526208 111978
rect 525888 111888 526208 111922
rect 458108 110068 458164 110078
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 439218 82350 439838 99922
rect 457884 101668 457940 101678
rect 457436 98868 457492 98878
rect 457324 98308 457380 98318
rect 457324 89796 457380 98252
rect 457324 89730 457380 89740
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 439218 64350 439838 81922
rect 457436 81060 457492 98812
rect 457772 98532 457828 98542
rect 457660 98420 457716 98430
rect 457660 98218 457716 98364
rect 457660 98152 457716 98162
rect 457548 97300 457604 97310
rect 457548 94798 457604 97244
rect 457660 95508 457716 95518
rect 457660 94978 457716 95452
rect 457660 94912 457716 94922
rect 457548 94742 457716 94798
rect 457660 86884 457716 94742
rect 457660 86818 457716 86828
rect 457436 80994 457492 81004
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 439218 46350 439838 63922
rect 457548 66388 457604 66398
rect 457548 60676 457604 66332
rect 457772 63588 457828 98476
rect 457884 69412 457940 101612
rect 457884 69346 457940 69356
rect 457996 98980 458052 98990
rect 457996 66500 458052 98924
rect 458108 83972 458164 110012
rect 553756 109228 553812 150002
rect 553420 109172 553812 109228
rect 553420 105868 553476 109172
rect 553868 105868 553924 157922
rect 553196 105812 553476 105868
rect 553756 105812 553924 105868
rect 458108 83906 458164 83916
rect 458220 105140 458276 105150
rect 458220 78148 458276 105084
rect 479808 100350 480128 100384
rect 479808 100294 479878 100350
rect 479934 100294 480002 100350
rect 480058 100294 480128 100350
rect 479808 100226 480128 100294
rect 479808 100170 479878 100226
rect 479934 100170 480002 100226
rect 480058 100170 480128 100226
rect 479808 100102 480128 100170
rect 479808 100046 479878 100102
rect 479934 100046 480002 100102
rect 480058 100046 480128 100102
rect 479808 99978 480128 100046
rect 479808 99922 479878 99978
rect 479934 99922 480002 99978
rect 480058 99922 480128 99978
rect 479808 99888 480128 99922
rect 510528 100350 510848 100384
rect 510528 100294 510598 100350
rect 510654 100294 510722 100350
rect 510778 100294 510848 100350
rect 510528 100226 510848 100294
rect 510528 100170 510598 100226
rect 510654 100170 510722 100226
rect 510778 100170 510848 100226
rect 510528 100102 510848 100170
rect 510528 100046 510598 100102
rect 510654 100046 510722 100102
rect 510778 100046 510848 100102
rect 510528 99978 510848 100046
rect 510528 99922 510598 99978
rect 510654 99922 510722 99978
rect 510778 99922 510848 99978
rect 510528 99888 510848 99922
rect 541248 100350 541568 100384
rect 541248 100294 541318 100350
rect 541374 100294 541442 100350
rect 541498 100294 541568 100350
rect 541248 100226 541568 100294
rect 541248 100170 541318 100226
rect 541374 100170 541442 100226
rect 541498 100170 541568 100226
rect 541248 100102 541568 100170
rect 541248 100046 541318 100102
rect 541374 100046 541442 100102
rect 541498 100046 541568 100102
rect 541248 99978 541568 100046
rect 541248 99922 541318 99978
rect 541374 99922 541442 99978
rect 541498 99922 541568 99978
rect 541248 99888 541568 99922
rect 553196 99658 553252 105812
rect 553196 99592 553252 99602
rect 553308 105418 553364 105428
rect 458220 78082 458276 78092
rect 458332 98644 458388 98654
rect 458332 75236 458388 98588
rect 464448 94350 464768 94384
rect 464448 94294 464518 94350
rect 464574 94294 464642 94350
rect 464698 94294 464768 94350
rect 464448 94226 464768 94294
rect 464448 94170 464518 94226
rect 464574 94170 464642 94226
rect 464698 94170 464768 94226
rect 464448 94102 464768 94170
rect 464448 94046 464518 94102
rect 464574 94046 464642 94102
rect 464698 94046 464768 94102
rect 464448 93978 464768 94046
rect 464448 93922 464518 93978
rect 464574 93922 464642 93978
rect 464698 93922 464768 93978
rect 464448 93888 464768 93922
rect 495168 94350 495488 94384
rect 495168 94294 495238 94350
rect 495294 94294 495362 94350
rect 495418 94294 495488 94350
rect 495168 94226 495488 94294
rect 495168 94170 495238 94226
rect 495294 94170 495362 94226
rect 495418 94170 495488 94226
rect 495168 94102 495488 94170
rect 495168 94046 495238 94102
rect 495294 94046 495362 94102
rect 495418 94046 495488 94102
rect 495168 93978 495488 94046
rect 495168 93922 495238 93978
rect 495294 93922 495362 93978
rect 495418 93922 495488 93978
rect 495168 93888 495488 93922
rect 525888 94350 526208 94384
rect 525888 94294 525958 94350
rect 526014 94294 526082 94350
rect 526138 94294 526208 94350
rect 525888 94226 526208 94294
rect 525888 94170 525958 94226
rect 526014 94170 526082 94226
rect 526138 94170 526208 94226
rect 525888 94102 526208 94170
rect 525888 94046 525958 94102
rect 526014 94046 526082 94102
rect 526138 94046 526208 94102
rect 553308 94108 553364 105362
rect 553756 103978 553812 105812
rect 553980 105364 554036 163100
rect 553756 103912 553812 103922
rect 553868 105308 554036 105364
rect 554092 148820 554148 148830
rect 554092 105418 554148 148764
rect 554316 114268 554372 163682
rect 556220 163044 556276 163054
rect 554652 161588 554708 161598
rect 554540 158878 554596 158888
rect 554204 114212 554372 114268
rect 554428 156358 554484 156368
rect 554204 109198 554260 114212
rect 554204 109142 554372 109198
rect 554092 105352 554148 105362
rect 553868 100660 553924 105308
rect 554316 104132 554372 109142
rect 554316 104066 554372 104076
rect 554316 103978 554372 103988
rect 554316 102228 554372 103922
rect 554316 102162 554372 102172
rect 554316 100660 554372 100670
rect 553868 100604 554316 100660
rect 554316 100594 554372 100604
rect 554316 99988 554372 99998
rect 554316 99838 554372 99932
rect 554204 99782 554372 99838
rect 553308 94052 553588 94108
rect 525888 93978 526208 94046
rect 525888 93922 525958 93978
rect 526014 93922 526082 93978
rect 526138 93922 526208 93978
rect 525888 93888 526208 93922
rect 553532 90748 553588 94052
rect 553532 90692 554148 90748
rect 479808 82350 480128 82384
rect 479808 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 480128 82350
rect 479808 82226 480128 82294
rect 479808 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 480128 82226
rect 479808 82102 480128 82170
rect 479808 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 480128 82102
rect 479808 81978 480128 82046
rect 479808 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 480128 81978
rect 479808 81888 480128 81922
rect 510528 82350 510848 82384
rect 510528 82294 510598 82350
rect 510654 82294 510722 82350
rect 510778 82294 510848 82350
rect 510528 82226 510848 82294
rect 510528 82170 510598 82226
rect 510654 82170 510722 82226
rect 510778 82170 510848 82226
rect 510528 82102 510848 82170
rect 510528 82046 510598 82102
rect 510654 82046 510722 82102
rect 510778 82046 510848 82102
rect 510528 81978 510848 82046
rect 510528 81922 510598 81978
rect 510654 81922 510722 81978
rect 510778 81922 510848 81978
rect 510528 81888 510848 81922
rect 541248 82350 541568 82384
rect 541248 82294 541318 82350
rect 541374 82294 541442 82350
rect 541498 82294 541568 82350
rect 554092 82348 554148 90692
rect 541248 82226 541568 82294
rect 541248 82170 541318 82226
rect 541374 82170 541442 82226
rect 541498 82170 541568 82226
rect 541248 82102 541568 82170
rect 541248 82046 541318 82102
rect 541374 82046 541442 82102
rect 541498 82046 541568 82102
rect 541248 81978 541568 82046
rect 541248 81922 541318 81978
rect 541374 81922 541442 81978
rect 541498 81922 541568 81978
rect 541248 81888 541568 81922
rect 553980 82292 554148 82348
rect 554204 82348 554260 99782
rect 554316 99658 554372 99668
rect 554316 94388 554372 99602
rect 554316 94322 554372 94332
rect 554316 82348 554372 82358
rect 554204 82292 554316 82348
rect 464448 76350 464768 76384
rect 464448 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 464768 76350
rect 464448 76226 464768 76294
rect 464448 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 464768 76226
rect 464448 76102 464768 76170
rect 464448 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 464768 76102
rect 464448 75978 464768 76046
rect 464448 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 464768 75978
rect 464448 75888 464768 75922
rect 495168 76350 495488 76384
rect 495168 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 495488 76350
rect 495168 76226 495488 76294
rect 495168 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 495488 76226
rect 495168 76102 495488 76170
rect 495168 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 495488 76102
rect 495168 75978 495488 76046
rect 495168 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 495488 75978
rect 495168 75888 495488 75922
rect 525888 76350 526208 76384
rect 525888 76294 525958 76350
rect 526014 76294 526082 76350
rect 526138 76294 526208 76350
rect 525888 76226 526208 76294
rect 525888 76170 525958 76226
rect 526014 76170 526082 76226
rect 526138 76170 526208 76226
rect 525888 76102 526208 76170
rect 525888 76046 525958 76102
rect 526014 76046 526082 76102
rect 526138 76046 526208 76102
rect 525888 75978 526208 76046
rect 525888 75922 525958 75978
rect 526014 75922 526082 75978
rect 526138 75922 526208 75978
rect 525888 75888 526208 75922
rect 458332 75170 458388 75180
rect 553980 74004 554036 82292
rect 554316 82282 554372 82292
rect 554316 74004 554372 74014
rect 553980 73948 554316 74004
rect 554316 73938 554372 73948
rect 554428 72436 554484 156302
rect 554540 80276 554596 158822
rect 554652 89684 554708 161532
rect 554764 160678 554820 160688
rect 554764 91252 554820 160622
rect 555212 160498 555268 160508
rect 555100 154738 555156 154748
rect 554988 150598 555044 150608
rect 554764 91186 554820 91196
rect 554876 149698 554932 149708
rect 554652 89618 554708 89628
rect 554540 80210 554596 80220
rect 554652 82292 554708 82302
rect 554428 72370 554484 72380
rect 554652 70588 554708 82236
rect 554876 81844 554932 149642
rect 554988 85316 555044 150542
rect 555100 92820 555156 154682
rect 555212 122612 555268 160442
rect 555212 122546 555268 122556
rect 556108 152938 556164 152948
rect 555212 116938 555268 116948
rect 555212 116834 555268 116844
rect 555100 92754 555156 92764
rect 554988 85250 555044 85260
rect 554876 81778 554932 81788
rect 556108 77140 556164 152882
rect 556220 95956 556276 162988
rect 556332 158698 556388 158708
rect 556332 117908 556388 158642
rect 557788 155458 557844 155468
rect 557788 151172 557844 155402
rect 557900 152852 557956 164780
rect 557900 152786 557956 152796
rect 558012 153188 558068 153198
rect 557788 151106 557844 151116
rect 557900 150418 557956 150428
rect 557788 148618 557844 148628
rect 557788 143892 557844 148562
rect 557788 143826 557844 143836
rect 557900 143758 557956 150362
rect 557788 143702 557956 143758
rect 557788 143444 557844 143702
rect 557788 143378 557844 143388
rect 557900 143556 557956 143566
rect 556332 117842 556388 117852
rect 557900 99092 557956 143500
rect 558012 103796 558068 153132
rect 558236 152218 558292 152228
rect 558124 152038 558180 152048
rect 558124 143668 558180 151982
rect 558236 147924 558292 152162
rect 558236 147858 558292 147868
rect 558378 148350 558998 164250
rect 558378 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 558998 148350
rect 558378 148226 558998 148294
rect 558378 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 558998 148226
rect 558378 148102 558998 148170
rect 558378 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 558998 148102
rect 558378 147978 558998 148046
rect 558378 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 558998 147978
rect 558124 143602 558180 143612
rect 558236 143892 558292 143902
rect 558124 143444 558180 143454
rect 558124 105364 558180 143388
rect 558236 106932 558292 143836
rect 558236 106866 558292 106876
rect 558378 130350 558998 147922
rect 558378 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 558998 130350
rect 558378 130226 558998 130294
rect 558378 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 558998 130226
rect 558378 130102 558998 130170
rect 558378 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 558998 130102
rect 558378 129978 558998 130046
rect 558378 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 558998 129978
rect 558378 112350 558998 129922
rect 558378 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 558998 112350
rect 558378 112226 558998 112294
rect 558378 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 558998 112226
rect 558378 112102 558998 112170
rect 558378 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 558998 112102
rect 558378 111978 558998 112046
rect 558378 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 558998 111978
rect 558124 105298 558180 105308
rect 558012 103730 558068 103740
rect 557900 99026 557956 99036
rect 556220 95890 556276 95900
rect 556108 77074 556164 77084
rect 558378 94350 558998 111922
rect 559132 162118 559188 162128
rect 559132 97524 559188 162062
rect 559132 97458 559188 97468
rect 562098 154350 562718 164250
rect 562098 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 562718 154350
rect 562098 154226 562718 154294
rect 562098 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 562718 154226
rect 562098 154102 562718 154170
rect 562098 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 562718 154102
rect 562098 153978 562718 154046
rect 562098 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 562718 153978
rect 562098 136350 562718 153922
rect 581756 153972 581812 406588
rect 589098 400350 589718 417922
rect 590492 562212 590548 562222
rect 590492 409078 590548 562156
rect 590604 549220 590660 567868
rect 590604 549154 590660 549164
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 590716 522564 590772 522574
rect 590492 409012 590548 409022
rect 590604 509348 590660 509358
rect 590604 402418 590660 509292
rect 590716 409618 590772 522508
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 590716 409552 590772 409562
rect 590828 469700 590884 469710
rect 590828 404038 590884 469644
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 590828 403972 590884 403982
rect 590940 430164 590996 430174
rect 590940 402598 590996 430108
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 590940 402532 590996 402542
rect 591164 403318 591220 403328
rect 590604 402352 590660 402362
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 586348 398638 586404 398648
rect 584780 395398 584836 395408
rect 581756 153906 581812 153916
rect 584668 394858 584724 394868
rect 562098 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 562718 136350
rect 562098 136226 562718 136294
rect 562098 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 562718 136226
rect 562098 136102 562718 136170
rect 562098 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 562718 136102
rect 562098 135978 562718 136046
rect 562098 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 562718 135978
rect 562098 118350 562718 135922
rect 562098 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 562718 118350
rect 562098 118226 562718 118294
rect 562098 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 562718 118226
rect 562098 118102 562718 118170
rect 562098 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 562718 118102
rect 562098 117978 562718 118046
rect 562098 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 562718 117978
rect 562098 100350 562718 117922
rect 562098 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 562718 100350
rect 562098 100226 562718 100294
rect 562098 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 562718 100226
rect 562098 100102 562718 100170
rect 562098 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 562718 100102
rect 562098 99978 562718 100046
rect 562098 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 562718 99978
rect 558378 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 558998 94350
rect 558378 94226 558998 94294
rect 558378 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 558998 94226
rect 558378 94102 558998 94170
rect 558378 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 558998 94102
rect 558378 93978 558998 94046
rect 558378 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 558998 93978
rect 554316 70532 554708 70588
rect 558378 76350 558998 93922
rect 558378 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 558998 76350
rect 558378 76226 558998 76294
rect 558378 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 558998 76226
rect 558378 76102 558998 76170
rect 558378 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 558998 76102
rect 558378 75978 558998 76046
rect 558378 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 558998 75978
rect 554316 67732 554372 70532
rect 554316 67666 554372 67676
rect 457996 66434 458052 66444
rect 557788 64596 557844 64606
rect 479808 64350 480128 64384
rect 479808 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 480128 64350
rect 479808 64226 480128 64294
rect 479808 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 480128 64226
rect 479808 64102 480128 64170
rect 479808 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 480128 64102
rect 479808 63978 480128 64046
rect 479808 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 480128 63978
rect 479808 63888 480128 63922
rect 510528 64350 510848 64384
rect 510528 64294 510598 64350
rect 510654 64294 510722 64350
rect 510778 64294 510848 64350
rect 510528 64226 510848 64294
rect 510528 64170 510598 64226
rect 510654 64170 510722 64226
rect 510778 64170 510848 64226
rect 510528 64102 510848 64170
rect 510528 64046 510598 64102
rect 510654 64046 510722 64102
rect 510778 64046 510848 64102
rect 510528 63978 510848 64046
rect 510528 63922 510598 63978
rect 510654 63922 510722 63978
rect 510778 63922 510848 63978
rect 510528 63888 510848 63922
rect 541248 64350 541568 64384
rect 541248 64294 541318 64350
rect 541374 64294 541442 64350
rect 541498 64294 541568 64350
rect 541248 64226 541568 64294
rect 541248 64170 541318 64226
rect 541374 64170 541442 64226
rect 541498 64170 541568 64226
rect 541248 64102 541568 64170
rect 541248 64046 541318 64102
rect 541374 64046 541442 64102
rect 541498 64046 541568 64102
rect 541248 63978 541568 64046
rect 541248 63922 541318 63978
rect 541374 63922 541442 63978
rect 541498 63922 541568 63978
rect 541248 63888 541568 63922
rect 457772 63522 457828 63532
rect 457548 60610 457604 60620
rect 457660 61348 457716 61358
rect 457660 57764 457716 61292
rect 464448 58350 464768 58384
rect 464448 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 464768 58350
rect 464448 58226 464768 58294
rect 464448 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 464768 58226
rect 464448 58102 464768 58170
rect 464448 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 464768 58102
rect 464448 57978 464768 58046
rect 464448 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 464768 57978
rect 464448 57888 464768 57922
rect 495168 58350 495488 58384
rect 495168 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 495488 58350
rect 495168 58226 495488 58294
rect 495168 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 495488 58226
rect 495168 58102 495488 58170
rect 495168 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 495488 58102
rect 495168 57978 495488 58046
rect 495168 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 495488 57978
rect 495168 57888 495488 57922
rect 525888 58350 526208 58384
rect 525888 58294 525958 58350
rect 526014 58294 526082 58350
rect 526138 58294 526208 58350
rect 525888 58226 526208 58294
rect 525888 58170 525958 58226
rect 526014 58170 526082 58226
rect 526138 58170 526208 58226
rect 525888 58102 526208 58170
rect 525888 58046 525958 58102
rect 526014 58046 526082 58102
rect 526138 58046 526208 58102
rect 525888 57978 526208 58046
rect 525888 57922 525958 57978
rect 526014 57922 526082 57978
rect 526138 57922 526208 57978
rect 525888 57888 526208 57922
rect 457660 57698 457716 57708
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 439218 28350 439838 45922
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 439218 10350 439838 27922
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 439218 -1120 439838 9922
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 40350 466838 48914
rect 466218 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 466838 40350
rect 466218 40226 466838 40294
rect 466218 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 466838 40226
rect 466218 40102 466838 40170
rect 466218 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 466838 40102
rect 466218 39978 466838 40046
rect 466218 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 466838 39978
rect 466218 22350 466838 39922
rect 466218 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 466838 22350
rect 466218 22226 466838 22294
rect 466218 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 466838 22226
rect 466218 22102 466838 22170
rect 466218 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 466838 22102
rect 466218 21978 466838 22046
rect 466218 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 466838 21978
rect 466218 4350 466838 21922
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 46350 470558 48914
rect 469938 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 470558 46350
rect 469938 46226 470558 46294
rect 469938 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 470558 46226
rect 469938 46102 470558 46170
rect 469938 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 470558 46102
rect 469938 45978 470558 46046
rect 469938 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 470558 45978
rect 469938 28350 470558 45922
rect 469938 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 470558 28350
rect 469938 28226 470558 28294
rect 469938 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 470558 28226
rect 469938 28102 470558 28170
rect 469938 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 470558 28102
rect 469938 27978 470558 28046
rect 469938 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 470558 27978
rect 469938 10350 470558 27922
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 469938 -1120 470558 9922
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 40350 497558 48914
rect 496938 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 497558 40350
rect 496938 40226 497558 40294
rect 496938 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 497558 40226
rect 496938 40102 497558 40170
rect 496938 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 497558 40102
rect 496938 39978 497558 40046
rect 496938 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 497558 39978
rect 496938 22350 497558 39922
rect 496938 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 497558 22350
rect 496938 22226 497558 22294
rect 496938 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 497558 22226
rect 496938 22102 497558 22170
rect 496938 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 497558 22102
rect 496938 21978 497558 22046
rect 496938 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 497558 21978
rect 496938 4350 497558 21922
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 496938 -160 497558 3922
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 46350 501278 48914
rect 500658 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 501278 46350
rect 500658 46226 501278 46294
rect 500658 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 501278 46226
rect 500658 46102 501278 46170
rect 500658 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 501278 46102
rect 500658 45978 501278 46046
rect 500658 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 501278 45978
rect 500658 28350 501278 45922
rect 500658 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 501278 28350
rect 500658 28226 501278 28294
rect 500658 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 501278 28226
rect 500658 28102 501278 28170
rect 500658 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 501278 28102
rect 500658 27978 501278 28046
rect 500658 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 501278 27978
rect 500658 10350 501278 27922
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 500658 -1120 501278 9922
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 40350 528278 48914
rect 527658 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 528278 40350
rect 527658 40226 528278 40294
rect 527658 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 528278 40226
rect 527658 40102 528278 40170
rect 527658 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 528278 40102
rect 527658 39978 528278 40046
rect 527658 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 528278 39978
rect 527658 22350 528278 39922
rect 527658 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 528278 22350
rect 527658 22226 528278 22294
rect 527658 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 528278 22226
rect 527658 22102 528278 22170
rect 527658 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 528278 22102
rect 527658 21978 528278 22046
rect 527658 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 528278 21978
rect 527658 4350 528278 21922
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 46350 531998 48914
rect 557788 48580 557844 64540
rect 557788 48514 557844 48524
rect 558378 58350 558998 75922
rect 558378 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 558998 58350
rect 558378 58226 558998 58294
rect 558378 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 558998 58226
rect 558378 58102 558998 58170
rect 558378 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 558998 58102
rect 558378 57978 558998 58046
rect 558378 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 558998 57978
rect 531378 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 531998 46350
rect 531378 46226 531998 46294
rect 531378 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 531998 46226
rect 531378 46102 531998 46170
rect 531378 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 531998 46102
rect 531378 45978 531998 46046
rect 531378 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 531998 45978
rect 531378 28350 531998 45922
rect 531378 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 531998 28350
rect 531378 28226 531998 28294
rect 531378 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 531998 28226
rect 531378 28102 531998 28170
rect 531378 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 531998 28102
rect 531378 27978 531998 28046
rect 531378 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 531998 27978
rect 531378 10350 531998 27922
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 531378 -1120 531998 9922
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 40350 558998 57922
rect 558378 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 558998 40350
rect 558378 40226 558998 40294
rect 558378 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 558998 40226
rect 558378 40102 558998 40170
rect 558378 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 558998 40102
rect 558378 39978 558998 40046
rect 558378 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 558998 39978
rect 558378 22350 558998 39922
rect 558378 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 558998 22350
rect 558378 22226 558998 22294
rect 558378 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 558998 22226
rect 558378 22102 558998 22170
rect 558378 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 558998 22102
rect 558378 21978 558998 22046
rect 558378 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 558998 21978
rect 558378 4350 558998 21922
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 558378 -160 558998 3922
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 82350 562718 99922
rect 562098 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 562718 82350
rect 562098 82226 562718 82294
rect 562098 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 562718 82226
rect 562098 82102 562718 82170
rect 562098 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 562718 82102
rect 562098 81978 562718 82046
rect 562098 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 562718 81978
rect 562098 64350 562718 81922
rect 562098 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 562718 64350
rect 562098 64226 562718 64294
rect 562098 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 562718 64226
rect 562098 64102 562718 64170
rect 562098 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 562718 64102
rect 562098 63978 562718 64046
rect 562098 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 562718 63978
rect 562098 46350 562718 63922
rect 562098 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 562718 46350
rect 562098 46226 562718 46294
rect 562098 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 562718 46226
rect 562098 46102 562718 46170
rect 562098 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 562718 46102
rect 562098 45978 562718 46046
rect 562098 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 562718 45978
rect 562098 28350 562718 45922
rect 562098 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 562718 28350
rect 562098 28226 562718 28294
rect 562098 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 562718 28226
rect 562098 28102 562718 28170
rect 562098 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 562718 28102
rect 562098 27978 562718 28046
rect 562098 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 562718 27978
rect 562098 10350 562718 27922
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 562098 -1120 562718 9922
rect 584668 5012 584724 394802
rect 584780 162596 584836 395342
rect 585452 393958 585508 393968
rect 585452 179172 585508 393902
rect 585452 179106 585508 179116
rect 586348 162708 586404 398582
rect 586460 395218 586516 395228
rect 586460 164724 586516 395162
rect 586460 164658 586516 164668
rect 587132 393778 587188 393788
rect 586348 162642 586404 162652
rect 584780 162530 584836 162540
rect 587132 99876 587188 393722
rect 587356 393418 587412 393428
rect 587356 139412 587412 393362
rect 587356 139346 587412 139356
rect 589098 382350 589718 399922
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 589098 364350 589718 381922
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 589098 292350 589718 309922
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 589098 274350 589718 291922
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 589098 256350 589718 273922
rect 590492 400618 590548 400628
rect 590492 258468 590548 400562
rect 591052 398458 591108 398468
rect 590828 398278 590884 398288
rect 590716 394660 590772 394670
rect 590604 393598 590660 393608
rect 590604 298116 590660 393542
rect 590716 311332 590772 394604
rect 590828 337652 590884 398222
rect 591052 350980 591108 398402
rect 591164 390628 591220 403262
rect 591164 390562 591220 390572
rect 592172 401698 592228 401708
rect 591052 350914 591108 350924
rect 590828 337586 590884 337596
rect 590716 311266 590772 311276
rect 590604 298050 590660 298060
rect 590492 258402 590548 258412
rect 590716 271460 590772 271470
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 589098 238350 589718 255922
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 589098 148350 589718 165922
rect 590492 192164 590548 192174
rect 590492 164638 590548 192108
rect 590716 165732 590772 271404
rect 590940 231924 590996 231934
rect 590940 166180 590996 231868
rect 590940 166114 590996 166124
rect 590716 165666 590772 165676
rect 590492 164572 590548 164582
rect 590156 152758 590212 152778
rect 590156 152674 590212 152684
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 587132 99810 587188 99820
rect 589098 130350 589718 147922
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 590492 151318 590548 151328
rect 590492 113092 590548 151262
rect 590492 113026 590548 113036
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 584668 4946 584724 4956
rect 589098 94350 589718 111922
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 589098 76350 589718 93922
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 589098 58350 589718 75922
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 589098 40350 589718 57922
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 589098 22350 589718 39922
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 4350 589718 21922
rect 592172 20580 592228 401642
rect 592284 393238 592340 393248
rect 592284 218820 592340 393182
rect 592284 218754 592340 218764
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 592172 20514 592228 20524
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect 4172 416762 4228 416818
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect 7532 409022 7588 409078
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect 4172 377162 4228 377218
rect 4172 376262 4228 376318
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect 4284 294722 4340 294778
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 36234 597156 36290 597212
rect 36358 597156 36414 597212
rect 36482 597156 36538 597212
rect 36606 597156 36662 597212
rect 36234 597032 36290 597088
rect 36358 597032 36414 597088
rect 36482 597032 36538 597088
rect 36606 597032 36662 597088
rect 36234 596908 36290 596964
rect 36358 596908 36414 596964
rect 36482 596908 36538 596964
rect 36606 596908 36662 596964
rect 36234 596784 36290 596840
rect 36358 596784 36414 596840
rect 36482 596784 36538 596840
rect 36606 596784 36662 596840
rect 36234 580294 36290 580350
rect 36358 580294 36414 580350
rect 36482 580294 36538 580350
rect 36606 580294 36662 580350
rect 36234 580170 36290 580226
rect 36358 580170 36414 580226
rect 36482 580170 36538 580226
rect 36606 580170 36662 580226
rect 36234 580046 36290 580102
rect 36358 580046 36414 580102
rect 36482 580046 36538 580102
rect 36606 580046 36662 580102
rect 36234 579922 36290 579978
rect 36358 579922 36414 579978
rect 36482 579922 36538 579978
rect 36606 579922 36662 579978
rect 36234 562294 36290 562350
rect 36358 562294 36414 562350
rect 36482 562294 36538 562350
rect 36606 562294 36662 562350
rect 36234 562170 36290 562226
rect 36358 562170 36414 562226
rect 36482 562170 36538 562226
rect 36606 562170 36662 562226
rect 36234 562046 36290 562102
rect 36358 562046 36414 562102
rect 36482 562046 36538 562102
rect 36606 562046 36662 562102
rect 36234 561922 36290 561978
rect 36358 561922 36414 561978
rect 36482 561922 36538 561978
rect 36606 561922 36662 561978
rect 36234 544294 36290 544350
rect 36358 544294 36414 544350
rect 36482 544294 36538 544350
rect 36606 544294 36662 544350
rect 36234 544170 36290 544226
rect 36358 544170 36414 544226
rect 36482 544170 36538 544226
rect 36606 544170 36662 544226
rect 36234 544046 36290 544102
rect 36358 544046 36414 544102
rect 36482 544046 36538 544102
rect 36606 544046 36662 544102
rect 36234 543922 36290 543978
rect 36358 543922 36414 543978
rect 36482 543922 36538 543978
rect 36606 543922 36662 543978
rect 36234 526294 36290 526350
rect 36358 526294 36414 526350
rect 36482 526294 36538 526350
rect 36606 526294 36662 526350
rect 36234 526170 36290 526226
rect 36358 526170 36414 526226
rect 36482 526170 36538 526226
rect 36606 526170 36662 526226
rect 36234 526046 36290 526102
rect 36358 526046 36414 526102
rect 36482 526046 36538 526102
rect 36606 526046 36662 526102
rect 36234 525922 36290 525978
rect 36358 525922 36414 525978
rect 36482 525922 36538 525978
rect 36606 525922 36662 525978
rect 36234 508294 36290 508350
rect 36358 508294 36414 508350
rect 36482 508294 36538 508350
rect 36606 508294 36662 508350
rect 36234 508170 36290 508226
rect 36358 508170 36414 508226
rect 36482 508170 36538 508226
rect 36606 508170 36662 508226
rect 36234 508046 36290 508102
rect 36358 508046 36414 508102
rect 36482 508046 36538 508102
rect 36606 508046 36662 508102
rect 36234 507922 36290 507978
rect 36358 507922 36414 507978
rect 36482 507922 36538 507978
rect 36606 507922 36662 507978
rect 36234 490294 36290 490350
rect 36358 490294 36414 490350
rect 36482 490294 36538 490350
rect 36606 490294 36662 490350
rect 36234 490170 36290 490226
rect 36358 490170 36414 490226
rect 36482 490170 36538 490226
rect 36606 490170 36662 490226
rect 36234 490046 36290 490102
rect 36358 490046 36414 490102
rect 36482 490046 36538 490102
rect 36606 490046 36662 490102
rect 36234 489922 36290 489978
rect 36358 489922 36414 489978
rect 36482 489922 36538 489978
rect 36606 489922 36662 489978
rect 36234 472294 36290 472350
rect 36358 472294 36414 472350
rect 36482 472294 36538 472350
rect 36606 472294 36662 472350
rect 36234 472170 36290 472226
rect 36358 472170 36414 472226
rect 36482 472170 36538 472226
rect 36606 472170 36662 472226
rect 36234 472046 36290 472102
rect 36358 472046 36414 472102
rect 36482 472046 36538 472102
rect 36606 472046 36662 472102
rect 36234 471922 36290 471978
rect 36358 471922 36414 471978
rect 36482 471922 36538 471978
rect 36606 471922 36662 471978
rect 36234 454294 36290 454350
rect 36358 454294 36414 454350
rect 36482 454294 36538 454350
rect 36606 454294 36662 454350
rect 36234 454170 36290 454226
rect 36358 454170 36414 454226
rect 36482 454170 36538 454226
rect 36606 454170 36662 454226
rect 36234 454046 36290 454102
rect 36358 454046 36414 454102
rect 36482 454046 36538 454102
rect 36606 454046 36662 454102
rect 36234 453922 36290 453978
rect 36358 453922 36414 453978
rect 36482 453922 36538 453978
rect 36606 453922 36662 453978
rect 36234 436294 36290 436350
rect 36358 436294 36414 436350
rect 36482 436294 36538 436350
rect 36606 436294 36662 436350
rect 36234 436170 36290 436226
rect 36358 436170 36414 436226
rect 36482 436170 36538 436226
rect 36606 436170 36662 436226
rect 36234 436046 36290 436102
rect 36358 436046 36414 436102
rect 36482 436046 36538 436102
rect 36606 436046 36662 436102
rect 36234 435922 36290 435978
rect 36358 435922 36414 435978
rect 36482 435922 36538 435978
rect 36606 435922 36662 435978
rect 36234 418294 36290 418350
rect 36358 418294 36414 418350
rect 36482 418294 36538 418350
rect 36606 418294 36662 418350
rect 36234 418170 36290 418226
rect 36358 418170 36414 418226
rect 36482 418170 36538 418226
rect 36606 418170 36662 418226
rect 36234 418046 36290 418102
rect 36358 418046 36414 418102
rect 36482 418046 36538 418102
rect 36606 418046 36662 418102
rect 36234 417922 36290 417978
rect 36358 417922 36414 417978
rect 36482 417922 36538 417978
rect 36606 417922 36662 417978
rect 36234 400294 36290 400350
rect 36358 400294 36414 400350
rect 36482 400294 36538 400350
rect 36606 400294 36662 400350
rect 36234 400170 36290 400226
rect 36358 400170 36414 400226
rect 36482 400170 36538 400226
rect 36606 400170 36662 400226
rect 36234 400046 36290 400102
rect 36358 400046 36414 400102
rect 36482 400046 36538 400102
rect 36606 400046 36662 400102
rect 36234 399922 36290 399978
rect 36358 399922 36414 399978
rect 36482 399922 36538 399978
rect 36606 399922 36662 399978
rect 36234 382294 36290 382350
rect 36358 382294 36414 382350
rect 36482 382294 36538 382350
rect 36606 382294 36662 382350
rect 36234 382170 36290 382226
rect 36358 382170 36414 382226
rect 36482 382170 36538 382226
rect 36606 382170 36662 382226
rect 36234 382046 36290 382102
rect 36358 382046 36414 382102
rect 36482 382046 36538 382102
rect 36606 382046 36662 382102
rect 36234 381922 36290 381978
rect 36358 381922 36414 381978
rect 36482 381922 36538 381978
rect 36606 381922 36662 381978
rect 31052 378782 31108 378838
rect 29372 377342 29428 377398
rect 9234 370294 9290 370350
rect 9358 370294 9414 370350
rect 9482 370294 9538 370350
rect 9606 370294 9662 370350
rect 9234 370170 9290 370226
rect 9358 370170 9414 370226
rect 9482 370170 9538 370226
rect 9606 370170 9662 370226
rect 9234 370046 9290 370102
rect 9358 370046 9414 370102
rect 9482 370046 9538 370102
rect 9606 370046 9662 370102
rect 9234 369922 9290 369978
rect 9358 369922 9414 369978
rect 9482 369922 9538 369978
rect 9606 369922 9662 369978
rect 9234 352294 9290 352350
rect 9358 352294 9414 352350
rect 9482 352294 9538 352350
rect 9606 352294 9662 352350
rect 9234 352170 9290 352226
rect 9358 352170 9414 352226
rect 9482 352170 9538 352226
rect 9606 352170 9662 352226
rect 9234 352046 9290 352102
rect 9358 352046 9414 352102
rect 9482 352046 9538 352102
rect 9606 352046 9662 352102
rect 9234 351922 9290 351978
rect 9358 351922 9414 351978
rect 9482 351922 9538 351978
rect 9606 351922 9662 351978
rect 9234 334294 9290 334350
rect 9358 334294 9414 334350
rect 9482 334294 9538 334350
rect 9606 334294 9662 334350
rect 9234 334170 9290 334226
rect 9358 334170 9414 334226
rect 9482 334170 9538 334226
rect 9606 334170 9662 334226
rect 9234 334046 9290 334102
rect 9358 334046 9414 334102
rect 9482 334046 9538 334102
rect 9606 334046 9662 334102
rect 9234 333922 9290 333978
rect 9358 333922 9414 333978
rect 9482 333922 9538 333978
rect 9606 333922 9662 333978
rect 9234 316294 9290 316350
rect 9358 316294 9414 316350
rect 9482 316294 9538 316350
rect 9606 316294 9662 316350
rect 9234 316170 9290 316226
rect 9358 316170 9414 316226
rect 9482 316170 9538 316226
rect 9606 316170 9662 316226
rect 9234 316046 9290 316102
rect 9358 316046 9414 316102
rect 9482 316046 9538 316102
rect 9606 316046 9662 316102
rect 9234 315922 9290 315978
rect 9358 315922 9414 315978
rect 9482 315922 9538 315978
rect 9606 315922 9662 315978
rect 9234 298294 9290 298350
rect 9358 298294 9414 298350
rect 9482 298294 9538 298350
rect 9606 298294 9662 298350
rect 9234 298170 9290 298226
rect 9358 298170 9414 298226
rect 9482 298170 9538 298226
rect 9606 298170 9662 298226
rect 9234 298046 9290 298102
rect 9358 298046 9414 298102
rect 9482 298046 9538 298102
rect 9606 298046 9662 298102
rect 9234 297922 9290 297978
rect 9358 297922 9414 297978
rect 9482 297922 9538 297978
rect 9606 297922 9662 297978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 12572 372122 12628 372178
rect 9234 280294 9290 280350
rect 9358 280294 9414 280350
rect 9482 280294 9538 280350
rect 9606 280294 9662 280350
rect 9234 280170 9290 280226
rect 9358 280170 9414 280226
rect 9482 280170 9538 280226
rect 9606 280170 9662 280226
rect 9234 280046 9290 280102
rect 9358 280046 9414 280102
rect 9482 280046 9538 280102
rect 9606 280046 9662 280102
rect 9234 279922 9290 279978
rect 9358 279922 9414 279978
rect 9482 279922 9538 279978
rect 9606 279922 9662 279978
rect 9234 262294 9290 262350
rect 9358 262294 9414 262350
rect 9482 262294 9538 262350
rect 9606 262294 9662 262350
rect 9234 262170 9290 262226
rect 9358 262170 9414 262226
rect 9482 262170 9538 262226
rect 9606 262170 9662 262226
rect 9234 262046 9290 262102
rect 9358 262046 9414 262102
rect 9482 262046 9538 262102
rect 9606 262046 9662 262102
rect 9234 261922 9290 261978
rect 9358 261922 9414 261978
rect 9482 261922 9538 261978
rect 9606 261922 9662 261978
rect 9234 244294 9290 244350
rect 9358 244294 9414 244350
rect 9482 244294 9538 244350
rect 9606 244294 9662 244350
rect 9234 244170 9290 244226
rect 9358 244170 9414 244226
rect 9482 244170 9538 244226
rect 9606 244170 9662 244226
rect 9234 244046 9290 244102
rect 9358 244046 9414 244102
rect 9482 244046 9538 244102
rect 9606 244046 9662 244102
rect 9234 243922 9290 243978
rect 9358 243922 9414 243978
rect 9482 243922 9538 243978
rect 9606 243922 9662 243978
rect 9234 226294 9290 226350
rect 9358 226294 9414 226350
rect 9482 226294 9538 226350
rect 9606 226294 9662 226350
rect 9234 226170 9290 226226
rect 9358 226170 9414 226226
rect 9482 226170 9538 226226
rect 9606 226170 9662 226226
rect 9234 226046 9290 226102
rect 9358 226046 9414 226102
rect 9482 226046 9538 226102
rect 9606 226046 9662 226102
rect 9234 225922 9290 225978
rect 9358 225922 9414 225978
rect 9482 225922 9538 225978
rect 9606 225922 9662 225978
rect 9234 208294 9290 208350
rect 9358 208294 9414 208350
rect 9482 208294 9538 208350
rect 9606 208294 9662 208350
rect 9234 208170 9290 208226
rect 9358 208170 9414 208226
rect 9482 208170 9538 208226
rect 9606 208170 9662 208226
rect 9234 208046 9290 208102
rect 9358 208046 9414 208102
rect 9482 208046 9538 208102
rect 9606 208046 9662 208102
rect 9234 207922 9290 207978
rect 9358 207922 9414 207978
rect 9482 207922 9538 207978
rect 9606 207922 9662 207978
rect 9234 190294 9290 190350
rect 9358 190294 9414 190350
rect 9482 190294 9538 190350
rect 9606 190294 9662 190350
rect 9234 190170 9290 190226
rect 9358 190170 9414 190226
rect 9482 190170 9538 190226
rect 9606 190170 9662 190226
rect 9234 190046 9290 190102
rect 9358 190046 9414 190102
rect 9482 190046 9538 190102
rect 9606 190046 9662 190102
rect 9234 189922 9290 189978
rect 9358 189922 9414 189978
rect 9482 189922 9538 189978
rect 9606 189922 9662 189978
rect 9234 172294 9290 172350
rect 9358 172294 9414 172350
rect 9482 172294 9538 172350
rect 9606 172294 9662 172350
rect 9234 172170 9290 172226
rect 9358 172170 9414 172226
rect 9482 172170 9538 172226
rect 9606 172170 9662 172226
rect 9234 172046 9290 172102
rect 9358 172046 9414 172102
rect 9482 172046 9538 172102
rect 9606 172046 9662 172102
rect 9234 171922 9290 171978
rect 9358 171922 9414 171978
rect 9482 171922 9538 171978
rect 9606 171922 9662 171978
rect 9234 154294 9290 154350
rect 9358 154294 9414 154350
rect 9482 154294 9538 154350
rect 9606 154294 9662 154350
rect 9234 154170 9290 154226
rect 9358 154170 9414 154226
rect 9482 154170 9538 154226
rect 9606 154170 9662 154226
rect 9234 154046 9290 154102
rect 9358 154046 9414 154102
rect 9482 154046 9538 154102
rect 9606 154046 9662 154102
rect 9234 153922 9290 153978
rect 9358 153922 9414 153978
rect 9482 153922 9538 153978
rect 9606 153922 9662 153978
rect 9234 136294 9290 136350
rect 9358 136294 9414 136350
rect 9482 136294 9538 136350
rect 9606 136294 9662 136350
rect 9234 136170 9290 136226
rect 9358 136170 9414 136226
rect 9482 136170 9538 136226
rect 9606 136170 9662 136226
rect 9234 136046 9290 136102
rect 9358 136046 9414 136102
rect 9482 136046 9538 136102
rect 9606 136046 9662 136102
rect 9234 135922 9290 135978
rect 9358 135922 9414 135978
rect 9482 135922 9538 135978
rect 9606 135922 9662 135978
rect 9234 118294 9290 118350
rect 9358 118294 9414 118350
rect 9482 118294 9538 118350
rect 9606 118294 9662 118350
rect 9234 118170 9290 118226
rect 9358 118170 9414 118226
rect 9482 118170 9538 118226
rect 9606 118170 9662 118226
rect 9234 118046 9290 118102
rect 9358 118046 9414 118102
rect 9482 118046 9538 118102
rect 9606 118046 9662 118102
rect 9234 117922 9290 117978
rect 9358 117922 9414 117978
rect 9482 117922 9538 117978
rect 9606 117922 9662 117978
rect 9234 100294 9290 100350
rect 9358 100294 9414 100350
rect 9482 100294 9538 100350
rect 9606 100294 9662 100350
rect 9234 100170 9290 100226
rect 9358 100170 9414 100226
rect 9482 100170 9538 100226
rect 9606 100170 9662 100226
rect 9234 100046 9290 100102
rect 9358 100046 9414 100102
rect 9482 100046 9538 100102
rect 9606 100046 9662 100102
rect 9234 99922 9290 99978
rect 9358 99922 9414 99978
rect 9482 99922 9538 99978
rect 9606 99922 9662 99978
rect 9234 82294 9290 82350
rect 9358 82294 9414 82350
rect 9482 82294 9538 82350
rect 9606 82294 9662 82350
rect 9234 82170 9290 82226
rect 9358 82170 9414 82226
rect 9482 82170 9538 82226
rect 9606 82170 9662 82226
rect 9234 82046 9290 82102
rect 9358 82046 9414 82102
rect 9482 82046 9538 82102
rect 9606 82046 9662 82102
rect 9234 81922 9290 81978
rect 9358 81922 9414 81978
rect 9482 81922 9538 81978
rect 9606 81922 9662 81978
rect 9234 64294 9290 64350
rect 9358 64294 9414 64350
rect 9482 64294 9538 64350
rect 9606 64294 9662 64350
rect 9234 64170 9290 64226
rect 9358 64170 9414 64226
rect 9482 64170 9538 64226
rect 9606 64170 9662 64226
rect 9234 64046 9290 64102
rect 9358 64046 9414 64102
rect 9482 64046 9538 64102
rect 9606 64046 9662 64102
rect 9234 63922 9290 63978
rect 9358 63922 9414 63978
rect 9482 63922 9538 63978
rect 9606 63922 9662 63978
rect 18396 238922 18452 238978
rect 16716 238742 16772 238798
rect 9234 46294 9290 46350
rect 9358 46294 9414 46350
rect 9482 46294 9538 46350
rect 9606 46294 9662 46350
rect 9234 46170 9290 46226
rect 9358 46170 9414 46226
rect 9482 46170 9538 46226
rect 9606 46170 9662 46226
rect 9234 46046 9290 46102
rect 9358 46046 9414 46102
rect 9482 46046 9538 46102
rect 9606 46046 9662 46102
rect 9234 45922 9290 45978
rect 9358 45922 9414 45978
rect 9482 45922 9538 45978
rect 9606 45922 9662 45978
rect 9234 28294 9290 28350
rect 9358 28294 9414 28350
rect 9482 28294 9538 28350
rect 9606 28294 9662 28350
rect 9234 28170 9290 28226
rect 9358 28170 9414 28226
rect 9482 28170 9538 28226
rect 9606 28170 9662 28226
rect 9234 28046 9290 28102
rect 9358 28046 9414 28102
rect 9482 28046 9538 28102
rect 9606 28046 9662 28102
rect 9234 27922 9290 27978
rect 9358 27922 9414 27978
rect 9482 27922 9538 27978
rect 9606 27922 9662 27978
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 21756 234422 21812 234478
rect 26796 234242 26852 234298
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 39954 568294 40010 568350
rect 40078 568294 40134 568350
rect 40202 568294 40258 568350
rect 40326 568294 40382 568350
rect 39954 568170 40010 568226
rect 40078 568170 40134 568226
rect 40202 568170 40258 568226
rect 40326 568170 40382 568226
rect 39954 568046 40010 568102
rect 40078 568046 40134 568102
rect 40202 568046 40258 568102
rect 40326 568046 40382 568102
rect 39954 567922 40010 567978
rect 40078 567922 40134 567978
rect 40202 567922 40258 567978
rect 40326 567922 40382 567978
rect 39954 550294 40010 550350
rect 40078 550294 40134 550350
rect 40202 550294 40258 550350
rect 40326 550294 40382 550350
rect 39954 550170 40010 550226
rect 40078 550170 40134 550226
rect 40202 550170 40258 550226
rect 40326 550170 40382 550226
rect 39954 550046 40010 550102
rect 40078 550046 40134 550102
rect 40202 550046 40258 550102
rect 40326 550046 40382 550102
rect 39954 549922 40010 549978
rect 40078 549922 40134 549978
rect 40202 549922 40258 549978
rect 40326 549922 40382 549978
rect 66954 597156 67010 597212
rect 67078 597156 67134 597212
rect 67202 597156 67258 597212
rect 67326 597156 67382 597212
rect 66954 597032 67010 597088
rect 67078 597032 67134 597088
rect 67202 597032 67258 597088
rect 67326 597032 67382 597088
rect 66954 596908 67010 596964
rect 67078 596908 67134 596964
rect 67202 596908 67258 596964
rect 67326 596908 67382 596964
rect 66954 596784 67010 596840
rect 67078 596784 67134 596840
rect 67202 596784 67258 596840
rect 67326 596784 67382 596840
rect 66954 580294 67010 580350
rect 67078 580294 67134 580350
rect 67202 580294 67258 580350
rect 67326 580294 67382 580350
rect 66954 580170 67010 580226
rect 67078 580170 67134 580226
rect 67202 580170 67258 580226
rect 67326 580170 67382 580226
rect 66954 580046 67010 580102
rect 67078 580046 67134 580102
rect 67202 580046 67258 580102
rect 67326 580046 67382 580102
rect 66954 579922 67010 579978
rect 67078 579922 67134 579978
rect 67202 579922 67258 579978
rect 67326 579922 67382 579978
rect 66954 562294 67010 562350
rect 67078 562294 67134 562350
rect 67202 562294 67258 562350
rect 67326 562294 67382 562350
rect 66954 562170 67010 562226
rect 67078 562170 67134 562226
rect 67202 562170 67258 562226
rect 67326 562170 67382 562226
rect 66954 562046 67010 562102
rect 67078 562046 67134 562102
rect 67202 562046 67258 562102
rect 67326 562046 67382 562102
rect 66954 561922 67010 561978
rect 67078 561922 67134 561978
rect 67202 561922 67258 561978
rect 67326 561922 67382 561978
rect 66954 544294 67010 544350
rect 67078 544294 67134 544350
rect 67202 544294 67258 544350
rect 67326 544294 67382 544350
rect 66954 544170 67010 544226
rect 67078 544170 67134 544226
rect 67202 544170 67258 544226
rect 67326 544170 67382 544226
rect 66954 544046 67010 544102
rect 67078 544046 67134 544102
rect 67202 544046 67258 544102
rect 67326 544046 67382 544102
rect 66954 543922 67010 543978
rect 67078 543922 67134 543978
rect 67202 543922 67258 543978
rect 67326 543922 67382 543978
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 70674 568294 70730 568350
rect 70798 568294 70854 568350
rect 70922 568294 70978 568350
rect 71046 568294 71102 568350
rect 70674 568170 70730 568226
rect 70798 568170 70854 568226
rect 70922 568170 70978 568226
rect 71046 568170 71102 568226
rect 70674 568046 70730 568102
rect 70798 568046 70854 568102
rect 70922 568046 70978 568102
rect 71046 568046 71102 568102
rect 70674 567922 70730 567978
rect 70798 567922 70854 567978
rect 70922 567922 70978 567978
rect 71046 567922 71102 567978
rect 70674 550294 70730 550350
rect 70798 550294 70854 550350
rect 70922 550294 70978 550350
rect 71046 550294 71102 550350
rect 70674 550170 70730 550226
rect 70798 550170 70854 550226
rect 70922 550170 70978 550226
rect 71046 550170 71102 550226
rect 70674 550046 70730 550102
rect 70798 550046 70854 550102
rect 70922 550046 70978 550102
rect 71046 550046 71102 550102
rect 70674 549922 70730 549978
rect 70798 549922 70854 549978
rect 70922 549922 70978 549978
rect 71046 549922 71102 549978
rect 97674 597156 97730 597212
rect 97798 597156 97854 597212
rect 97922 597156 97978 597212
rect 98046 597156 98102 597212
rect 97674 597032 97730 597088
rect 97798 597032 97854 597088
rect 97922 597032 97978 597088
rect 98046 597032 98102 597088
rect 97674 596908 97730 596964
rect 97798 596908 97854 596964
rect 97922 596908 97978 596964
rect 98046 596908 98102 596964
rect 97674 596784 97730 596840
rect 97798 596784 97854 596840
rect 97922 596784 97978 596840
rect 98046 596784 98102 596840
rect 97674 580294 97730 580350
rect 97798 580294 97854 580350
rect 97922 580294 97978 580350
rect 98046 580294 98102 580350
rect 97674 580170 97730 580226
rect 97798 580170 97854 580226
rect 97922 580170 97978 580226
rect 98046 580170 98102 580226
rect 97674 580046 97730 580102
rect 97798 580046 97854 580102
rect 97922 580046 97978 580102
rect 98046 580046 98102 580102
rect 97674 579922 97730 579978
rect 97798 579922 97854 579978
rect 97922 579922 97978 579978
rect 98046 579922 98102 579978
rect 97674 562294 97730 562350
rect 97798 562294 97854 562350
rect 97922 562294 97978 562350
rect 98046 562294 98102 562350
rect 97674 562170 97730 562226
rect 97798 562170 97854 562226
rect 97922 562170 97978 562226
rect 98046 562170 98102 562226
rect 97674 562046 97730 562102
rect 97798 562046 97854 562102
rect 97922 562046 97978 562102
rect 98046 562046 98102 562102
rect 97674 561922 97730 561978
rect 97798 561922 97854 561978
rect 97922 561922 97978 561978
rect 98046 561922 98102 561978
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 159114 597156 159170 597212
rect 159238 597156 159294 597212
rect 159362 597156 159418 597212
rect 159486 597156 159542 597212
rect 159114 597032 159170 597088
rect 159238 597032 159294 597088
rect 159362 597032 159418 597088
rect 159486 597032 159542 597088
rect 159114 596908 159170 596964
rect 159238 596908 159294 596964
rect 159362 596908 159418 596964
rect 159486 596908 159542 596964
rect 159114 596784 159170 596840
rect 159238 596784 159294 596840
rect 159362 596784 159418 596840
rect 159486 596784 159542 596840
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 130346 580007 130402 580063
rect 130470 580007 130526 580063
rect 130594 580007 130650 580063
rect 130718 580007 130774 580063
rect 130346 579883 130402 579939
rect 130470 579883 130526 579939
rect 130594 579883 130650 579939
rect 130718 579883 130774 579939
rect 101394 568294 101450 568350
rect 101518 568294 101574 568350
rect 101642 568294 101698 568350
rect 101766 568294 101822 568350
rect 101394 568170 101450 568226
rect 101518 568170 101574 568226
rect 101642 568170 101698 568226
rect 101766 568170 101822 568226
rect 101394 568046 101450 568102
rect 101518 568046 101574 568102
rect 101642 568046 101698 568102
rect 101766 568046 101822 568102
rect 101394 567922 101450 567978
rect 101518 567922 101574 567978
rect 101642 567922 101698 567978
rect 101766 567922 101822 567978
rect 116228 562216 116284 562272
rect 116352 562216 116408 562272
rect 116476 562216 116532 562272
rect 116600 562216 116656 562272
rect 116724 562216 116780 562272
rect 116848 562216 116904 562272
rect 116972 562216 117028 562272
rect 117096 562216 117152 562272
rect 117220 562216 117276 562272
rect 117344 562216 117400 562272
rect 117468 562216 117524 562272
rect 117592 562216 117648 562272
rect 117716 562216 117772 562272
rect 117840 562216 117896 562272
rect 117964 562216 118020 562272
rect 118088 562216 118144 562272
rect 118212 562216 118268 562272
rect 118336 562216 118392 562272
rect 118460 562216 118516 562272
rect 118584 562216 118640 562272
rect 118708 562216 118764 562272
rect 118832 562216 118888 562272
rect 118956 562216 119012 562272
rect 119080 562216 119136 562272
rect 119204 562216 119260 562272
rect 119328 562216 119384 562272
rect 119452 562216 119508 562272
rect 119576 562216 119632 562272
rect 119700 562216 119756 562272
rect 119824 562216 119880 562272
rect 119948 562216 120004 562272
rect 120072 562216 120128 562272
rect 120196 562216 120252 562272
rect 120320 562216 120376 562272
rect 120444 562216 120500 562272
rect 120568 562216 120624 562272
rect 120692 562216 120748 562272
rect 120816 562216 120872 562272
rect 120940 562216 120996 562272
rect 121064 562216 121120 562272
rect 121188 562216 121244 562272
rect 121312 562216 121368 562272
rect 121436 562216 121492 562272
rect 121560 562216 121616 562272
rect 121684 562216 121740 562272
rect 121808 562216 121864 562272
rect 121932 562216 121988 562272
rect 122056 562216 122112 562272
rect 122180 562216 122236 562272
rect 122304 562216 122360 562272
rect 122428 562216 122484 562272
rect 122552 562216 122608 562272
rect 122676 562216 122732 562272
rect 122800 562216 122856 562272
rect 122924 562216 122980 562272
rect 123048 562216 123104 562272
rect 123172 562216 123228 562272
rect 123296 562216 123352 562272
rect 123420 562216 123476 562272
rect 123544 562216 123600 562272
rect 123668 562216 123724 562272
rect 123792 562216 123848 562272
rect 123916 562216 123972 562272
rect 124040 562216 124096 562272
rect 124164 562216 124220 562272
rect 124288 562216 124344 562272
rect 124412 562216 124468 562272
rect 124536 562216 124592 562272
rect 124660 562216 124716 562272
rect 124784 562216 124840 562272
rect 124908 562216 124964 562272
rect 125032 562216 125088 562272
rect 125156 562216 125212 562272
rect 125280 562216 125336 562272
rect 125404 562216 125460 562272
rect 125528 562216 125584 562272
rect 125652 562216 125708 562272
rect 125776 562216 125832 562272
rect 125900 562216 125956 562272
rect 126024 562216 126080 562272
rect 126148 562216 126204 562272
rect 126272 562216 126328 562272
rect 126396 562216 126452 562272
rect 126520 562216 126576 562272
rect 126644 562216 126700 562272
rect 126768 562216 126824 562272
rect 126892 562216 126948 562272
rect 127016 562216 127072 562272
rect 127140 562216 127196 562272
rect 127264 562216 127320 562272
rect 127388 562216 127444 562272
rect 127512 562216 127568 562272
rect 127636 562216 127692 562272
rect 127760 562216 127816 562272
rect 127884 562216 127940 562272
rect 128008 562216 128064 562272
rect 128132 562216 128188 562272
rect 128256 562216 128312 562272
rect 128380 562216 128436 562272
rect 128504 562216 128560 562272
rect 128628 562216 128684 562272
rect 128752 562216 128808 562272
rect 128876 562216 128932 562272
rect 129000 562216 129056 562272
rect 129124 562216 129180 562272
rect 129248 562216 129304 562272
rect 129372 562216 129428 562272
rect 129496 562216 129552 562272
rect 129620 562216 129676 562272
rect 129744 562216 129800 562272
rect 129868 562216 129924 562272
rect 129992 562216 130048 562272
rect 130116 562216 130172 562272
rect 130240 562216 130296 562272
rect 130364 562216 130420 562272
rect 130488 562216 130544 562272
rect 130612 562216 130668 562272
rect 130736 562216 130792 562272
rect 130860 562216 130916 562272
rect 130984 562216 131040 562272
rect 131108 562216 131164 562272
rect 131232 562216 131288 562272
rect 131356 562216 131412 562272
rect 131480 562216 131536 562272
rect 131604 562216 131660 562272
rect 131728 562216 131784 562272
rect 131852 562216 131908 562272
rect 131976 562216 132032 562272
rect 132100 562216 132156 562272
rect 132224 562216 132280 562272
rect 132348 562216 132404 562272
rect 132472 562216 132528 562272
rect 132596 562216 132652 562272
rect 116228 562092 116284 562148
rect 116352 562092 116408 562148
rect 116476 562092 116532 562148
rect 116600 562092 116656 562148
rect 116724 562092 116780 562148
rect 116848 562092 116904 562148
rect 116972 562092 117028 562148
rect 117096 562092 117152 562148
rect 117220 562092 117276 562148
rect 117344 562092 117400 562148
rect 117468 562092 117524 562148
rect 117592 562092 117648 562148
rect 117716 562092 117772 562148
rect 117840 562092 117896 562148
rect 117964 562092 118020 562148
rect 118088 562092 118144 562148
rect 118212 562092 118268 562148
rect 118336 562092 118392 562148
rect 118460 562092 118516 562148
rect 118584 562092 118640 562148
rect 118708 562092 118764 562148
rect 118832 562092 118888 562148
rect 118956 562092 119012 562148
rect 119080 562092 119136 562148
rect 119204 562092 119260 562148
rect 119328 562092 119384 562148
rect 119452 562092 119508 562148
rect 119576 562092 119632 562148
rect 119700 562092 119756 562148
rect 119824 562092 119880 562148
rect 119948 562092 120004 562148
rect 120072 562092 120128 562148
rect 120196 562092 120252 562148
rect 120320 562092 120376 562148
rect 120444 562092 120500 562148
rect 120568 562092 120624 562148
rect 120692 562092 120748 562148
rect 120816 562092 120872 562148
rect 120940 562092 120996 562148
rect 121064 562092 121120 562148
rect 121188 562092 121244 562148
rect 121312 562092 121368 562148
rect 121436 562092 121492 562148
rect 121560 562092 121616 562148
rect 121684 562092 121740 562148
rect 121808 562092 121864 562148
rect 121932 562092 121988 562148
rect 122056 562092 122112 562148
rect 122180 562092 122236 562148
rect 122304 562092 122360 562148
rect 122428 562092 122484 562148
rect 122552 562092 122608 562148
rect 122676 562092 122732 562148
rect 122800 562092 122856 562148
rect 122924 562092 122980 562148
rect 123048 562092 123104 562148
rect 123172 562092 123228 562148
rect 123296 562092 123352 562148
rect 123420 562092 123476 562148
rect 123544 562092 123600 562148
rect 123668 562092 123724 562148
rect 123792 562092 123848 562148
rect 123916 562092 123972 562148
rect 124040 562092 124096 562148
rect 124164 562092 124220 562148
rect 124288 562092 124344 562148
rect 124412 562092 124468 562148
rect 124536 562092 124592 562148
rect 124660 562092 124716 562148
rect 124784 562092 124840 562148
rect 124908 562092 124964 562148
rect 125032 562092 125088 562148
rect 125156 562092 125212 562148
rect 125280 562092 125336 562148
rect 125404 562092 125460 562148
rect 125528 562092 125584 562148
rect 125652 562092 125708 562148
rect 125776 562092 125832 562148
rect 125900 562092 125956 562148
rect 126024 562092 126080 562148
rect 126148 562092 126204 562148
rect 126272 562092 126328 562148
rect 126396 562092 126452 562148
rect 126520 562092 126576 562148
rect 126644 562092 126700 562148
rect 126768 562092 126824 562148
rect 126892 562092 126948 562148
rect 127016 562092 127072 562148
rect 127140 562092 127196 562148
rect 127264 562092 127320 562148
rect 127388 562092 127444 562148
rect 127512 562092 127568 562148
rect 127636 562092 127692 562148
rect 127760 562092 127816 562148
rect 127884 562092 127940 562148
rect 128008 562092 128064 562148
rect 128132 562092 128188 562148
rect 128256 562092 128312 562148
rect 128380 562092 128436 562148
rect 128504 562092 128560 562148
rect 128628 562092 128684 562148
rect 128752 562092 128808 562148
rect 128876 562092 128932 562148
rect 129000 562092 129056 562148
rect 129124 562092 129180 562148
rect 129248 562092 129304 562148
rect 129372 562092 129428 562148
rect 129496 562092 129552 562148
rect 129620 562092 129676 562148
rect 129744 562092 129800 562148
rect 129868 562092 129924 562148
rect 129992 562092 130048 562148
rect 130116 562092 130172 562148
rect 130240 562092 130296 562148
rect 130364 562092 130420 562148
rect 130488 562092 130544 562148
rect 130612 562092 130668 562148
rect 130736 562092 130792 562148
rect 130860 562092 130916 562148
rect 130984 562092 131040 562148
rect 131108 562092 131164 562148
rect 131232 562092 131288 562148
rect 131356 562092 131412 562148
rect 131480 562092 131536 562148
rect 131604 562092 131660 562148
rect 131728 562092 131784 562148
rect 131852 562092 131908 562148
rect 131976 562092 132032 562148
rect 132100 562092 132156 562148
rect 132224 562092 132280 562148
rect 132348 562092 132404 562148
rect 132472 562092 132528 562148
rect 132596 562092 132652 562148
rect 116228 561968 116284 562024
rect 116352 561968 116408 562024
rect 116476 561968 116532 562024
rect 116600 561968 116656 562024
rect 116724 561968 116780 562024
rect 116848 561968 116904 562024
rect 116972 561968 117028 562024
rect 117096 561968 117152 562024
rect 117220 561968 117276 562024
rect 117344 561968 117400 562024
rect 117468 561968 117524 562024
rect 117592 561968 117648 562024
rect 117716 561968 117772 562024
rect 117840 561968 117896 562024
rect 117964 561968 118020 562024
rect 118088 561968 118144 562024
rect 118212 561968 118268 562024
rect 118336 561968 118392 562024
rect 118460 561968 118516 562024
rect 118584 561968 118640 562024
rect 118708 561968 118764 562024
rect 118832 561968 118888 562024
rect 118956 561968 119012 562024
rect 119080 561968 119136 562024
rect 119204 561968 119260 562024
rect 119328 561968 119384 562024
rect 119452 561968 119508 562024
rect 119576 561968 119632 562024
rect 119700 561968 119756 562024
rect 119824 561968 119880 562024
rect 119948 561968 120004 562024
rect 120072 561968 120128 562024
rect 120196 561968 120252 562024
rect 120320 561968 120376 562024
rect 120444 561968 120500 562024
rect 120568 561968 120624 562024
rect 120692 561968 120748 562024
rect 120816 561968 120872 562024
rect 120940 561968 120996 562024
rect 121064 561968 121120 562024
rect 121188 561968 121244 562024
rect 121312 561968 121368 562024
rect 121436 561968 121492 562024
rect 121560 561968 121616 562024
rect 121684 561968 121740 562024
rect 121808 561968 121864 562024
rect 121932 561968 121988 562024
rect 122056 561968 122112 562024
rect 122180 561968 122236 562024
rect 122304 561968 122360 562024
rect 122428 561968 122484 562024
rect 122552 561968 122608 562024
rect 122676 561968 122732 562024
rect 122800 561968 122856 562024
rect 122924 561968 122980 562024
rect 123048 561968 123104 562024
rect 123172 561968 123228 562024
rect 123296 561968 123352 562024
rect 123420 561968 123476 562024
rect 123544 561968 123600 562024
rect 123668 561968 123724 562024
rect 123792 561968 123848 562024
rect 123916 561968 123972 562024
rect 124040 561968 124096 562024
rect 124164 561968 124220 562024
rect 124288 561968 124344 562024
rect 124412 561968 124468 562024
rect 124536 561968 124592 562024
rect 124660 561968 124716 562024
rect 124784 561968 124840 562024
rect 124908 561968 124964 562024
rect 125032 561968 125088 562024
rect 125156 561968 125212 562024
rect 125280 561968 125336 562024
rect 125404 561968 125460 562024
rect 125528 561968 125584 562024
rect 125652 561968 125708 562024
rect 125776 561968 125832 562024
rect 125900 561968 125956 562024
rect 126024 561968 126080 562024
rect 126148 561968 126204 562024
rect 126272 561968 126328 562024
rect 126396 561968 126452 562024
rect 126520 561968 126576 562024
rect 126644 561968 126700 562024
rect 126768 561968 126824 562024
rect 126892 561968 126948 562024
rect 127016 561968 127072 562024
rect 127140 561968 127196 562024
rect 127264 561968 127320 562024
rect 127388 561968 127444 562024
rect 127512 561968 127568 562024
rect 127636 561968 127692 562024
rect 127760 561968 127816 562024
rect 127884 561968 127940 562024
rect 128008 561968 128064 562024
rect 128132 561968 128188 562024
rect 128256 561968 128312 562024
rect 128380 561968 128436 562024
rect 128504 561968 128560 562024
rect 128628 561968 128684 562024
rect 128752 561968 128808 562024
rect 128876 561968 128932 562024
rect 129000 561968 129056 562024
rect 129124 561968 129180 562024
rect 129248 561968 129304 562024
rect 129372 561968 129428 562024
rect 129496 561968 129552 562024
rect 129620 561968 129676 562024
rect 129744 561968 129800 562024
rect 129868 561968 129924 562024
rect 129992 561968 130048 562024
rect 130116 561968 130172 562024
rect 130240 561968 130296 562024
rect 130364 561968 130420 562024
rect 130488 561968 130544 562024
rect 130612 561968 130668 562024
rect 130736 561968 130792 562024
rect 130860 561968 130916 562024
rect 130984 561968 131040 562024
rect 131108 561968 131164 562024
rect 131232 561968 131288 562024
rect 131356 561968 131412 562024
rect 131480 561968 131536 562024
rect 131604 561968 131660 562024
rect 131728 561968 131784 562024
rect 131852 561968 131908 562024
rect 131976 561968 132032 562024
rect 132100 561968 132156 562024
rect 132224 561968 132280 562024
rect 132348 561968 132404 562024
rect 132472 561968 132528 562024
rect 132596 561968 132652 562024
rect 101394 550294 101450 550350
rect 101518 550294 101574 550350
rect 101642 550294 101698 550350
rect 101766 550294 101822 550350
rect 101394 550170 101450 550226
rect 101518 550170 101574 550226
rect 101642 550170 101698 550226
rect 101766 550170 101822 550226
rect 101394 550046 101450 550102
rect 101518 550046 101574 550102
rect 101642 550046 101698 550102
rect 101766 550046 101822 550102
rect 101394 549922 101450 549978
rect 101518 549922 101574 549978
rect 101642 549922 101698 549978
rect 101766 549922 101822 549978
rect 104348 544002 104404 544058
rect 104472 544002 104528 544058
rect 104596 544002 104652 544058
rect 104720 544002 104776 544058
rect 104844 544002 104900 544058
rect 104968 544002 105024 544058
rect 105092 544002 105148 544058
rect 105216 544002 105272 544058
rect 105340 544002 105396 544058
rect 105464 544002 105520 544058
rect 105588 544002 105644 544058
rect 105712 544002 105768 544058
rect 105836 544002 105892 544058
rect 105960 544002 106016 544058
rect 106084 544002 106140 544058
rect 106208 544002 106264 544058
rect 106332 544002 106388 544058
rect 106456 544002 106512 544058
rect 106580 544002 106636 544058
rect 106704 544002 106760 544058
rect 106828 544002 106884 544058
rect 106952 544002 107008 544058
rect 107076 544002 107132 544058
rect 107200 544002 107256 544058
rect 107324 544002 107380 544058
rect 107448 544002 107504 544058
rect 107572 544002 107628 544058
rect 107696 544002 107752 544058
rect 107820 544002 107876 544058
rect 107944 544002 108000 544058
rect 108068 544002 108124 544058
rect 108192 544002 108248 544058
rect 108316 544002 108372 544058
rect 108440 544002 108496 544058
rect 108564 544002 108620 544058
rect 108688 544002 108744 544058
rect 108812 544002 108868 544058
rect 108936 544002 108992 544058
rect 109060 544002 109116 544058
rect 109184 544002 109240 544058
rect 109308 544002 109364 544058
rect 109432 544002 109488 544058
rect 109556 544002 109612 544058
rect 109680 544002 109736 544058
rect 109804 544002 109860 544058
rect 109928 544002 109984 544058
rect 110052 544002 110108 544058
rect 110176 544002 110232 544058
rect 110300 544002 110356 544058
rect 110424 544002 110480 544058
rect 110548 544002 110604 544058
rect 110672 544002 110728 544058
rect 110796 544002 110852 544058
rect 110920 544002 110976 544058
rect 111044 544002 111100 544058
rect 111168 544002 111224 544058
rect 111292 544002 111348 544058
rect 111416 544002 111472 544058
rect 111540 544002 111596 544058
rect 111664 544002 111720 544058
rect 111788 544002 111844 544058
rect 111912 544002 111968 544058
rect 112036 544002 112092 544058
rect 112160 544002 112216 544058
rect 112284 544002 112340 544058
rect 112408 544002 112464 544058
rect 112532 544002 112588 544058
rect 112656 544002 112712 544058
rect 112780 544002 112836 544058
rect 112904 544002 112960 544058
rect 113028 544002 113084 544058
rect 113152 544002 113208 544058
rect 113276 544002 113332 544058
rect 113400 544002 113456 544058
rect 113524 544002 113580 544058
rect 113648 544002 113704 544058
rect 113772 544002 113828 544058
rect 113896 544002 113952 544058
rect 114020 544002 114076 544058
rect 114144 544002 114200 544058
rect 114268 544002 114324 544058
rect 114392 544002 114448 544058
rect 114516 544002 114572 544058
rect 114640 544002 114696 544058
rect 114764 544002 114820 544058
rect 114888 544002 114944 544058
rect 115012 544002 115068 544058
rect 115136 544002 115192 544058
rect 115260 544002 115316 544058
rect 115384 544002 115440 544058
rect 115508 544002 115564 544058
rect 115632 544002 115688 544058
rect 115756 544002 115812 544058
rect 115880 544002 115936 544058
rect 116004 544002 116060 544058
rect 116128 544002 116184 544058
rect 116252 544002 116308 544058
rect 116376 544002 116432 544058
rect 116500 544002 116556 544058
rect 116624 544002 116680 544058
rect 116748 544002 116804 544058
rect 116872 544002 116928 544058
rect 116996 544002 117052 544058
rect 117120 544002 117176 544058
rect 117244 544002 117300 544058
rect 117368 544002 117424 544058
rect 117492 544002 117548 544058
rect 117616 544002 117672 544058
rect 117740 544002 117796 544058
rect 117864 544002 117920 544058
rect 117988 544002 118044 544058
rect 118112 544002 118168 544058
rect 118236 544002 118292 544058
rect 118360 544002 118416 544058
rect 118484 544002 118540 544058
rect 118608 544002 118664 544058
rect 118732 544002 118788 544058
rect 118856 544002 118912 544058
rect 118980 544002 119036 544058
rect 119104 544002 119160 544058
rect 119228 544002 119284 544058
rect 119352 544002 119408 544058
rect 119476 544002 119532 544058
rect 119600 544002 119656 544058
rect 119724 544002 119780 544058
rect 119848 544002 119904 544058
rect 119972 544002 120028 544058
rect 120096 544002 120152 544058
rect 120220 544002 120276 544058
rect 120344 544002 120400 544058
rect 120468 544002 120524 544058
rect 120592 544002 120648 544058
rect 120716 544002 120772 544058
rect 120840 544002 120896 544058
rect 120964 544002 121020 544058
rect 121088 544002 121144 544058
rect 121212 544002 121268 544058
rect 121336 544002 121392 544058
rect 121460 544002 121516 544058
rect 121584 544002 121640 544058
rect 121708 544002 121764 544058
rect 121832 544002 121888 544058
rect 121956 544002 122012 544058
rect 122080 544002 122136 544058
rect 122204 544002 122260 544058
rect 122328 544002 122384 544058
rect 122452 544002 122508 544058
rect 122576 544002 122632 544058
rect 122700 544002 122756 544058
rect 122824 544002 122880 544058
rect 122948 544002 123004 544058
rect 123072 544002 123128 544058
rect 123196 544002 123252 544058
rect 123320 544002 123376 544058
rect 123444 544002 123500 544058
rect 123568 544002 123624 544058
rect 123692 544002 123748 544058
rect 123816 544002 123872 544058
rect 123940 544002 123996 544058
rect 124064 544002 124120 544058
rect 124188 544002 124244 544058
rect 124312 544002 124368 544058
rect 124436 544002 124492 544058
rect 124560 544002 124616 544058
rect 124684 544002 124740 544058
rect 124808 544002 124864 544058
rect 124932 544002 124988 544058
rect 125056 544002 125112 544058
rect 125180 544002 125236 544058
rect 125304 544002 125360 544058
rect 125428 544002 125484 544058
rect 125552 544002 125608 544058
rect 125676 544002 125732 544058
rect 125800 544002 125856 544058
rect 125924 544002 125980 544058
rect 126048 544002 126104 544058
rect 126172 544002 126228 544058
rect 126296 544002 126352 544058
rect 39954 532294 40010 532350
rect 40078 532294 40134 532350
rect 40202 532294 40258 532350
rect 40326 532294 40382 532350
rect 66714 532302 66770 532358
rect 66838 532302 66894 532358
rect 66962 532302 67018 532358
rect 67086 532302 67142 532358
rect 67210 532302 67266 532358
rect 67334 532302 67390 532358
rect 67458 532302 67514 532358
rect 67582 532302 67638 532358
rect 67706 532302 67762 532358
rect 67830 532302 67886 532358
rect 67954 532302 68010 532358
rect 68078 532302 68134 532358
rect 68202 532302 68258 532358
rect 68326 532302 68382 532358
rect 68450 532302 68506 532358
rect 68574 532302 68630 532358
rect 68698 532302 68754 532358
rect 68822 532302 68878 532358
rect 68946 532302 69002 532358
rect 69070 532302 69126 532358
rect 69194 532302 69250 532358
rect 69318 532302 69374 532358
rect 69442 532302 69498 532358
rect 69566 532302 69622 532358
rect 69690 532302 69746 532358
rect 69814 532302 69870 532358
rect 69938 532302 69994 532358
rect 70062 532302 70118 532358
rect 70186 532302 70242 532358
rect 70310 532302 70366 532358
rect 70434 532302 70490 532358
rect 70558 532302 70614 532358
rect 70682 532302 70738 532358
rect 70806 532302 70862 532358
rect 70930 532302 70986 532358
rect 71054 532302 71110 532358
rect 71178 532302 71234 532358
rect 71302 532302 71358 532358
rect 71426 532302 71482 532358
rect 71550 532302 71606 532358
rect 71674 532302 71730 532358
rect 71798 532302 71854 532358
rect 71922 532302 71978 532358
rect 72046 532302 72102 532358
rect 72170 532302 72226 532358
rect 72294 532302 72350 532358
rect 72418 532302 72474 532358
rect 72542 532302 72598 532358
rect 72666 532302 72722 532358
rect 72790 532302 72846 532358
rect 72914 532302 72970 532358
rect 73038 532302 73094 532358
rect 73162 532302 73218 532358
rect 73286 532302 73342 532358
rect 73410 532302 73466 532358
rect 73534 532302 73590 532358
rect 73658 532302 73714 532358
rect 73782 532302 73838 532358
rect 73906 532302 73962 532358
rect 74030 532302 74086 532358
rect 74154 532302 74210 532358
rect 74278 532302 74334 532358
rect 74402 532302 74458 532358
rect 74526 532302 74582 532358
rect 74650 532302 74706 532358
rect 39954 532170 40010 532226
rect 40078 532170 40134 532226
rect 40202 532170 40258 532226
rect 40326 532170 40382 532226
rect 39954 532046 40010 532102
rect 40078 532046 40134 532102
rect 40202 532046 40258 532102
rect 40326 532046 40382 532102
rect 39954 531922 40010 531978
rect 40078 531922 40134 531978
rect 40202 531922 40258 531978
rect 40326 531922 40382 531978
rect 66506 531942 66562 531998
rect 66630 531942 66686 531998
rect 66754 531942 66810 531998
rect 66878 531942 66934 531998
rect 67002 531942 67058 531998
rect 67126 531942 67182 531998
rect 67250 531942 67306 531998
rect 67374 531942 67430 531998
rect 67498 531942 67554 531998
rect 67622 531942 67678 531998
rect 67746 531942 67802 531998
rect 67870 531942 67926 531998
rect 67994 531942 68050 531998
rect 68118 531942 68174 531998
rect 68242 531942 68298 531998
rect 68366 531942 68422 531998
rect 68490 531942 68546 531998
rect 68614 531942 68670 531998
rect 68738 531942 68794 531998
rect 68862 531942 68918 531998
rect 68986 531942 69042 531998
rect 69110 531942 69166 531998
rect 69234 531942 69290 531998
rect 69358 531942 69414 531998
rect 69482 531942 69538 531998
rect 69606 531942 69662 531998
rect 69730 531942 69786 531998
rect 69854 531942 69910 531998
rect 69978 531942 70034 531998
rect 70102 531942 70158 531998
rect 70226 531942 70282 531998
rect 70350 531942 70406 531998
rect 70474 531942 70530 531998
rect 70598 531942 70654 531998
rect 70722 531942 70778 531998
rect 70846 531942 70902 531998
rect 70970 531942 71026 531998
rect 71094 531942 71150 531998
rect 71218 531942 71274 531998
rect 71342 531942 71398 531998
rect 71466 531942 71522 531998
rect 71590 531942 71646 531998
rect 71714 531942 71770 531998
rect 71838 531942 71894 531998
rect 71962 531942 72018 531998
rect 72086 531942 72142 531998
rect 72210 531942 72266 531998
rect 72334 531942 72390 531998
rect 72458 531942 72514 531998
rect 72582 531942 72638 531998
rect 72706 531942 72762 531998
rect 72830 531942 72886 531998
rect 72954 531942 73010 531998
rect 73078 531942 73134 531998
rect 73202 531942 73258 531998
rect 73326 531942 73382 531998
rect 73450 531942 73506 531998
rect 73574 531942 73630 531998
rect 73698 531942 73754 531998
rect 73822 531942 73878 531998
rect 73946 531942 74002 531998
rect 74070 531942 74126 531998
rect 74194 531942 74250 531998
rect 74318 531942 74374 531998
rect 96026 526182 96082 526238
rect 96150 526182 96206 526238
rect 96274 526182 96330 526238
rect 96398 526182 96454 526238
rect 96522 526182 96578 526238
rect 96646 526182 96702 526238
rect 96770 526182 96826 526238
rect 96894 526182 96950 526238
rect 97018 526182 97074 526238
rect 97142 526182 97198 526238
rect 97266 526182 97322 526238
rect 97390 526182 97446 526238
rect 97514 526182 97570 526238
rect 97638 526182 97694 526238
rect 97762 526182 97818 526238
rect 97886 526182 97942 526238
rect 98010 526182 98066 526238
rect 98134 526182 98190 526238
rect 98258 526182 98314 526238
rect 98382 526182 98438 526238
rect 98506 526182 98562 526238
rect 98630 526182 98686 526238
rect 98754 526182 98810 526238
rect 98878 526182 98934 526238
rect 99002 526182 99058 526238
rect 99126 526182 99182 526238
rect 99250 526182 99306 526238
rect 99374 526182 99430 526238
rect 99498 526182 99554 526238
rect 99622 526182 99678 526238
rect 99746 526182 99802 526238
rect 99870 526182 99926 526238
rect 99994 526182 100050 526238
rect 100118 526182 100174 526238
rect 100242 526182 100298 526238
rect 100366 526182 100422 526238
rect 100490 526182 100546 526238
rect 100614 526182 100670 526238
rect 100738 526182 100794 526238
rect 100862 526182 100918 526238
rect 100986 526182 101042 526238
rect 101110 526182 101166 526238
rect 101234 526182 101290 526238
rect 101358 526182 101414 526238
rect 101482 526182 101538 526238
rect 101606 526182 101662 526238
rect 101730 526182 101786 526238
rect 101854 526182 101910 526238
rect 101978 526182 102034 526238
rect 102102 526182 102158 526238
rect 102226 526182 102282 526238
rect 102350 526182 102406 526238
rect 102474 526182 102530 526238
rect 102598 526182 102654 526238
rect 102722 526182 102778 526238
rect 102846 526182 102902 526238
rect 102970 526182 103026 526238
rect 103094 526182 103150 526238
rect 103218 526182 103274 526238
rect 103342 526182 103398 526238
rect 103466 526182 103522 526238
rect 103590 526182 103646 526238
rect 103714 526182 103770 526238
rect 103838 526182 103894 526238
rect 103962 526182 104018 526238
rect 104086 526182 104142 526238
rect 104210 526182 104266 526238
rect 104334 526182 104390 526238
rect 104458 526182 104514 526238
rect 104582 526182 104638 526238
rect 104706 526182 104762 526238
rect 104830 526182 104886 526238
rect 104954 526182 105010 526238
rect 105078 526182 105134 526238
rect 105202 526182 105258 526238
rect 105326 526182 105382 526238
rect 105450 526182 105506 526238
rect 105574 526182 105630 526238
rect 105698 526182 105754 526238
rect 105822 526182 105878 526238
rect 105946 526182 106002 526238
rect 106070 526182 106126 526238
rect 106194 526182 106250 526238
rect 106318 526182 106374 526238
rect 106442 526182 106498 526238
rect 106566 526182 106622 526238
rect 106690 526182 106746 526238
rect 106814 526182 106870 526238
rect 106938 526182 106994 526238
rect 107062 526182 107118 526238
rect 107186 526182 107242 526238
rect 107310 526182 107366 526238
rect 107434 526182 107490 526238
rect 107558 526182 107614 526238
rect 107682 526182 107738 526238
rect 107806 526182 107862 526238
rect 107930 526182 107986 526238
rect 108054 526182 108110 526238
rect 108178 526182 108234 526238
rect 108302 526182 108358 526238
rect 108426 526182 108482 526238
rect 108550 526182 108606 526238
rect 108674 526182 108730 526238
rect 108798 526182 108854 526238
rect 108922 526182 108978 526238
rect 109046 526182 109102 526238
rect 109170 526182 109226 526238
rect 109294 526182 109350 526238
rect 109418 526182 109474 526238
rect 109542 526182 109598 526238
rect 109666 526182 109722 526238
rect 109790 526182 109846 526238
rect 109914 526182 109970 526238
rect 110038 526182 110094 526238
rect 110162 526182 110218 526238
rect 110286 526182 110342 526238
rect 110410 526182 110466 526238
rect 110534 526182 110590 526238
rect 110658 526182 110714 526238
rect 110782 526182 110838 526238
rect 110906 526182 110962 526238
rect 111030 526182 111086 526238
rect 111154 526182 111210 526238
rect 111278 526182 111334 526238
rect 111402 526182 111458 526238
rect 111526 526182 111582 526238
rect 111650 526182 111706 526238
rect 111774 526182 111830 526238
rect 111898 526182 111954 526238
rect 112022 526182 112078 526238
rect 112146 526182 112202 526238
rect 112270 526182 112326 526238
rect 112394 526182 112450 526238
rect 112518 526182 112574 526238
rect 112642 526182 112698 526238
rect 112766 526182 112822 526238
rect 112890 526182 112946 526238
rect 113014 526182 113070 526238
rect 113138 526182 113194 526238
rect 113262 526182 113318 526238
rect 113386 526182 113442 526238
rect 113510 526182 113566 526238
rect 113634 526182 113690 526238
rect 113758 526182 113814 526238
rect 113882 526182 113938 526238
rect 114006 526182 114062 526238
rect 114130 526182 114186 526238
rect 114254 526182 114310 526238
rect 114378 526182 114434 526238
rect 114502 526182 114558 526238
rect 114626 526182 114682 526238
rect 114750 526182 114806 526238
rect 114874 526182 114930 526238
rect 114998 526182 115054 526238
rect 95880 525855 95936 525911
rect 96004 525855 96060 525911
rect 96128 525855 96184 525911
rect 96252 525855 96308 525911
rect 96376 525855 96432 525911
rect 96500 525855 96556 525911
rect 96624 525855 96680 525911
rect 96748 525855 96804 525911
rect 96872 525855 96928 525911
rect 96996 525855 97052 525911
rect 97120 525855 97176 525911
rect 97244 525855 97300 525911
rect 97368 525855 97424 525911
rect 97492 525855 97548 525911
rect 97616 525855 97672 525911
rect 97740 525855 97796 525911
rect 97864 525855 97920 525911
rect 97988 525855 98044 525911
rect 98112 525855 98168 525911
rect 98236 525855 98292 525911
rect 98360 525855 98416 525911
rect 98484 525855 98540 525911
rect 98608 525855 98664 525911
rect 98732 525855 98788 525911
rect 98856 525855 98912 525911
rect 98980 525855 99036 525911
rect 99104 525855 99160 525911
rect 99228 525855 99284 525911
rect 99352 525855 99408 525911
rect 99476 525855 99532 525911
rect 99600 525855 99656 525911
rect 99724 525855 99780 525911
rect 99848 525855 99904 525911
rect 99972 525855 100028 525911
rect 100096 525855 100152 525911
rect 100220 525855 100276 525911
rect 100344 525855 100400 525911
rect 100468 525855 100524 525911
rect 100592 525855 100648 525911
rect 100716 525855 100772 525911
rect 100840 525855 100896 525911
rect 100964 525855 101020 525911
rect 101088 525855 101144 525911
rect 101212 525855 101268 525911
rect 101336 525855 101392 525911
rect 101460 525855 101516 525911
rect 101584 525855 101640 525911
rect 101708 525855 101764 525911
rect 101832 525855 101888 525911
rect 101956 525855 102012 525911
rect 102080 525855 102136 525911
rect 102204 525855 102260 525911
rect 102328 525855 102384 525911
rect 102452 525855 102508 525911
rect 102576 525855 102632 525911
rect 102700 525855 102756 525911
rect 102824 525855 102880 525911
rect 102948 525855 103004 525911
rect 103072 525855 103128 525911
rect 103196 525855 103252 525911
rect 103320 525855 103376 525911
rect 103444 525855 103500 525911
rect 103568 525855 103624 525911
rect 103692 525855 103748 525911
rect 103816 525855 103872 525911
rect 103940 525855 103996 525911
rect 104064 525855 104120 525911
rect 104188 525855 104244 525911
rect 104312 525855 104368 525911
rect 104436 525855 104492 525911
rect 104560 525855 104616 525911
rect 104684 525855 104740 525911
rect 104808 525855 104864 525911
rect 104932 525855 104988 525911
rect 105056 525855 105112 525911
rect 105180 525855 105236 525911
rect 105304 525855 105360 525911
rect 105428 525855 105484 525911
rect 105552 525855 105608 525911
rect 105676 525855 105732 525911
rect 105800 525855 105856 525911
rect 105924 525855 105980 525911
rect 106048 525855 106104 525911
rect 106172 525855 106228 525911
rect 106296 525855 106352 525911
rect 106420 525855 106476 525911
rect 106544 525855 106600 525911
rect 106668 525855 106724 525911
rect 106792 525855 106848 525911
rect 106916 525855 106972 525911
rect 107040 525855 107096 525911
rect 107164 525855 107220 525911
rect 107288 525855 107344 525911
rect 107412 525855 107468 525911
rect 107536 525855 107592 525911
rect 107660 525855 107716 525911
rect 107784 525855 107840 525911
rect 107908 525855 107964 525911
rect 108032 525855 108088 525911
rect 108156 525855 108212 525911
rect 108280 525855 108336 525911
rect 108404 525855 108460 525911
rect 108528 525855 108584 525911
rect 108652 525855 108708 525911
rect 108776 525855 108832 525911
rect 108900 525855 108956 525911
rect 109024 525855 109080 525911
rect 109148 525855 109204 525911
rect 109272 525855 109328 525911
rect 109396 525855 109452 525911
rect 109520 525855 109576 525911
rect 109644 525855 109700 525911
rect 109768 525855 109824 525911
rect 109892 525855 109948 525911
rect 110016 525855 110072 525911
rect 110140 525855 110196 525911
rect 110264 525855 110320 525911
rect 110388 525855 110444 525911
rect 110512 525855 110568 525911
rect 110636 525855 110692 525911
rect 110760 525855 110816 525911
rect 110884 525855 110940 525911
rect 111008 525855 111064 525911
rect 111132 525855 111188 525911
rect 111256 525855 111312 525911
rect 111380 525855 111436 525911
rect 111504 525855 111560 525911
rect 111628 525855 111684 525911
rect 111752 525855 111808 525911
rect 111876 525855 111932 525911
rect 112000 525855 112056 525911
rect 112124 525855 112180 525911
rect 112248 525855 112304 525911
rect 112372 525855 112428 525911
rect 112496 525855 112552 525911
rect 112620 525855 112676 525911
rect 112744 525855 112800 525911
rect 112868 525855 112924 525911
rect 112992 525855 113048 525911
rect 113116 525855 113172 525911
rect 113240 525855 113296 525911
rect 113364 525855 113420 525911
rect 113488 525855 113544 525911
rect 113612 525855 113668 525911
rect 113736 525855 113792 525911
rect 113860 525855 113916 525911
rect 113984 525855 114040 525911
rect 114108 525855 114164 525911
rect 114232 525855 114288 525911
rect 114356 525855 114412 525911
rect 114480 525855 114536 525911
rect 114604 525855 114660 525911
rect 39954 514294 40010 514350
rect 40078 514294 40134 514350
rect 40202 514294 40258 514350
rect 40326 514294 40382 514350
rect 39954 514170 40010 514226
rect 40078 514170 40134 514226
rect 40202 514170 40258 514226
rect 40326 514170 40382 514226
rect 39954 514046 40010 514102
rect 40078 514046 40134 514102
rect 40202 514046 40258 514102
rect 40326 514046 40382 514102
rect 39954 513922 40010 513978
rect 40078 513922 40134 513978
rect 40202 513922 40258 513978
rect 40326 513922 40382 513978
rect 60202 514356 60258 514412
rect 60326 514356 60382 514412
rect 60450 514356 60506 514412
rect 60202 514232 60258 514288
rect 60326 514232 60382 514288
rect 60450 514232 60506 514288
rect 60202 514108 60258 514164
rect 60326 514108 60382 514164
rect 60450 514108 60506 514164
rect 60202 513984 60258 514040
rect 60326 513984 60382 514040
rect 60450 513984 60506 514040
rect 60202 513860 60258 513916
rect 60326 513860 60382 513916
rect 60450 513860 60506 513916
rect 60574 514356 60630 514412
rect 60698 514356 60754 514412
rect 60822 514356 60878 514412
rect 60946 514356 61002 514412
rect 60574 514232 60630 514288
rect 60698 514232 60754 514288
rect 60822 514232 60878 514288
rect 60946 514232 61002 514288
rect 60574 514108 60630 514164
rect 60698 514108 60754 514164
rect 60822 514108 60878 514164
rect 60946 514108 61002 514164
rect 60574 513984 60630 514040
rect 60698 513984 60754 514040
rect 60822 513984 60878 514040
rect 60946 513984 61002 514040
rect 60574 513860 60630 513916
rect 60698 513860 60754 513916
rect 60822 513860 60878 513916
rect 60946 513860 61002 513916
rect 61070 514356 61126 514412
rect 61194 514356 61250 514412
rect 61318 514356 61374 514412
rect 61442 514356 61498 514412
rect 61070 514232 61126 514288
rect 61194 514232 61250 514288
rect 61318 514232 61374 514288
rect 61442 514232 61498 514288
rect 61070 514108 61126 514164
rect 61194 514108 61250 514164
rect 61318 514108 61374 514164
rect 61442 514108 61498 514164
rect 61070 513984 61126 514040
rect 61194 513984 61250 514040
rect 61318 513984 61374 514040
rect 61442 513984 61498 514040
rect 61070 513860 61126 513916
rect 61194 513860 61250 513916
rect 61318 513860 61374 513916
rect 61442 513860 61498 513916
rect 61566 514356 61622 514412
rect 61690 514356 61746 514412
rect 61814 514356 61870 514412
rect 61938 514356 61994 514412
rect 61566 514232 61622 514288
rect 61690 514232 61746 514288
rect 61814 514232 61870 514288
rect 61938 514232 61994 514288
rect 61566 514108 61622 514164
rect 61690 514108 61746 514164
rect 61814 514108 61870 514164
rect 61938 514108 61994 514164
rect 61566 513984 61622 514040
rect 61690 513984 61746 514040
rect 61814 513984 61870 514040
rect 61938 513984 61994 514040
rect 61566 513860 61622 513916
rect 61690 513860 61746 513916
rect 61814 513860 61870 513916
rect 61938 513860 61994 513916
rect 62062 514356 62118 514412
rect 62186 514356 62242 514412
rect 62310 514356 62366 514412
rect 62434 514356 62490 514412
rect 62062 514232 62118 514288
rect 62186 514232 62242 514288
rect 62310 514232 62366 514288
rect 62434 514232 62490 514288
rect 62062 514108 62118 514164
rect 62186 514108 62242 514164
rect 62310 514108 62366 514164
rect 62434 514108 62490 514164
rect 62062 513984 62118 514040
rect 62186 513984 62242 514040
rect 62310 513984 62366 514040
rect 62434 513984 62490 514040
rect 62062 513860 62118 513916
rect 62186 513860 62242 513916
rect 62310 513860 62366 513916
rect 62434 513860 62490 513916
rect 62558 514356 62614 514412
rect 62682 514356 62738 514412
rect 62806 514356 62862 514412
rect 62930 514356 62986 514412
rect 62558 514232 62614 514288
rect 62682 514232 62738 514288
rect 62806 514232 62862 514288
rect 62930 514232 62986 514288
rect 62558 514108 62614 514164
rect 62682 514108 62738 514164
rect 62806 514108 62862 514164
rect 62930 514108 62986 514164
rect 62558 513984 62614 514040
rect 62682 513984 62738 514040
rect 62806 513984 62862 514040
rect 62930 513984 62986 514040
rect 62558 513860 62614 513916
rect 62682 513860 62738 513916
rect 62806 513860 62862 513916
rect 62930 513860 62986 513916
rect 63054 514356 63110 514412
rect 63178 514356 63234 514412
rect 63302 514356 63358 514412
rect 63426 514356 63482 514412
rect 63054 514232 63110 514288
rect 63178 514232 63234 514288
rect 63302 514232 63358 514288
rect 63426 514232 63482 514288
rect 63054 514108 63110 514164
rect 63178 514108 63234 514164
rect 63302 514108 63358 514164
rect 63426 514108 63482 514164
rect 63054 513984 63110 514040
rect 63178 513984 63234 514040
rect 63302 513984 63358 514040
rect 63426 513984 63482 514040
rect 63054 513860 63110 513916
rect 63178 513860 63234 513916
rect 63302 513860 63358 513916
rect 63426 513860 63482 513916
rect 63550 514356 63606 514412
rect 63674 514356 63730 514412
rect 63798 514356 63854 514412
rect 63922 514356 63978 514412
rect 63550 514232 63606 514288
rect 63674 514232 63730 514288
rect 63798 514232 63854 514288
rect 63922 514232 63978 514288
rect 63550 514108 63606 514164
rect 63674 514108 63730 514164
rect 63798 514108 63854 514164
rect 63922 514108 63978 514164
rect 63550 513984 63606 514040
rect 63674 513984 63730 514040
rect 63798 513984 63854 514040
rect 63922 513984 63978 514040
rect 63550 513860 63606 513916
rect 63674 513860 63730 513916
rect 63798 513860 63854 513916
rect 63922 513860 63978 513916
rect 64046 514356 64102 514412
rect 64170 514356 64226 514412
rect 64294 514356 64350 514412
rect 64418 514356 64474 514412
rect 64046 514232 64102 514288
rect 64170 514232 64226 514288
rect 64294 514232 64350 514288
rect 64418 514232 64474 514288
rect 64046 514108 64102 514164
rect 64170 514108 64226 514164
rect 64294 514108 64350 514164
rect 64418 514108 64474 514164
rect 64046 513984 64102 514040
rect 64170 513984 64226 514040
rect 64294 513984 64350 514040
rect 64418 513984 64474 514040
rect 64046 513860 64102 513916
rect 64170 513860 64226 513916
rect 64294 513860 64350 513916
rect 64418 513860 64474 513916
rect 64542 514356 64598 514412
rect 64666 514356 64722 514412
rect 64790 514356 64846 514412
rect 64914 514356 64970 514412
rect 64542 514232 64598 514288
rect 64666 514232 64722 514288
rect 64790 514232 64846 514288
rect 64914 514232 64970 514288
rect 64542 514108 64598 514164
rect 64666 514108 64722 514164
rect 64790 514108 64846 514164
rect 64914 514108 64970 514164
rect 64542 513984 64598 514040
rect 64666 513984 64722 514040
rect 64790 513984 64846 514040
rect 64914 513984 64970 514040
rect 64542 513860 64598 513916
rect 64666 513860 64722 513916
rect 64790 513860 64846 513916
rect 64914 513860 64970 513916
rect 65038 514356 65094 514412
rect 65162 514356 65218 514412
rect 65286 514356 65342 514412
rect 65410 514356 65466 514412
rect 65038 514232 65094 514288
rect 65162 514232 65218 514288
rect 65286 514232 65342 514288
rect 65410 514232 65466 514288
rect 65038 514108 65094 514164
rect 65162 514108 65218 514164
rect 65286 514108 65342 514164
rect 65410 514108 65466 514164
rect 65038 513984 65094 514040
rect 65162 513984 65218 514040
rect 65286 513984 65342 514040
rect 65410 513984 65466 514040
rect 65038 513860 65094 513916
rect 65162 513860 65218 513916
rect 65286 513860 65342 513916
rect 65410 513860 65466 513916
rect 65534 514356 65590 514412
rect 65658 514356 65714 514412
rect 65782 514356 65838 514412
rect 65906 514356 65962 514412
rect 65534 514232 65590 514288
rect 65658 514232 65714 514288
rect 65782 514232 65838 514288
rect 65906 514232 65962 514288
rect 65534 514108 65590 514164
rect 65658 514108 65714 514164
rect 65782 514108 65838 514164
rect 65906 514108 65962 514164
rect 65534 513984 65590 514040
rect 65658 513984 65714 514040
rect 65782 513984 65838 514040
rect 65906 513984 65962 514040
rect 65534 513860 65590 513916
rect 65658 513860 65714 513916
rect 65782 513860 65838 513916
rect 65906 513860 65962 513916
rect 66030 514356 66086 514412
rect 66154 514356 66210 514412
rect 66278 514356 66334 514412
rect 66402 514356 66458 514412
rect 66030 514232 66086 514288
rect 66154 514232 66210 514288
rect 66278 514232 66334 514288
rect 66402 514232 66458 514288
rect 66030 514108 66086 514164
rect 66154 514108 66210 514164
rect 66278 514108 66334 514164
rect 66402 514108 66458 514164
rect 66030 513984 66086 514040
rect 66154 513984 66210 514040
rect 66278 513984 66334 514040
rect 66402 513984 66458 514040
rect 66030 513860 66086 513916
rect 66154 513860 66210 513916
rect 66278 513860 66334 513916
rect 66402 513860 66458 513916
rect 90112 508379 90168 508435
rect 90236 508379 90292 508435
rect 90360 508379 90416 508435
rect 90484 508379 90540 508435
rect 90608 508379 90664 508435
rect 90732 508379 90788 508435
rect 90856 508379 90912 508435
rect 90980 508379 91036 508435
rect 91104 508379 91160 508435
rect 91228 508379 91284 508435
rect 91352 508379 91408 508435
rect 91476 508379 91532 508435
rect 91600 508379 91656 508435
rect 91724 508379 91780 508435
rect 91848 508379 91904 508435
rect 91972 508379 92028 508435
rect 92096 508379 92152 508435
rect 92220 508379 92276 508435
rect 92344 508379 92400 508435
rect 92468 508379 92524 508435
rect 92592 508379 92648 508435
rect 92716 508379 92772 508435
rect 92840 508379 92896 508435
rect 92964 508379 93020 508435
rect 93088 508379 93144 508435
rect 93212 508379 93268 508435
rect 93336 508379 93392 508435
rect 93460 508379 93516 508435
rect 93584 508379 93640 508435
rect 93708 508379 93764 508435
rect 93832 508379 93888 508435
rect 93956 508379 94012 508435
rect 94080 508379 94136 508435
rect 94204 508379 94260 508435
rect 94328 508379 94384 508435
rect 94452 508379 94508 508435
rect 94576 508379 94632 508435
rect 94700 508379 94756 508435
rect 94824 508379 94880 508435
rect 94948 508379 95004 508435
rect 95072 508379 95128 508435
rect 95196 508379 95252 508435
rect 95320 508379 95376 508435
rect 95444 508379 95500 508435
rect 95568 508379 95624 508435
rect 95692 508379 95748 508435
rect 95816 508379 95872 508435
rect 95940 508379 95996 508435
rect 96064 508379 96120 508435
rect 96188 508379 96244 508435
rect 96312 508379 96368 508435
rect 96436 508379 96492 508435
rect 96560 508379 96616 508435
rect 96684 508379 96740 508435
rect 96808 508379 96864 508435
rect 96932 508379 96988 508435
rect 97056 508379 97112 508435
rect 97180 508379 97236 508435
rect 97304 508379 97360 508435
rect 97428 508379 97484 508435
rect 97552 508379 97608 508435
rect 97676 508379 97732 508435
rect 97800 508379 97856 508435
rect 97924 508379 97980 508435
rect 98048 508379 98104 508435
rect 98172 508379 98228 508435
rect 98296 508379 98352 508435
rect 98420 508379 98476 508435
rect 98544 508379 98600 508435
rect 98668 508379 98724 508435
rect 98792 508379 98848 508435
rect 98916 508379 98972 508435
rect 99040 508379 99096 508435
rect 99164 508379 99220 508435
rect 99288 508379 99344 508435
rect 99412 508379 99468 508435
rect 99536 508379 99592 508435
rect 99660 508379 99716 508435
rect 99784 508379 99840 508435
rect 99908 508379 99964 508435
rect 100032 508379 100088 508435
rect 90112 508255 90168 508311
rect 90236 508255 90292 508311
rect 90360 508255 90416 508311
rect 90484 508255 90540 508311
rect 90608 508255 90664 508311
rect 90732 508255 90788 508311
rect 90856 508255 90912 508311
rect 90980 508255 91036 508311
rect 91104 508255 91160 508311
rect 91228 508255 91284 508311
rect 91352 508255 91408 508311
rect 91476 508255 91532 508311
rect 91600 508255 91656 508311
rect 91724 508255 91780 508311
rect 91848 508255 91904 508311
rect 91972 508255 92028 508311
rect 92096 508255 92152 508311
rect 92220 508255 92276 508311
rect 92344 508255 92400 508311
rect 92468 508255 92524 508311
rect 92592 508255 92648 508311
rect 92716 508255 92772 508311
rect 92840 508255 92896 508311
rect 92964 508255 93020 508311
rect 93088 508255 93144 508311
rect 93212 508255 93268 508311
rect 93336 508255 93392 508311
rect 93460 508255 93516 508311
rect 93584 508255 93640 508311
rect 93708 508255 93764 508311
rect 93832 508255 93888 508311
rect 93956 508255 94012 508311
rect 94080 508255 94136 508311
rect 94204 508255 94260 508311
rect 94328 508255 94384 508311
rect 94452 508255 94508 508311
rect 94576 508255 94632 508311
rect 94700 508255 94756 508311
rect 94824 508255 94880 508311
rect 94948 508255 95004 508311
rect 95072 508255 95128 508311
rect 95196 508255 95252 508311
rect 95320 508255 95376 508311
rect 95444 508255 95500 508311
rect 95568 508255 95624 508311
rect 95692 508255 95748 508311
rect 95816 508255 95872 508311
rect 95940 508255 95996 508311
rect 96064 508255 96120 508311
rect 96188 508255 96244 508311
rect 96312 508255 96368 508311
rect 96436 508255 96492 508311
rect 96560 508255 96616 508311
rect 96684 508255 96740 508311
rect 96808 508255 96864 508311
rect 96932 508255 96988 508311
rect 97056 508255 97112 508311
rect 97180 508255 97236 508311
rect 97304 508255 97360 508311
rect 97428 508255 97484 508311
rect 97552 508255 97608 508311
rect 97676 508255 97732 508311
rect 97800 508255 97856 508311
rect 97924 508255 97980 508311
rect 98048 508255 98104 508311
rect 98172 508255 98228 508311
rect 98296 508255 98352 508311
rect 98420 508255 98476 508311
rect 98544 508255 98600 508311
rect 98668 508255 98724 508311
rect 98792 508255 98848 508311
rect 98916 508255 98972 508311
rect 99040 508255 99096 508311
rect 99164 508255 99220 508311
rect 99288 508255 99344 508311
rect 99412 508255 99468 508311
rect 99536 508255 99592 508311
rect 99660 508255 99716 508311
rect 99784 508255 99840 508311
rect 99908 508255 99964 508311
rect 100032 508255 100088 508311
rect 90112 508131 90168 508187
rect 90236 508131 90292 508187
rect 90360 508131 90416 508187
rect 90484 508131 90540 508187
rect 90608 508131 90664 508187
rect 90732 508131 90788 508187
rect 90856 508131 90912 508187
rect 90980 508131 91036 508187
rect 91104 508131 91160 508187
rect 91228 508131 91284 508187
rect 91352 508131 91408 508187
rect 91476 508131 91532 508187
rect 91600 508131 91656 508187
rect 91724 508131 91780 508187
rect 91848 508131 91904 508187
rect 91972 508131 92028 508187
rect 92096 508131 92152 508187
rect 92220 508131 92276 508187
rect 92344 508131 92400 508187
rect 92468 508131 92524 508187
rect 92592 508131 92648 508187
rect 92716 508131 92772 508187
rect 92840 508131 92896 508187
rect 92964 508131 93020 508187
rect 93088 508131 93144 508187
rect 93212 508131 93268 508187
rect 93336 508131 93392 508187
rect 93460 508131 93516 508187
rect 93584 508131 93640 508187
rect 93708 508131 93764 508187
rect 93832 508131 93888 508187
rect 93956 508131 94012 508187
rect 94080 508131 94136 508187
rect 94204 508131 94260 508187
rect 94328 508131 94384 508187
rect 94452 508131 94508 508187
rect 94576 508131 94632 508187
rect 94700 508131 94756 508187
rect 94824 508131 94880 508187
rect 94948 508131 95004 508187
rect 95072 508131 95128 508187
rect 95196 508131 95252 508187
rect 95320 508131 95376 508187
rect 95444 508131 95500 508187
rect 95568 508131 95624 508187
rect 95692 508131 95748 508187
rect 95816 508131 95872 508187
rect 95940 508131 95996 508187
rect 96064 508131 96120 508187
rect 96188 508131 96244 508187
rect 96312 508131 96368 508187
rect 96436 508131 96492 508187
rect 96560 508131 96616 508187
rect 96684 508131 96740 508187
rect 96808 508131 96864 508187
rect 96932 508131 96988 508187
rect 97056 508131 97112 508187
rect 97180 508131 97236 508187
rect 97304 508131 97360 508187
rect 97428 508131 97484 508187
rect 97552 508131 97608 508187
rect 97676 508131 97732 508187
rect 97800 508131 97856 508187
rect 97924 508131 97980 508187
rect 98048 508131 98104 508187
rect 98172 508131 98228 508187
rect 98296 508131 98352 508187
rect 98420 508131 98476 508187
rect 98544 508131 98600 508187
rect 98668 508131 98724 508187
rect 98792 508131 98848 508187
rect 98916 508131 98972 508187
rect 99040 508131 99096 508187
rect 99164 508131 99220 508187
rect 99288 508131 99344 508187
rect 99412 508131 99468 508187
rect 99536 508131 99592 508187
rect 99660 508131 99716 508187
rect 99784 508131 99840 508187
rect 99908 508131 99964 508187
rect 100032 508131 100088 508187
rect 39954 496294 40010 496350
rect 40078 496294 40134 496350
rect 40202 496294 40258 496350
rect 40326 496294 40382 496350
rect 39954 496170 40010 496226
rect 40078 496170 40134 496226
rect 40202 496170 40258 496226
rect 40326 496170 40382 496226
rect 39954 496046 40010 496102
rect 40078 496046 40134 496102
rect 40202 496046 40258 496102
rect 40326 496046 40382 496102
rect 39954 495922 40010 495978
rect 40078 495922 40134 495978
rect 40202 495922 40258 495978
rect 40326 495922 40382 495978
rect 63430 496156 63486 496212
rect 63430 496032 63486 496088
rect 63430 495908 63486 495964
rect 63554 496156 63610 496212
rect 63678 496156 63734 496212
rect 63802 496156 63858 496212
rect 63926 496156 63982 496212
rect 63554 496032 63610 496088
rect 63678 496032 63734 496088
rect 63802 496032 63858 496088
rect 63926 496032 63982 496088
rect 63554 495908 63610 495964
rect 63678 495908 63734 495964
rect 63802 495908 63858 495964
rect 63926 495908 63982 495964
rect 64050 496156 64106 496212
rect 64174 496156 64230 496212
rect 64298 496156 64354 496212
rect 64422 496156 64478 496212
rect 64050 496032 64106 496088
rect 64174 496032 64230 496088
rect 64298 496032 64354 496088
rect 64422 496032 64478 496088
rect 64050 495908 64106 495964
rect 64174 495908 64230 495964
rect 64298 495908 64354 495964
rect 64422 495908 64478 495964
rect 64546 496156 64602 496212
rect 64670 496156 64726 496212
rect 64794 496156 64850 496212
rect 64918 496156 64974 496212
rect 64546 496032 64602 496088
rect 64670 496032 64726 496088
rect 64794 496032 64850 496088
rect 64918 496032 64974 496088
rect 64546 495908 64602 495964
rect 64670 495908 64726 495964
rect 64794 495908 64850 495964
rect 64918 495908 64974 495964
rect 65042 496156 65098 496212
rect 65166 496156 65222 496212
rect 65290 496156 65346 496212
rect 65414 496156 65470 496212
rect 65042 496032 65098 496088
rect 65166 496032 65222 496088
rect 65290 496032 65346 496088
rect 65414 496032 65470 496088
rect 65042 495908 65098 495964
rect 65166 495908 65222 495964
rect 65290 495908 65346 495964
rect 65414 495908 65470 495964
rect 65538 496156 65594 496212
rect 65662 496156 65718 496212
rect 65786 496156 65842 496212
rect 65910 496156 65966 496212
rect 65538 496032 65594 496088
rect 65662 496032 65718 496088
rect 65786 496032 65842 496088
rect 65910 496032 65966 496088
rect 65538 495908 65594 495964
rect 65662 495908 65718 495964
rect 65786 495908 65842 495964
rect 65910 495908 65966 495964
rect 66034 496156 66090 496212
rect 66158 496156 66214 496212
rect 66282 496156 66338 496212
rect 66406 496156 66462 496212
rect 66034 496032 66090 496088
rect 66158 496032 66214 496088
rect 66282 496032 66338 496088
rect 66406 496032 66462 496088
rect 66034 495908 66090 495964
rect 66158 495908 66214 495964
rect 66282 495908 66338 495964
rect 66406 495908 66462 495964
rect 66530 496156 66586 496212
rect 66654 496156 66710 496212
rect 66778 496156 66834 496212
rect 66902 496156 66958 496212
rect 66530 496032 66586 496088
rect 66654 496032 66710 496088
rect 66778 496032 66834 496088
rect 66902 496032 66958 496088
rect 66530 495908 66586 495964
rect 66654 495908 66710 495964
rect 66778 495908 66834 495964
rect 66902 495908 66958 495964
rect 67026 496156 67082 496212
rect 67150 496156 67206 496212
rect 67274 496156 67330 496212
rect 67398 496156 67454 496212
rect 67026 496032 67082 496088
rect 67150 496032 67206 496088
rect 67274 496032 67330 496088
rect 67398 496032 67454 496088
rect 67026 495908 67082 495964
rect 67150 495908 67206 495964
rect 67274 495908 67330 495964
rect 67398 495908 67454 495964
rect 67522 496156 67578 496212
rect 67646 496156 67702 496212
rect 67770 496156 67826 496212
rect 67894 496156 67950 496212
rect 67522 496032 67578 496088
rect 67646 496032 67702 496088
rect 67770 496032 67826 496088
rect 67894 496032 67950 496088
rect 67522 495908 67578 495964
rect 67646 495908 67702 495964
rect 67770 495908 67826 495964
rect 67894 495908 67950 495964
rect 68018 496156 68074 496212
rect 68142 496156 68198 496212
rect 68266 496156 68322 496212
rect 68390 496156 68446 496212
rect 68018 496032 68074 496088
rect 68142 496032 68198 496088
rect 68266 496032 68322 496088
rect 68390 496032 68446 496088
rect 68018 495908 68074 495964
rect 68142 495908 68198 495964
rect 68266 495908 68322 495964
rect 68390 495908 68446 495964
rect 68514 496156 68570 496212
rect 68638 496156 68694 496212
rect 68762 496156 68818 496212
rect 68886 496156 68942 496212
rect 68514 496032 68570 496088
rect 68638 496032 68694 496088
rect 68762 496032 68818 496088
rect 68886 496032 68942 496088
rect 68514 495908 68570 495964
rect 68638 495908 68694 495964
rect 68762 495908 68818 495964
rect 68886 495908 68942 495964
rect 69010 496156 69066 496212
rect 69134 496156 69190 496212
rect 69258 496156 69314 496212
rect 69382 496156 69438 496212
rect 69010 496032 69066 496088
rect 69134 496032 69190 496088
rect 69258 496032 69314 496088
rect 69382 496032 69438 496088
rect 69010 495908 69066 495964
rect 69134 495908 69190 495964
rect 69258 495908 69314 495964
rect 69382 495908 69438 495964
rect 69506 496156 69562 496212
rect 69630 496156 69686 496212
rect 69754 496156 69810 496212
rect 69878 496156 69934 496212
rect 69506 496032 69562 496088
rect 69630 496032 69686 496088
rect 69754 496032 69810 496088
rect 69878 496032 69934 496088
rect 69506 495908 69562 495964
rect 69630 495908 69686 495964
rect 69754 495908 69810 495964
rect 69878 495908 69934 495964
rect 70002 496156 70058 496212
rect 70126 496156 70182 496212
rect 70250 496156 70306 496212
rect 70374 496156 70430 496212
rect 70002 496032 70058 496088
rect 70126 496032 70182 496088
rect 70250 496032 70306 496088
rect 70374 496032 70430 496088
rect 70002 495908 70058 495964
rect 70126 495908 70182 495964
rect 70250 495908 70306 495964
rect 70374 495908 70430 495964
rect 85236 490216 85292 490272
rect 85360 490216 85416 490272
rect 85484 490216 85540 490272
rect 85608 490216 85664 490272
rect 85732 490216 85788 490272
rect 85856 490216 85912 490272
rect 85980 490216 86036 490272
rect 86104 490216 86160 490272
rect 86228 490216 86284 490272
rect 86352 490216 86408 490272
rect 86476 490216 86532 490272
rect 86600 490216 86656 490272
rect 86724 490216 86780 490272
rect 86848 490216 86904 490272
rect 86972 490216 87028 490272
rect 87096 490216 87152 490272
rect 87220 490216 87276 490272
rect 87344 490216 87400 490272
rect 87468 490216 87524 490272
rect 87592 490216 87648 490272
rect 87716 490216 87772 490272
rect 87840 490216 87896 490272
rect 87964 490216 88020 490272
rect 88088 490216 88144 490272
rect 88212 490216 88268 490272
rect 88336 490216 88392 490272
rect 88460 490216 88516 490272
rect 88584 490216 88640 490272
rect 88708 490216 88764 490272
rect 85236 490092 85292 490148
rect 85360 490092 85416 490148
rect 85484 490092 85540 490148
rect 85608 490092 85664 490148
rect 85732 490092 85788 490148
rect 85856 490092 85912 490148
rect 85980 490092 86036 490148
rect 86104 490092 86160 490148
rect 86228 490092 86284 490148
rect 86352 490092 86408 490148
rect 86476 490092 86532 490148
rect 86600 490092 86656 490148
rect 86724 490092 86780 490148
rect 86848 490092 86904 490148
rect 86972 490092 87028 490148
rect 87096 490092 87152 490148
rect 87220 490092 87276 490148
rect 87344 490092 87400 490148
rect 87468 490092 87524 490148
rect 87592 490092 87648 490148
rect 87716 490092 87772 490148
rect 87840 490092 87896 490148
rect 87964 490092 88020 490148
rect 88088 490092 88144 490148
rect 88212 490092 88268 490148
rect 88336 490092 88392 490148
rect 88460 490092 88516 490148
rect 88584 490092 88640 490148
rect 88708 490092 88764 490148
rect 85236 489968 85292 490024
rect 85360 489968 85416 490024
rect 85484 489968 85540 490024
rect 85608 489968 85664 490024
rect 85732 489968 85788 490024
rect 85856 489968 85912 490024
rect 85980 489968 86036 490024
rect 86104 489968 86160 490024
rect 86228 489968 86284 490024
rect 86352 489968 86408 490024
rect 86476 489968 86532 490024
rect 86600 489968 86656 490024
rect 86724 489968 86780 490024
rect 86848 489968 86904 490024
rect 86972 489968 87028 490024
rect 87096 489968 87152 490024
rect 87220 489968 87276 490024
rect 87344 489968 87400 490024
rect 87468 489968 87524 490024
rect 87592 489968 87648 490024
rect 87716 489968 87772 490024
rect 87840 489968 87896 490024
rect 87964 489968 88020 490024
rect 88088 489968 88144 490024
rect 88212 489968 88268 490024
rect 88336 489968 88392 490024
rect 88460 489968 88516 490024
rect 88584 489968 88640 490024
rect 88708 489968 88764 490024
rect 39954 478294 40010 478350
rect 40078 478294 40134 478350
rect 40202 478294 40258 478350
rect 40326 478294 40382 478350
rect 39954 478170 40010 478226
rect 40078 478170 40134 478226
rect 40202 478170 40258 478226
rect 40326 478170 40382 478226
rect 39954 478046 40010 478102
rect 40078 478046 40134 478102
rect 40202 478046 40258 478102
rect 40326 478046 40382 478102
rect 39954 477922 40010 477978
rect 40078 477922 40134 477978
rect 40202 477922 40258 477978
rect 40326 477922 40382 477978
rect 39954 460294 40010 460350
rect 40078 460294 40134 460350
rect 40202 460294 40258 460350
rect 40326 460294 40382 460350
rect 39954 460170 40010 460226
rect 40078 460170 40134 460226
rect 40202 460170 40258 460226
rect 40326 460170 40382 460226
rect 39954 460046 40010 460102
rect 40078 460046 40134 460102
rect 40202 460046 40258 460102
rect 40326 460046 40382 460102
rect 39954 459922 40010 459978
rect 40078 459922 40134 459978
rect 40202 459922 40258 459978
rect 40326 459922 40382 459978
rect 39954 442294 40010 442350
rect 40078 442294 40134 442350
rect 40202 442294 40258 442350
rect 40326 442294 40382 442350
rect 39954 442170 40010 442226
rect 40078 442170 40134 442226
rect 40202 442170 40258 442226
rect 40326 442170 40382 442226
rect 39954 442046 40010 442102
rect 40078 442046 40134 442102
rect 40202 442046 40258 442102
rect 40326 442046 40382 442102
rect 39954 441922 40010 441978
rect 40078 441922 40134 441978
rect 40202 441922 40258 441978
rect 40326 441922 40382 441978
rect 39954 424294 40010 424350
rect 40078 424294 40134 424350
rect 40202 424294 40258 424350
rect 40326 424294 40382 424350
rect 39954 424170 40010 424226
rect 40078 424170 40134 424226
rect 40202 424170 40258 424226
rect 40326 424170 40382 424226
rect 39954 424046 40010 424102
rect 40078 424046 40134 424102
rect 40202 424046 40258 424102
rect 40326 424046 40382 424102
rect 39954 423922 40010 423978
rect 40078 423922 40134 423978
rect 40202 423922 40258 423978
rect 40326 423922 40382 423978
rect 66954 472294 67010 472350
rect 67078 472294 67134 472350
rect 67202 472294 67258 472350
rect 67326 472294 67382 472350
rect 66954 472170 67010 472226
rect 67078 472170 67134 472226
rect 67202 472170 67258 472226
rect 67326 472170 67382 472226
rect 66954 472046 67010 472102
rect 67078 472046 67134 472102
rect 67202 472046 67258 472102
rect 67326 472046 67382 472102
rect 66954 471922 67010 471978
rect 67078 471922 67134 471978
rect 67202 471922 67258 471978
rect 67326 471922 67382 471978
rect 66954 454294 67010 454350
rect 67078 454294 67134 454350
rect 67202 454294 67258 454350
rect 67326 454294 67382 454350
rect 66954 454170 67010 454226
rect 67078 454170 67134 454226
rect 67202 454170 67258 454226
rect 67326 454170 67382 454226
rect 66954 454046 67010 454102
rect 67078 454046 67134 454102
rect 67202 454046 67258 454102
rect 67326 454046 67382 454102
rect 66954 453922 67010 453978
rect 67078 453922 67134 453978
rect 67202 453922 67258 453978
rect 67326 453922 67382 453978
rect 66954 436294 67010 436350
rect 67078 436294 67134 436350
rect 67202 436294 67258 436350
rect 67326 436294 67382 436350
rect 66954 436170 67010 436226
rect 67078 436170 67134 436226
rect 67202 436170 67258 436226
rect 67326 436170 67382 436226
rect 66954 436046 67010 436102
rect 67078 436046 67134 436102
rect 67202 436046 67258 436102
rect 67326 436046 67382 436102
rect 66954 435922 67010 435978
rect 67078 435922 67134 435978
rect 67202 435922 67258 435978
rect 67326 435922 67382 435978
rect 66954 418294 67010 418350
rect 67078 418294 67134 418350
rect 67202 418294 67258 418350
rect 67326 418294 67382 418350
rect 66954 418170 67010 418226
rect 67078 418170 67134 418226
rect 67202 418170 67258 418226
rect 67326 418170 67382 418226
rect 66954 418046 67010 418102
rect 67078 418046 67134 418102
rect 67202 418046 67258 418102
rect 67326 418046 67382 418102
rect 66954 417922 67010 417978
rect 67078 417922 67134 417978
rect 67202 417922 67258 417978
rect 67326 417922 67382 417978
rect 70674 478294 70730 478350
rect 70798 478294 70854 478350
rect 70922 478294 70978 478350
rect 71046 478294 71102 478350
rect 80936 478302 80992 478358
rect 81060 478302 81116 478358
rect 81184 478302 81240 478358
rect 81308 478302 81364 478358
rect 70674 478170 70730 478226
rect 70798 478170 70854 478226
rect 70922 478170 70978 478226
rect 71046 478170 71102 478226
rect 70674 478046 70730 478102
rect 70798 478046 70854 478102
rect 70922 478046 70978 478102
rect 71046 478046 71102 478102
rect 70674 477922 70730 477978
rect 70798 477922 70854 477978
rect 70922 477922 70978 477978
rect 71046 477922 71102 477978
rect 70674 460294 70730 460350
rect 70798 460294 70854 460350
rect 70922 460294 70978 460350
rect 71046 460294 71102 460350
rect 70674 460170 70730 460226
rect 70798 460170 70854 460226
rect 70922 460170 70978 460226
rect 71046 460170 71102 460226
rect 70674 460046 70730 460102
rect 70798 460046 70854 460102
rect 70922 460046 70978 460102
rect 71046 460046 71102 460102
rect 70674 459922 70730 459978
rect 70798 459922 70854 459978
rect 70922 459922 70978 459978
rect 71046 459922 71102 459978
rect 70674 442294 70730 442350
rect 70798 442294 70854 442350
rect 70922 442294 70978 442350
rect 71046 442294 71102 442350
rect 70674 442170 70730 442226
rect 70798 442170 70854 442226
rect 70922 442170 70978 442226
rect 71046 442170 71102 442226
rect 70674 442046 70730 442102
rect 70798 442046 70854 442102
rect 70922 442046 70978 442102
rect 71046 442046 71102 442102
rect 70674 441922 70730 441978
rect 70798 441922 70854 441978
rect 70922 441922 70978 441978
rect 71046 441922 71102 441978
rect 70674 424294 70730 424350
rect 70798 424294 70854 424350
rect 70922 424294 70978 424350
rect 71046 424294 71102 424350
rect 70674 424170 70730 424226
rect 70798 424170 70854 424226
rect 70922 424170 70978 424226
rect 71046 424170 71102 424226
rect 70674 424046 70730 424102
rect 70798 424046 70854 424102
rect 70922 424046 70978 424102
rect 71046 424046 71102 424102
rect 70674 423922 70730 423978
rect 70798 423922 70854 423978
rect 70922 423922 70978 423978
rect 71046 423922 71102 423978
rect 97674 472294 97730 472350
rect 97798 472294 97854 472350
rect 97922 472294 97978 472350
rect 98046 472294 98102 472350
rect 97674 472170 97730 472226
rect 97798 472170 97854 472226
rect 97922 472170 97978 472226
rect 98046 472170 98102 472226
rect 97674 472046 97730 472102
rect 97798 472046 97854 472102
rect 97922 472046 97978 472102
rect 98046 472046 98102 472102
rect 97674 471922 97730 471978
rect 97798 471922 97854 471978
rect 97922 471922 97978 471978
rect 98046 471922 98102 471978
rect 97674 454294 97730 454350
rect 97798 454294 97854 454350
rect 97922 454294 97978 454350
rect 98046 454294 98102 454350
rect 97674 454170 97730 454226
rect 97798 454170 97854 454226
rect 97922 454170 97978 454226
rect 98046 454170 98102 454226
rect 97674 454046 97730 454102
rect 97798 454046 97854 454102
rect 97922 454046 97978 454102
rect 98046 454046 98102 454102
rect 97674 453922 97730 453978
rect 97798 453922 97854 453978
rect 97922 453922 97978 453978
rect 98046 453922 98102 453978
rect 97674 436294 97730 436350
rect 97798 436294 97854 436350
rect 97922 436294 97978 436350
rect 98046 436294 98102 436350
rect 97674 436170 97730 436226
rect 97798 436170 97854 436226
rect 97922 436170 97978 436226
rect 98046 436170 98102 436226
rect 97674 436046 97730 436102
rect 97798 436046 97854 436102
rect 97922 436046 97978 436102
rect 98046 436046 98102 436102
rect 97674 435922 97730 435978
rect 97798 435922 97854 435978
rect 97922 435922 97978 435978
rect 98046 435922 98102 435978
rect 97674 418294 97730 418350
rect 97798 418294 97854 418350
rect 97922 418294 97978 418350
rect 98046 418294 98102 418350
rect 97674 418170 97730 418226
rect 97798 418170 97854 418226
rect 97922 418170 97978 418226
rect 98046 418170 98102 418226
rect 97674 418046 97730 418102
rect 97798 418046 97854 418102
rect 97922 418046 97978 418102
rect 98046 418046 98102 418102
rect 97674 417922 97730 417978
rect 97798 417922 97854 417978
rect 97922 417922 97978 417978
rect 98046 417922 98102 417978
rect 83916 416762 83972 416818
rect 39954 406294 40010 406350
rect 40078 406294 40134 406350
rect 40202 406294 40258 406350
rect 40326 406294 40382 406350
rect 39954 406170 40010 406226
rect 40078 406170 40134 406226
rect 40202 406170 40258 406226
rect 40326 406170 40382 406226
rect 39954 406046 40010 406102
rect 40078 406046 40134 406102
rect 40202 406046 40258 406102
rect 40326 406046 40382 406102
rect 39954 405922 40010 405978
rect 40078 405922 40134 405978
rect 40202 405922 40258 405978
rect 40326 405922 40382 405978
rect 66574 406294 66630 406350
rect 66698 406294 66754 406350
rect 66574 406170 66630 406226
rect 66698 406170 66754 406226
rect 66574 406046 66630 406102
rect 66698 406046 66754 406102
rect 66574 405922 66630 405978
rect 66698 405922 66754 405978
rect 71894 406294 71950 406350
rect 72018 406294 72074 406350
rect 71894 406170 71950 406226
rect 72018 406170 72074 406226
rect 71894 406046 71950 406102
rect 72018 406046 72074 406102
rect 71894 405922 71950 405978
rect 72018 405922 72074 405978
rect 77214 406294 77270 406350
rect 77338 406294 77394 406350
rect 77214 406170 77270 406226
rect 77338 406170 77394 406226
rect 77214 406046 77270 406102
rect 77338 406046 77394 406102
rect 77214 405922 77270 405978
rect 77338 405922 77394 405978
rect 82534 406294 82590 406350
rect 82658 406294 82714 406350
rect 82534 406170 82590 406226
rect 82658 406170 82714 406226
rect 82534 406046 82590 406102
rect 82658 406046 82714 406102
rect 82534 405922 82590 405978
rect 82658 405922 82714 405978
rect 63914 400294 63970 400350
rect 64038 400294 64094 400350
rect 63914 400170 63970 400226
rect 64038 400170 64094 400226
rect 63914 400046 63970 400102
rect 64038 400046 64094 400102
rect 63914 399922 63970 399978
rect 64038 399922 64094 399978
rect 69234 400294 69290 400350
rect 69358 400294 69414 400350
rect 69234 400170 69290 400226
rect 69358 400170 69414 400226
rect 69234 400046 69290 400102
rect 69358 400046 69414 400102
rect 69234 399922 69290 399978
rect 69358 399922 69414 399978
rect 74554 400294 74610 400350
rect 74678 400294 74734 400350
rect 74554 400170 74610 400226
rect 74678 400170 74734 400226
rect 74554 400046 74610 400102
rect 74678 400046 74734 400102
rect 74554 399922 74610 399978
rect 74678 399922 74734 399978
rect 79874 400294 79930 400350
rect 79998 400294 80054 400350
rect 79874 400170 79930 400226
rect 79998 400170 80054 400226
rect 79874 400046 79930 400102
rect 79998 400046 80054 400102
rect 79874 399922 79930 399978
rect 79998 399922 80054 399978
rect 62076 390482 62132 390538
rect 39954 388294 40010 388350
rect 40078 388294 40134 388350
rect 40202 388294 40258 388350
rect 40326 388294 40382 388350
rect 39954 388170 40010 388226
rect 40078 388170 40134 388226
rect 40202 388170 40258 388226
rect 40326 388170 40382 388226
rect 39954 388046 40010 388102
rect 40078 388046 40134 388102
rect 40202 388046 40258 388102
rect 40326 388046 40382 388102
rect 39954 387922 40010 387978
rect 40078 387922 40134 387978
rect 40202 387922 40258 387978
rect 40326 387922 40382 387978
rect 36234 364294 36290 364350
rect 36358 364294 36414 364350
rect 36482 364294 36538 364350
rect 36606 364294 36662 364350
rect 36234 364170 36290 364226
rect 36358 364170 36414 364226
rect 36482 364170 36538 364226
rect 36606 364170 36662 364226
rect 36234 364046 36290 364102
rect 36358 364046 36414 364102
rect 36482 364046 36538 364102
rect 36606 364046 36662 364102
rect 36234 363922 36290 363978
rect 36358 363922 36414 363978
rect 36482 363922 36538 363978
rect 36606 363922 36662 363978
rect 36234 346294 36290 346350
rect 36358 346294 36414 346350
rect 36482 346294 36538 346350
rect 36606 346294 36662 346350
rect 36234 346170 36290 346226
rect 36358 346170 36414 346226
rect 36482 346170 36538 346226
rect 36606 346170 36662 346226
rect 36234 346046 36290 346102
rect 36358 346046 36414 346102
rect 36482 346046 36538 346102
rect 36606 346046 36662 346102
rect 36234 345922 36290 345978
rect 36358 345922 36414 345978
rect 36482 345922 36538 345978
rect 36606 345922 36662 345978
rect 36234 328294 36290 328350
rect 36358 328294 36414 328350
rect 36482 328294 36538 328350
rect 36606 328294 36662 328350
rect 36234 328170 36290 328226
rect 36358 328170 36414 328226
rect 36482 328170 36538 328226
rect 36606 328170 36662 328226
rect 36234 328046 36290 328102
rect 36358 328046 36414 328102
rect 36482 328046 36538 328102
rect 36606 328046 36662 328102
rect 36234 327922 36290 327978
rect 36358 327922 36414 327978
rect 36482 327922 36538 327978
rect 36606 327922 36662 327978
rect 36234 310294 36290 310350
rect 36358 310294 36414 310350
rect 36482 310294 36538 310350
rect 36606 310294 36662 310350
rect 36234 310170 36290 310226
rect 36358 310170 36414 310226
rect 36482 310170 36538 310226
rect 36606 310170 36662 310226
rect 36234 310046 36290 310102
rect 36358 310046 36414 310102
rect 36482 310046 36538 310102
rect 36606 310046 36662 310102
rect 36234 309922 36290 309978
rect 36358 309922 36414 309978
rect 36482 309922 36538 309978
rect 36606 309922 36662 309978
rect 36234 292294 36290 292350
rect 36358 292294 36414 292350
rect 36482 292294 36538 292350
rect 36606 292294 36662 292350
rect 36234 292170 36290 292226
rect 36358 292170 36414 292226
rect 36482 292170 36538 292226
rect 36606 292170 36662 292226
rect 36234 292046 36290 292102
rect 36358 292046 36414 292102
rect 36482 292046 36538 292102
rect 36606 292046 36662 292102
rect 36234 291922 36290 291978
rect 36358 291922 36414 291978
rect 36482 291922 36538 291978
rect 36606 291922 36662 291978
rect 36234 274294 36290 274350
rect 36358 274294 36414 274350
rect 36482 274294 36538 274350
rect 36606 274294 36662 274350
rect 36234 274170 36290 274226
rect 36358 274170 36414 274226
rect 36482 274170 36538 274226
rect 36606 274170 36662 274226
rect 36234 274046 36290 274102
rect 36358 274046 36414 274102
rect 36482 274046 36538 274102
rect 36606 274046 36662 274102
rect 36234 273922 36290 273978
rect 36358 273922 36414 273978
rect 36482 273922 36538 273978
rect 36606 273922 36662 273978
rect 36234 256294 36290 256350
rect 36358 256294 36414 256350
rect 36482 256294 36538 256350
rect 36606 256294 36662 256350
rect 36234 256170 36290 256226
rect 36358 256170 36414 256226
rect 36482 256170 36538 256226
rect 36606 256170 36662 256226
rect 36234 256046 36290 256102
rect 36358 256046 36414 256102
rect 36482 256046 36538 256102
rect 36606 256046 36662 256102
rect 36234 255922 36290 255978
rect 36358 255922 36414 255978
rect 36482 255922 36538 255978
rect 36606 255922 36662 255978
rect 36234 238294 36290 238350
rect 36358 238294 36414 238350
rect 36482 238294 36538 238350
rect 36606 238294 36662 238350
rect 36234 238170 36290 238226
rect 36358 238170 36414 238226
rect 36482 238170 36538 238226
rect 36606 238170 36662 238226
rect 36234 238046 36290 238102
rect 36358 238046 36414 238102
rect 36482 238046 36538 238102
rect 36606 238046 36662 238102
rect 36234 237922 36290 237978
rect 36358 237922 36414 237978
rect 36482 237922 36538 237978
rect 36606 237922 36662 237978
rect 33404 224162 33460 224218
rect 39676 373742 39732 373798
rect 39954 370294 40010 370350
rect 40078 370294 40134 370350
rect 40202 370294 40258 370350
rect 40326 370294 40382 370350
rect 39954 370170 40010 370226
rect 40078 370170 40134 370226
rect 40202 370170 40258 370226
rect 40326 370170 40382 370226
rect 39954 370046 40010 370102
rect 40078 370046 40134 370102
rect 40202 370046 40258 370102
rect 40326 370046 40382 370102
rect 39954 369922 40010 369978
rect 40078 369922 40134 369978
rect 40202 369922 40258 369978
rect 40326 369922 40382 369978
rect 66954 382294 67010 382350
rect 67078 382294 67134 382350
rect 67202 382294 67258 382350
rect 67326 382294 67382 382350
rect 66954 382170 67010 382226
rect 67078 382170 67134 382226
rect 67202 382170 67258 382226
rect 67326 382170 67382 382226
rect 66954 382046 67010 382102
rect 67078 382046 67134 382102
rect 67202 382046 67258 382102
rect 67326 382046 67382 382102
rect 66954 381922 67010 381978
rect 67078 381922 67134 381978
rect 67202 381922 67258 381978
rect 67326 381922 67382 381978
rect 66954 364294 67010 364350
rect 67078 364294 67134 364350
rect 67202 364294 67258 364350
rect 67326 364294 67382 364350
rect 66954 364170 67010 364226
rect 67078 364170 67134 364226
rect 67202 364170 67258 364226
rect 67326 364170 67382 364226
rect 66954 364046 67010 364102
rect 67078 364046 67134 364102
rect 67202 364046 67258 364102
rect 67326 364046 67382 364102
rect 66954 363922 67010 363978
rect 67078 363922 67134 363978
rect 67202 363922 67258 363978
rect 67326 363922 67382 363978
rect 70674 388294 70730 388350
rect 70798 388294 70854 388350
rect 70922 388294 70978 388350
rect 71046 388294 71102 388350
rect 70674 388170 70730 388226
rect 70798 388170 70854 388226
rect 70922 388170 70978 388226
rect 71046 388170 71102 388226
rect 70674 388046 70730 388102
rect 70798 388046 70854 388102
rect 70922 388046 70978 388102
rect 71046 388046 71102 388102
rect 70674 387922 70730 387978
rect 70798 387922 70854 387978
rect 70922 387922 70978 387978
rect 71046 387922 71102 387978
rect 70674 370294 70730 370350
rect 70798 370294 70854 370350
rect 70922 370294 70978 370350
rect 71046 370294 71102 370350
rect 70674 370170 70730 370226
rect 70798 370170 70854 370226
rect 70922 370170 70978 370226
rect 71046 370170 71102 370226
rect 70674 370046 70730 370102
rect 70798 370046 70854 370102
rect 70922 370046 70978 370102
rect 71046 370046 71102 370102
rect 70674 369922 70730 369978
rect 70798 369922 70854 369978
rect 70922 369922 70978 369978
rect 71046 369922 71102 369978
rect 86492 356102 86548 356158
rect 89852 354302 89908 354358
rect 39954 352294 40010 352350
rect 40078 352294 40134 352350
rect 40202 352294 40258 352350
rect 40326 352294 40382 352350
rect 39954 352170 40010 352226
rect 40078 352170 40134 352226
rect 40202 352170 40258 352226
rect 40326 352170 40382 352226
rect 39954 352046 40010 352102
rect 40078 352046 40134 352102
rect 40202 352046 40258 352102
rect 40326 352046 40382 352102
rect 39954 351922 40010 351978
rect 40078 351922 40134 351978
rect 40202 351922 40258 351978
rect 40326 351922 40382 351978
rect 69878 352294 69934 352350
rect 70002 352294 70058 352350
rect 69878 352170 69934 352226
rect 70002 352170 70058 352226
rect 69878 352046 69934 352102
rect 70002 352046 70058 352102
rect 69878 351922 69934 351978
rect 70002 351922 70058 351978
rect 54518 346294 54574 346350
rect 54642 346294 54698 346350
rect 54518 346170 54574 346226
rect 54642 346170 54698 346226
rect 54518 346046 54574 346102
rect 54642 346046 54698 346102
rect 54518 345922 54574 345978
rect 54642 345922 54698 345978
rect 85238 346294 85294 346350
rect 85362 346294 85418 346350
rect 85238 346170 85294 346226
rect 85362 346170 85418 346226
rect 85238 346046 85294 346102
rect 85362 346046 85418 346102
rect 85238 345922 85294 345978
rect 85362 345922 85418 345978
rect 39954 334294 40010 334350
rect 40078 334294 40134 334350
rect 40202 334294 40258 334350
rect 40326 334294 40382 334350
rect 39954 334170 40010 334226
rect 40078 334170 40134 334226
rect 40202 334170 40258 334226
rect 40326 334170 40382 334226
rect 39954 334046 40010 334102
rect 40078 334046 40134 334102
rect 40202 334046 40258 334102
rect 40326 334046 40382 334102
rect 39954 333922 40010 333978
rect 40078 333922 40134 333978
rect 40202 333922 40258 333978
rect 40326 333922 40382 333978
rect 54518 328294 54574 328350
rect 54642 328294 54698 328350
rect 54518 328170 54574 328226
rect 54642 328170 54698 328226
rect 54518 328046 54574 328102
rect 54642 328046 54698 328102
rect 54518 327922 54574 327978
rect 54642 327922 54698 327978
rect 69878 334294 69934 334350
rect 70002 334294 70058 334350
rect 69878 334170 69934 334226
rect 70002 334170 70058 334226
rect 69878 334046 69934 334102
rect 70002 334046 70058 334102
rect 69878 333922 69934 333978
rect 70002 333922 70058 333978
rect 70674 334294 70730 334350
rect 70798 334294 70854 334350
rect 70922 334294 70978 334350
rect 71046 334294 71102 334350
rect 70674 334170 70730 334226
rect 70798 334170 70854 334226
rect 70922 334170 70978 334226
rect 71046 334170 71102 334226
rect 70674 334046 70730 334102
rect 70798 334046 70854 334102
rect 70922 334046 70978 334102
rect 71046 334046 71102 334102
rect 70674 333922 70730 333978
rect 70798 333922 70854 333978
rect 70922 333922 70978 333978
rect 71046 333922 71102 333978
rect 66954 328294 67010 328350
rect 67078 328294 67134 328350
rect 67202 328294 67258 328350
rect 67326 328294 67382 328350
rect 66954 328170 67010 328226
rect 67078 328170 67134 328226
rect 67202 328170 67258 328226
rect 67326 328170 67382 328226
rect 66954 328046 67010 328102
rect 67078 328046 67134 328102
rect 67202 328046 67258 328102
rect 67326 328046 67382 328102
rect 66954 327922 67010 327978
rect 67078 327922 67134 327978
rect 67202 327922 67258 327978
rect 67326 327922 67382 327978
rect 39954 316294 40010 316350
rect 40078 316294 40134 316350
rect 40202 316294 40258 316350
rect 40326 316294 40382 316350
rect 39954 316170 40010 316226
rect 40078 316170 40134 316226
rect 40202 316170 40258 316226
rect 40326 316170 40382 316226
rect 39954 316046 40010 316102
rect 40078 316046 40134 316102
rect 40202 316046 40258 316102
rect 40326 316046 40382 316102
rect 39954 315922 40010 315978
rect 40078 315922 40134 315978
rect 40202 315922 40258 315978
rect 40326 315922 40382 315978
rect 39954 298294 40010 298350
rect 40078 298294 40134 298350
rect 40202 298294 40258 298350
rect 40326 298294 40382 298350
rect 39954 298170 40010 298226
rect 40078 298170 40134 298226
rect 40202 298170 40258 298226
rect 40326 298170 40382 298226
rect 39954 298046 40010 298102
rect 40078 298046 40134 298102
rect 40202 298046 40258 298102
rect 40326 298046 40382 298102
rect 39954 297922 40010 297978
rect 40078 297922 40134 297978
rect 40202 297922 40258 297978
rect 40326 297922 40382 297978
rect 60396 311642 60452 311698
rect 66954 310294 67010 310350
rect 67078 310294 67134 310350
rect 67202 310294 67258 310350
rect 67326 310294 67382 310350
rect 66954 310170 67010 310226
rect 67078 310170 67134 310226
rect 67202 310170 67258 310226
rect 67326 310170 67382 310226
rect 66954 310046 67010 310102
rect 67078 310046 67134 310102
rect 67202 310046 67258 310102
rect 67326 310046 67382 310102
rect 66954 309922 67010 309978
rect 67078 309922 67134 309978
rect 67202 309922 67258 309978
rect 67326 309922 67382 309978
rect 66954 292294 67010 292350
rect 67078 292294 67134 292350
rect 67202 292294 67258 292350
rect 67326 292294 67382 292350
rect 66954 292170 67010 292226
rect 67078 292170 67134 292226
rect 67202 292170 67258 292226
rect 67326 292170 67382 292226
rect 66954 292046 67010 292102
rect 67078 292046 67134 292102
rect 67202 292046 67258 292102
rect 67326 292046 67382 292102
rect 66954 291922 67010 291978
rect 67078 291922 67134 291978
rect 67202 291922 67258 291978
rect 67326 291922 67382 291978
rect 91644 356102 91700 356158
rect 91644 332702 91700 332758
rect 91532 330902 91588 330958
rect 85238 328294 85294 328350
rect 85362 328294 85418 328350
rect 85238 328170 85294 328226
rect 85362 328170 85418 328226
rect 85238 328046 85294 328102
rect 85362 328046 85418 328102
rect 85238 327922 85294 327978
rect 85362 327922 85418 327978
rect 70674 316294 70730 316350
rect 70798 316294 70854 316350
rect 70922 316294 70978 316350
rect 71046 316294 71102 316350
rect 70674 316170 70730 316226
rect 70798 316170 70854 316226
rect 70922 316170 70978 316226
rect 71046 316170 71102 316226
rect 70674 316046 70730 316102
rect 70798 316046 70854 316102
rect 70922 316046 70978 316102
rect 71046 316046 71102 316102
rect 70674 315922 70730 315978
rect 70798 315922 70854 315978
rect 70922 315922 70978 315978
rect 71046 315922 71102 315978
rect 70674 298294 70730 298350
rect 70798 298294 70854 298350
rect 70922 298294 70978 298350
rect 71046 298294 71102 298350
rect 70674 298170 70730 298226
rect 70798 298170 70854 298226
rect 70922 298170 70978 298226
rect 71046 298170 71102 298226
rect 70674 298046 70730 298102
rect 70798 298046 70854 298102
rect 70922 298046 70978 298102
rect 71046 298046 71102 298102
rect 70674 297922 70730 297978
rect 70798 297922 70854 297978
rect 70922 297922 70978 297978
rect 71046 297922 71102 297978
rect 71820 294002 71876 294058
rect 84588 293822 84644 293878
rect 39954 280294 40010 280350
rect 40078 280294 40134 280350
rect 40202 280294 40258 280350
rect 40326 280294 40382 280350
rect 39954 280170 40010 280226
rect 40078 280170 40134 280226
rect 40202 280170 40258 280226
rect 40326 280170 40382 280226
rect 39954 280046 40010 280102
rect 40078 280046 40134 280102
rect 40202 280046 40258 280102
rect 40326 280046 40382 280102
rect 39954 279922 40010 279978
rect 40078 279922 40134 279978
rect 40202 279922 40258 279978
rect 40326 279922 40382 279978
rect 59878 280294 59934 280350
rect 60002 280294 60058 280350
rect 59878 280170 59934 280226
rect 60002 280170 60058 280226
rect 59878 280046 59934 280102
rect 60002 280046 60058 280102
rect 59878 279922 59934 279978
rect 60002 279922 60058 279978
rect 44518 274294 44574 274350
rect 44642 274294 44698 274350
rect 44518 274170 44574 274226
rect 44642 274170 44698 274226
rect 44518 274046 44574 274102
rect 44642 274046 44698 274102
rect 44518 273922 44574 273978
rect 44642 273922 44698 273978
rect 75238 274294 75294 274350
rect 75362 274294 75418 274350
rect 75238 274170 75294 274226
rect 75362 274170 75418 274226
rect 75238 274046 75294 274102
rect 75362 274046 75418 274102
rect 75238 273922 75294 273978
rect 75362 273922 75418 273978
rect 39954 262294 40010 262350
rect 40078 262294 40134 262350
rect 40202 262294 40258 262350
rect 40326 262294 40382 262350
rect 39954 262170 40010 262226
rect 40078 262170 40134 262226
rect 40202 262170 40258 262226
rect 40326 262170 40382 262226
rect 39954 262046 40010 262102
rect 40078 262046 40134 262102
rect 40202 262046 40258 262102
rect 40326 262046 40382 262102
rect 39954 261922 40010 261978
rect 40078 261922 40134 261978
rect 40202 261922 40258 261978
rect 40326 261922 40382 261978
rect 59878 262294 59934 262350
rect 60002 262294 60058 262350
rect 59878 262170 59934 262226
rect 60002 262170 60058 262226
rect 59878 262046 59934 262102
rect 60002 262046 60058 262102
rect 59878 261922 59934 261978
rect 60002 261922 60058 261978
rect 97674 400294 97730 400350
rect 97798 400294 97854 400350
rect 97922 400294 97978 400350
rect 98046 400294 98102 400350
rect 97674 400170 97730 400226
rect 97798 400170 97854 400226
rect 97922 400170 97978 400226
rect 98046 400170 98102 400226
rect 97674 400046 97730 400102
rect 97798 400046 97854 400102
rect 97922 400046 97978 400102
rect 98046 400046 98102 400102
rect 97674 399922 97730 399978
rect 97798 399922 97854 399978
rect 97922 399922 97978 399978
rect 98046 399922 98102 399978
rect 101394 460294 101450 460350
rect 101518 460294 101574 460350
rect 101642 460294 101698 460350
rect 101766 460294 101822 460350
rect 101394 460170 101450 460226
rect 101518 460170 101574 460226
rect 101642 460170 101698 460226
rect 101766 460170 101822 460226
rect 101394 460046 101450 460102
rect 101518 460046 101574 460102
rect 101642 460046 101698 460102
rect 101766 460046 101822 460102
rect 101394 459922 101450 459978
rect 101518 459922 101574 459978
rect 101642 459922 101698 459978
rect 101766 459922 101822 459978
rect 101394 442294 101450 442350
rect 101518 442294 101574 442350
rect 101642 442294 101698 442350
rect 101766 442294 101822 442350
rect 101394 442170 101450 442226
rect 101518 442170 101574 442226
rect 101642 442170 101698 442226
rect 101766 442170 101822 442226
rect 101394 442046 101450 442102
rect 101518 442046 101574 442102
rect 101642 442046 101698 442102
rect 101766 442046 101822 442102
rect 101394 441922 101450 441978
rect 101518 441922 101574 441978
rect 101642 441922 101698 441978
rect 101766 441922 101822 441978
rect 101394 424294 101450 424350
rect 101518 424294 101574 424350
rect 101642 424294 101698 424350
rect 101766 424294 101822 424350
rect 101394 424170 101450 424226
rect 101518 424170 101574 424226
rect 101642 424170 101698 424226
rect 101766 424170 101822 424226
rect 101394 424046 101450 424102
rect 101518 424046 101574 424102
rect 101642 424046 101698 424102
rect 101766 424046 101822 424102
rect 101394 423922 101450 423978
rect 101518 423922 101574 423978
rect 101642 423922 101698 423978
rect 101766 423922 101822 423978
rect 101394 406294 101450 406350
rect 101518 406294 101574 406350
rect 101642 406294 101698 406350
rect 101766 406294 101822 406350
rect 101394 406170 101450 406226
rect 101518 406170 101574 406226
rect 101642 406170 101698 406226
rect 101766 406170 101822 406226
rect 101394 406046 101450 406102
rect 101518 406046 101574 406102
rect 101642 406046 101698 406102
rect 101766 406046 101822 406102
rect 101394 405922 101450 405978
rect 101518 405922 101574 405978
rect 101642 405922 101698 405978
rect 101766 405922 101822 405978
rect 101394 388294 101450 388350
rect 101518 388294 101574 388350
rect 101642 388294 101698 388350
rect 101766 388294 101822 388350
rect 101394 388170 101450 388226
rect 101518 388170 101574 388226
rect 101642 388170 101698 388226
rect 101766 388170 101822 388226
rect 101394 388046 101450 388102
rect 101518 388046 101574 388102
rect 101642 388046 101698 388102
rect 101766 388046 101822 388102
rect 101394 387922 101450 387978
rect 101518 387922 101574 387978
rect 101642 387922 101698 387978
rect 101766 387922 101822 387978
rect 97674 382294 97730 382350
rect 97798 382294 97854 382350
rect 97922 382294 97978 382350
rect 98046 382294 98102 382350
rect 97674 382170 97730 382226
rect 97798 382170 97854 382226
rect 97922 382170 97978 382226
rect 98046 382170 98102 382226
rect 97674 382046 97730 382102
rect 97798 382046 97854 382102
rect 97922 382046 97978 382102
rect 98046 382046 98102 382102
rect 97674 381922 97730 381978
rect 97798 381922 97854 381978
rect 97922 381922 97978 381978
rect 98046 381922 98102 381978
rect 97674 364294 97730 364350
rect 97798 364294 97854 364350
rect 97922 364294 97978 364350
rect 98046 364294 98102 364350
rect 97674 364170 97730 364226
rect 97798 364170 97854 364226
rect 97922 364170 97978 364226
rect 98046 364170 98102 364226
rect 97674 364046 97730 364102
rect 97798 364046 97854 364102
rect 97922 364046 97978 364102
rect 98046 364046 98102 364102
rect 97674 363922 97730 363978
rect 97798 363922 97854 363978
rect 97922 363922 97978 363978
rect 98046 363922 98102 363978
rect 93212 330902 93268 330958
rect 93212 320822 93268 320878
rect 44518 256294 44574 256350
rect 44642 256294 44698 256350
rect 44518 256170 44574 256226
rect 44642 256170 44698 256226
rect 44518 256046 44574 256102
rect 44642 256046 44698 256102
rect 44518 255922 44574 255978
rect 44642 255922 44698 255978
rect 75238 256294 75294 256350
rect 75362 256294 75418 256350
rect 75238 256170 75294 256226
rect 75362 256170 75418 256226
rect 75238 256046 75294 256102
rect 75362 256046 75418 256102
rect 75238 255922 75294 255978
rect 75362 255922 75418 255978
rect 39954 244294 40010 244350
rect 40078 244294 40134 244350
rect 40202 244294 40258 244350
rect 40326 244294 40382 244350
rect 39954 244170 40010 244226
rect 40078 244170 40134 244226
rect 40202 244170 40258 244226
rect 40326 244170 40382 244226
rect 39954 244046 40010 244102
rect 40078 244046 40134 244102
rect 40202 244046 40258 244102
rect 40326 244046 40382 244102
rect 39954 243922 40010 243978
rect 40078 243922 40134 243978
rect 40202 243922 40258 243978
rect 40326 243922 40382 243978
rect 36234 220294 36290 220350
rect 36358 220294 36414 220350
rect 36482 220294 36538 220350
rect 36606 220294 36662 220350
rect 36234 220170 36290 220226
rect 36358 220170 36414 220226
rect 36482 220170 36538 220226
rect 36606 220170 36662 220226
rect 36234 220046 36290 220102
rect 36358 220046 36414 220102
rect 36482 220046 36538 220102
rect 36606 220046 36662 220102
rect 36234 219922 36290 219978
rect 36358 219922 36414 219978
rect 36482 219922 36538 219978
rect 36606 219922 36662 219978
rect 33516 4922 33572 4978
rect 35196 4742 35252 4798
rect 36234 202294 36290 202350
rect 36358 202294 36414 202350
rect 36482 202294 36538 202350
rect 36606 202294 36662 202350
rect 36234 202170 36290 202226
rect 36358 202170 36414 202226
rect 36482 202170 36538 202226
rect 36606 202170 36662 202226
rect 36234 202046 36290 202102
rect 36358 202046 36414 202102
rect 36482 202046 36538 202102
rect 36606 202046 36662 202102
rect 36234 201922 36290 201978
rect 36358 201922 36414 201978
rect 36482 201922 36538 201978
rect 36606 201922 36662 201978
rect 36234 184294 36290 184350
rect 36358 184294 36414 184350
rect 36482 184294 36538 184350
rect 36606 184294 36662 184350
rect 36234 184170 36290 184226
rect 36358 184170 36414 184226
rect 36482 184170 36538 184226
rect 36606 184170 36662 184226
rect 36234 184046 36290 184102
rect 36358 184046 36414 184102
rect 36482 184046 36538 184102
rect 36606 184046 36662 184102
rect 36234 183922 36290 183978
rect 36358 183922 36414 183978
rect 36482 183922 36538 183978
rect 36606 183922 36662 183978
rect 36234 166294 36290 166350
rect 36358 166294 36414 166350
rect 36482 166294 36538 166350
rect 36606 166294 36662 166350
rect 36234 166170 36290 166226
rect 36358 166170 36414 166226
rect 36482 166170 36538 166226
rect 36606 166170 36662 166226
rect 36234 166046 36290 166102
rect 36358 166046 36414 166102
rect 36482 166046 36538 166102
rect 36606 166046 36662 166102
rect 36234 165922 36290 165978
rect 36358 165922 36414 165978
rect 36482 165922 36538 165978
rect 36606 165922 36662 165978
rect 36234 148294 36290 148350
rect 36358 148294 36414 148350
rect 36482 148294 36538 148350
rect 36606 148294 36662 148350
rect 36234 148170 36290 148226
rect 36358 148170 36414 148226
rect 36482 148170 36538 148226
rect 36606 148170 36662 148226
rect 36234 148046 36290 148102
rect 36358 148046 36414 148102
rect 36482 148046 36538 148102
rect 36606 148046 36662 148102
rect 36234 147922 36290 147978
rect 36358 147922 36414 147978
rect 36482 147922 36538 147978
rect 36606 147922 36662 147978
rect 36234 130294 36290 130350
rect 36358 130294 36414 130350
rect 36482 130294 36538 130350
rect 36606 130294 36662 130350
rect 36234 130170 36290 130226
rect 36358 130170 36414 130226
rect 36482 130170 36538 130226
rect 36606 130170 36662 130226
rect 36234 130046 36290 130102
rect 36358 130046 36414 130102
rect 36482 130046 36538 130102
rect 36606 130046 36662 130102
rect 36234 129922 36290 129978
rect 36358 129922 36414 129978
rect 36482 129922 36538 129978
rect 36606 129922 36662 129978
rect 36234 112294 36290 112350
rect 36358 112294 36414 112350
rect 36482 112294 36538 112350
rect 36606 112294 36662 112350
rect 36234 112170 36290 112226
rect 36358 112170 36414 112226
rect 36482 112170 36538 112226
rect 36606 112170 36662 112226
rect 36234 112046 36290 112102
rect 36358 112046 36414 112102
rect 36482 112046 36538 112102
rect 36606 112046 36662 112102
rect 36234 111922 36290 111978
rect 36358 111922 36414 111978
rect 36482 111922 36538 111978
rect 36606 111922 36662 111978
rect 36234 94294 36290 94350
rect 36358 94294 36414 94350
rect 36482 94294 36538 94350
rect 36606 94294 36662 94350
rect 36234 94170 36290 94226
rect 36358 94170 36414 94226
rect 36482 94170 36538 94226
rect 36606 94170 36662 94226
rect 36234 94046 36290 94102
rect 36358 94046 36414 94102
rect 36482 94046 36538 94102
rect 36606 94046 36662 94102
rect 36234 93922 36290 93978
rect 36358 93922 36414 93978
rect 36482 93922 36538 93978
rect 36606 93922 36662 93978
rect 36234 76294 36290 76350
rect 36358 76294 36414 76350
rect 36482 76294 36538 76350
rect 36606 76294 36662 76350
rect 36234 76170 36290 76226
rect 36358 76170 36414 76226
rect 36482 76170 36538 76226
rect 36606 76170 36662 76226
rect 36234 76046 36290 76102
rect 36358 76046 36414 76102
rect 36482 76046 36538 76102
rect 36606 76046 36662 76102
rect 36234 75922 36290 75978
rect 36358 75922 36414 75978
rect 36482 75922 36538 75978
rect 36606 75922 36662 75978
rect 36234 58294 36290 58350
rect 36358 58294 36414 58350
rect 36482 58294 36538 58350
rect 36606 58294 36662 58350
rect 36234 58170 36290 58226
rect 36358 58170 36414 58226
rect 36482 58170 36538 58226
rect 36606 58170 36662 58226
rect 36234 58046 36290 58102
rect 36358 58046 36414 58102
rect 36482 58046 36538 58102
rect 36606 58046 36662 58102
rect 36234 57922 36290 57978
rect 36358 57922 36414 57978
rect 36482 57922 36538 57978
rect 36606 57922 36662 57978
rect 36234 40294 36290 40350
rect 36358 40294 36414 40350
rect 36482 40294 36538 40350
rect 36606 40294 36662 40350
rect 36234 40170 36290 40226
rect 36358 40170 36414 40226
rect 36482 40170 36538 40226
rect 36606 40170 36662 40226
rect 36234 40046 36290 40102
rect 36358 40046 36414 40102
rect 36482 40046 36538 40102
rect 36606 40046 36662 40102
rect 36234 39922 36290 39978
rect 36358 39922 36414 39978
rect 36482 39922 36538 39978
rect 36606 39922 36662 39978
rect 36234 22294 36290 22350
rect 36358 22294 36414 22350
rect 36482 22294 36538 22350
rect 36606 22294 36662 22350
rect 36234 22170 36290 22226
rect 36358 22170 36414 22226
rect 36482 22170 36538 22226
rect 36606 22170 36662 22226
rect 36234 22046 36290 22102
rect 36358 22046 36414 22102
rect 36482 22046 36538 22102
rect 36606 22046 36662 22102
rect 36234 21922 36290 21978
rect 36358 21922 36414 21978
rect 36482 21922 36538 21978
rect 36606 21922 36662 21978
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 59878 244294 59934 244350
rect 60002 244294 60058 244350
rect 59878 244170 59934 244226
rect 60002 244170 60058 244226
rect 59878 244046 59934 244102
rect 60002 244046 60058 244102
rect 59878 243922 59934 243978
rect 60002 243922 60058 243978
rect 93660 354302 93716 354358
rect 93324 322442 93380 322498
rect 93436 332702 93492 332758
rect 93436 320642 93492 320698
rect 93660 320462 93716 320518
rect 97674 346294 97730 346350
rect 97798 346294 97854 346350
rect 97922 346294 97978 346350
rect 98046 346294 98102 346350
rect 97674 346170 97730 346226
rect 97798 346170 97854 346226
rect 97922 346170 97978 346226
rect 98046 346170 98102 346226
rect 97674 346046 97730 346102
rect 97798 346046 97854 346102
rect 97922 346046 97978 346102
rect 98046 346046 98102 346102
rect 97674 345922 97730 345978
rect 97798 345922 97854 345978
rect 97922 345922 97978 345978
rect 98046 345922 98102 345978
rect 97674 328294 97730 328350
rect 97798 328294 97854 328350
rect 97922 328294 97978 328350
rect 98046 328294 98102 328350
rect 97674 328170 97730 328226
rect 97798 328170 97854 328226
rect 97922 328170 97978 328226
rect 98046 328170 98102 328226
rect 97674 328046 97730 328102
rect 97798 328046 97854 328102
rect 97922 328046 97978 328102
rect 98046 328046 98102 328102
rect 97674 327922 97730 327978
rect 97798 327922 97854 327978
rect 97922 327922 97978 327978
rect 98046 327922 98102 327978
rect 97674 310294 97730 310350
rect 97798 310294 97854 310350
rect 97922 310294 97978 310350
rect 98046 310294 98102 310350
rect 97674 310170 97730 310226
rect 97798 310170 97854 310226
rect 97922 310170 97978 310226
rect 98046 310170 98102 310226
rect 97674 310046 97730 310102
rect 97798 310046 97854 310102
rect 97922 310046 97978 310102
rect 98046 310046 98102 310102
rect 97674 309922 97730 309978
rect 97798 309922 97854 309978
rect 97922 309922 97978 309978
rect 98046 309922 98102 309978
rect 97674 292294 97730 292350
rect 97798 292294 97854 292350
rect 97922 292294 97978 292350
rect 98046 292294 98102 292350
rect 97674 292170 97730 292226
rect 97798 292170 97854 292226
rect 97922 292170 97978 292226
rect 98046 292170 98102 292226
rect 97674 292046 97730 292102
rect 97798 292046 97854 292102
rect 97922 292046 97978 292102
rect 98046 292046 98102 292102
rect 97674 291922 97730 291978
rect 97798 291922 97854 291978
rect 97922 291922 97978 291978
rect 98046 291922 98102 291978
rect 93996 275642 94052 275698
rect 97674 274294 97730 274350
rect 97798 274294 97854 274350
rect 97922 274294 97978 274350
rect 98046 274294 98102 274350
rect 97674 274170 97730 274226
rect 97798 274170 97854 274226
rect 97922 274170 97978 274226
rect 98046 274170 98102 274226
rect 97674 274046 97730 274102
rect 97798 274046 97854 274102
rect 97922 274046 97978 274102
rect 98046 274046 98102 274102
rect 97674 273922 97730 273978
rect 97798 273922 97854 273978
rect 97922 273922 97978 273978
rect 98046 273922 98102 273978
rect 93996 270602 94052 270658
rect 97674 256294 97730 256350
rect 97798 256294 97854 256350
rect 97922 256294 97978 256350
rect 98046 256294 98102 256350
rect 97674 256170 97730 256226
rect 97798 256170 97854 256226
rect 97922 256170 97978 256226
rect 98046 256170 98102 256226
rect 97674 256046 97730 256102
rect 97798 256046 97854 256102
rect 97922 256046 97978 256102
rect 98046 256046 98102 256102
rect 97674 255922 97730 255978
rect 97798 255922 97854 255978
rect 97922 255922 97978 255978
rect 98046 255922 98102 255978
rect 62636 237662 62692 237718
rect 64428 237482 64484 237538
rect 66954 238294 67010 238350
rect 67078 238294 67134 238350
rect 67202 238294 67258 238350
rect 67326 238294 67382 238350
rect 66954 238170 67010 238226
rect 67078 238170 67134 238226
rect 67202 238170 67258 238226
rect 67326 238170 67382 238226
rect 66954 238046 67010 238102
rect 67078 238046 67134 238102
rect 67202 238046 67258 238102
rect 67326 238046 67382 238102
rect 66954 237922 67010 237978
rect 67078 237922 67134 237978
rect 67202 237922 67258 237978
rect 67326 237922 67382 237978
rect 39954 226294 40010 226350
rect 40078 226294 40134 226350
rect 40202 226294 40258 226350
rect 40326 226294 40382 226350
rect 39954 226170 40010 226226
rect 40078 226170 40134 226226
rect 40202 226170 40258 226226
rect 40326 226170 40382 226226
rect 39954 226046 40010 226102
rect 40078 226046 40134 226102
rect 40202 226046 40258 226102
rect 40326 226046 40382 226102
rect 39954 225922 40010 225978
rect 40078 225922 40134 225978
rect 40202 225922 40258 225978
rect 40326 225922 40382 225978
rect 39954 208294 40010 208350
rect 40078 208294 40134 208350
rect 40202 208294 40258 208350
rect 40326 208294 40382 208350
rect 39954 208170 40010 208226
rect 40078 208170 40134 208226
rect 40202 208170 40258 208226
rect 40326 208170 40382 208226
rect 39954 208046 40010 208102
rect 40078 208046 40134 208102
rect 40202 208046 40258 208102
rect 40326 208046 40382 208102
rect 39954 207922 40010 207978
rect 40078 207922 40134 207978
rect 40202 207922 40258 207978
rect 40326 207922 40382 207978
rect 39954 190294 40010 190350
rect 40078 190294 40134 190350
rect 40202 190294 40258 190350
rect 40326 190294 40382 190350
rect 39954 190170 40010 190226
rect 40078 190170 40134 190226
rect 40202 190170 40258 190226
rect 40326 190170 40382 190226
rect 39954 190046 40010 190102
rect 40078 190046 40134 190102
rect 40202 190046 40258 190102
rect 40326 190046 40382 190102
rect 39954 189922 40010 189978
rect 40078 189922 40134 189978
rect 40202 189922 40258 189978
rect 40326 189922 40382 189978
rect 39954 172294 40010 172350
rect 40078 172294 40134 172350
rect 40202 172294 40258 172350
rect 40326 172294 40382 172350
rect 39954 172170 40010 172226
rect 40078 172170 40134 172226
rect 40202 172170 40258 172226
rect 40326 172170 40382 172226
rect 39954 172046 40010 172102
rect 40078 172046 40134 172102
rect 40202 172046 40258 172102
rect 40326 172046 40382 172102
rect 39954 171922 40010 171978
rect 40078 171922 40134 171978
rect 40202 171922 40258 171978
rect 40326 171922 40382 171978
rect 39954 154294 40010 154350
rect 40078 154294 40134 154350
rect 40202 154294 40258 154350
rect 40326 154294 40382 154350
rect 39954 154170 40010 154226
rect 40078 154170 40134 154226
rect 40202 154170 40258 154226
rect 40326 154170 40382 154226
rect 39954 154046 40010 154102
rect 40078 154046 40134 154102
rect 40202 154046 40258 154102
rect 40326 154046 40382 154102
rect 39954 153922 40010 153978
rect 40078 153922 40134 153978
rect 40202 153922 40258 153978
rect 40326 153922 40382 153978
rect 39954 136294 40010 136350
rect 40078 136294 40134 136350
rect 40202 136294 40258 136350
rect 40326 136294 40382 136350
rect 39954 136170 40010 136226
rect 40078 136170 40134 136226
rect 40202 136170 40258 136226
rect 40326 136170 40382 136226
rect 39954 136046 40010 136102
rect 40078 136046 40134 136102
rect 40202 136046 40258 136102
rect 40326 136046 40382 136102
rect 39954 135922 40010 135978
rect 40078 135922 40134 135978
rect 40202 135922 40258 135978
rect 40326 135922 40382 135978
rect 39954 118294 40010 118350
rect 40078 118294 40134 118350
rect 40202 118294 40258 118350
rect 40326 118294 40382 118350
rect 39954 118170 40010 118226
rect 40078 118170 40134 118226
rect 40202 118170 40258 118226
rect 40326 118170 40382 118226
rect 39954 118046 40010 118102
rect 40078 118046 40134 118102
rect 40202 118046 40258 118102
rect 40326 118046 40382 118102
rect 39954 117922 40010 117978
rect 40078 117922 40134 117978
rect 40202 117922 40258 117978
rect 40326 117922 40382 117978
rect 39954 100294 40010 100350
rect 40078 100294 40134 100350
rect 40202 100294 40258 100350
rect 40326 100294 40382 100350
rect 39954 100170 40010 100226
rect 40078 100170 40134 100226
rect 40202 100170 40258 100226
rect 40326 100170 40382 100226
rect 39954 100046 40010 100102
rect 40078 100046 40134 100102
rect 40202 100046 40258 100102
rect 40326 100046 40382 100102
rect 39954 99922 40010 99978
rect 40078 99922 40134 99978
rect 40202 99922 40258 99978
rect 40326 99922 40382 99978
rect 39954 82294 40010 82350
rect 40078 82294 40134 82350
rect 40202 82294 40258 82350
rect 40326 82294 40382 82350
rect 39954 82170 40010 82226
rect 40078 82170 40134 82226
rect 40202 82170 40258 82226
rect 40326 82170 40382 82226
rect 39954 82046 40010 82102
rect 40078 82046 40134 82102
rect 40202 82046 40258 82102
rect 40326 82046 40382 82102
rect 39954 81922 40010 81978
rect 40078 81922 40134 81978
rect 40202 81922 40258 81978
rect 40326 81922 40382 81978
rect 39954 64294 40010 64350
rect 40078 64294 40134 64350
rect 40202 64294 40258 64350
rect 40326 64294 40382 64350
rect 39954 64170 40010 64226
rect 40078 64170 40134 64226
rect 40202 64170 40258 64226
rect 40326 64170 40382 64226
rect 39954 64046 40010 64102
rect 40078 64046 40134 64102
rect 40202 64046 40258 64102
rect 40326 64046 40382 64102
rect 39954 63922 40010 63978
rect 40078 63922 40134 63978
rect 40202 63922 40258 63978
rect 40326 63922 40382 63978
rect 39954 46294 40010 46350
rect 40078 46294 40134 46350
rect 40202 46294 40258 46350
rect 40326 46294 40382 46350
rect 39954 46170 40010 46226
rect 40078 46170 40134 46226
rect 40202 46170 40258 46226
rect 40326 46170 40382 46226
rect 39954 46046 40010 46102
rect 40078 46046 40134 46102
rect 40202 46046 40258 46102
rect 40326 46046 40382 46102
rect 39954 45922 40010 45978
rect 40078 45922 40134 45978
rect 40202 45922 40258 45978
rect 40326 45922 40382 45978
rect 39954 28294 40010 28350
rect 40078 28294 40134 28350
rect 40202 28294 40258 28350
rect 40326 28294 40382 28350
rect 39954 28170 40010 28226
rect 40078 28170 40134 28226
rect 40202 28170 40258 28226
rect 40326 28170 40382 28226
rect 39954 28046 40010 28102
rect 40078 28046 40134 28102
rect 40202 28046 40258 28102
rect 40326 28046 40382 28102
rect 39954 27922 40010 27978
rect 40078 27922 40134 27978
rect 40202 27922 40258 27978
rect 40326 27922 40382 27978
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 41132 210122 41188 210178
rect 41468 208682 41524 208738
rect 66954 220294 67010 220350
rect 67078 220294 67134 220350
rect 67202 220294 67258 220350
rect 67326 220294 67382 220350
rect 66954 220170 67010 220226
rect 67078 220170 67134 220226
rect 67202 220170 67258 220226
rect 67326 220170 67382 220226
rect 66954 220046 67010 220102
rect 67078 220046 67134 220102
rect 67202 220046 67258 220102
rect 67326 220046 67382 220102
rect 66954 219922 67010 219978
rect 67078 219922 67134 219978
rect 67202 219922 67258 219978
rect 67326 219922 67382 219978
rect 97674 238294 97730 238350
rect 97798 238294 97854 238350
rect 97922 238294 97978 238350
rect 98046 238294 98102 238350
rect 97674 238170 97730 238226
rect 97798 238170 97854 238226
rect 97922 238170 97978 238226
rect 98046 238170 98102 238226
rect 97674 238046 97730 238102
rect 97798 238046 97854 238102
rect 97922 238046 97978 238102
rect 98046 238046 98102 238102
rect 97674 237922 97730 237978
rect 97798 237922 97854 237978
rect 97922 237922 97978 237978
rect 98046 237922 98102 237978
rect 100156 237482 100212 237538
rect 101394 370294 101450 370350
rect 101518 370294 101574 370350
rect 101642 370294 101698 370350
rect 101766 370294 101822 370350
rect 101394 370170 101450 370226
rect 101518 370170 101574 370226
rect 101642 370170 101698 370226
rect 101766 370170 101822 370226
rect 101394 370046 101450 370102
rect 101518 370046 101574 370102
rect 101642 370046 101698 370102
rect 101766 370046 101822 370102
rect 101394 369922 101450 369978
rect 101518 369922 101574 369978
rect 101642 369922 101698 369978
rect 101766 369922 101822 369978
rect 101394 352294 101450 352350
rect 101518 352294 101574 352350
rect 101642 352294 101698 352350
rect 101766 352294 101822 352350
rect 101394 352170 101450 352226
rect 101518 352170 101574 352226
rect 101642 352170 101698 352226
rect 101766 352170 101822 352226
rect 101394 352046 101450 352102
rect 101518 352046 101574 352102
rect 101642 352046 101698 352102
rect 101766 352046 101822 352102
rect 101394 351922 101450 351978
rect 101518 351922 101574 351978
rect 101642 351922 101698 351978
rect 101766 351922 101822 351978
rect 128394 472294 128450 472350
rect 128518 472294 128574 472350
rect 128642 472294 128698 472350
rect 128766 472294 128822 472350
rect 128394 472170 128450 472226
rect 128518 472170 128574 472226
rect 128642 472170 128698 472226
rect 128766 472170 128822 472226
rect 128394 472046 128450 472102
rect 128518 472046 128574 472102
rect 128642 472046 128698 472102
rect 128766 472046 128822 472102
rect 128394 471922 128450 471978
rect 128518 471922 128574 471978
rect 128642 471922 128698 471978
rect 128766 471922 128822 471978
rect 128394 454294 128450 454350
rect 128518 454294 128574 454350
rect 128642 454294 128698 454350
rect 128766 454294 128822 454350
rect 128394 454170 128450 454226
rect 128518 454170 128574 454226
rect 128642 454170 128698 454226
rect 128766 454170 128822 454226
rect 128394 454046 128450 454102
rect 128518 454046 128574 454102
rect 128642 454046 128698 454102
rect 128766 454046 128822 454102
rect 128394 453922 128450 453978
rect 128518 453922 128574 453978
rect 128642 453922 128698 453978
rect 128766 453922 128822 453978
rect 128394 436294 128450 436350
rect 128518 436294 128574 436350
rect 128642 436294 128698 436350
rect 128766 436294 128822 436350
rect 128394 436170 128450 436226
rect 128518 436170 128574 436226
rect 128642 436170 128698 436226
rect 128766 436170 128822 436226
rect 128394 436046 128450 436102
rect 128518 436046 128574 436102
rect 128642 436046 128698 436102
rect 128766 436046 128822 436102
rect 128394 435922 128450 435978
rect 128518 435922 128574 435978
rect 128642 435922 128698 435978
rect 128766 435922 128822 435978
rect 128394 418294 128450 418350
rect 128518 418294 128574 418350
rect 128642 418294 128698 418350
rect 128766 418294 128822 418350
rect 128394 418170 128450 418226
rect 128518 418170 128574 418226
rect 128642 418170 128698 418226
rect 128766 418170 128822 418226
rect 128394 418046 128450 418102
rect 128518 418046 128574 418102
rect 128642 418046 128698 418102
rect 128766 418046 128822 418102
rect 128394 417922 128450 417978
rect 128518 417922 128574 417978
rect 128642 417922 128698 417978
rect 128766 417922 128822 417978
rect 128394 400294 128450 400350
rect 128518 400294 128574 400350
rect 128642 400294 128698 400350
rect 128766 400294 128822 400350
rect 128394 400170 128450 400226
rect 128518 400170 128574 400226
rect 128642 400170 128698 400226
rect 128766 400170 128822 400226
rect 128394 400046 128450 400102
rect 128518 400046 128574 400102
rect 128642 400046 128698 400102
rect 128766 400046 128822 400102
rect 128394 399922 128450 399978
rect 128518 399922 128574 399978
rect 128642 399922 128698 399978
rect 128766 399922 128822 399978
rect 128394 382294 128450 382350
rect 128518 382294 128574 382350
rect 128642 382294 128698 382350
rect 128766 382294 128822 382350
rect 128394 382170 128450 382226
rect 128518 382170 128574 382226
rect 128642 382170 128698 382226
rect 128766 382170 128822 382226
rect 128394 382046 128450 382102
rect 128518 382046 128574 382102
rect 128642 382046 128698 382102
rect 128766 382046 128822 382102
rect 128394 381922 128450 381978
rect 128518 381922 128574 381978
rect 128642 381922 128698 381978
rect 128766 381922 128822 381978
rect 128394 364294 128450 364350
rect 128518 364294 128574 364350
rect 128642 364294 128698 364350
rect 128766 364294 128822 364350
rect 128394 364170 128450 364226
rect 128518 364170 128574 364226
rect 128642 364170 128698 364226
rect 128766 364170 128822 364226
rect 128394 364046 128450 364102
rect 128518 364046 128574 364102
rect 128642 364046 128698 364102
rect 128766 364046 128822 364102
rect 128394 363922 128450 363978
rect 128518 363922 128574 363978
rect 128642 363922 128698 363978
rect 128766 363922 128822 363978
rect 124518 346294 124574 346350
rect 124642 346294 124698 346350
rect 124518 346170 124574 346226
rect 124642 346170 124698 346226
rect 124518 346046 124574 346102
rect 124642 346046 124698 346102
rect 124518 345922 124574 345978
rect 124642 345922 124698 345978
rect 128394 346294 128450 346350
rect 128518 346294 128574 346350
rect 128642 346294 128698 346350
rect 128766 346294 128822 346350
rect 128394 346170 128450 346226
rect 128518 346170 128574 346226
rect 128642 346170 128698 346226
rect 128766 346170 128822 346226
rect 128394 346046 128450 346102
rect 128518 346046 128574 346102
rect 128642 346046 128698 346102
rect 128766 346046 128822 346102
rect 128394 345922 128450 345978
rect 128518 345922 128574 345978
rect 128642 345922 128698 345978
rect 128766 345922 128822 345978
rect 101394 334294 101450 334350
rect 101518 334294 101574 334350
rect 101642 334294 101698 334350
rect 101766 334294 101822 334350
rect 101394 334170 101450 334226
rect 101518 334170 101574 334226
rect 101642 334170 101698 334226
rect 101766 334170 101822 334226
rect 101394 334046 101450 334102
rect 101518 334046 101574 334102
rect 101642 334046 101698 334102
rect 101766 334046 101822 334102
rect 101394 333922 101450 333978
rect 101518 333922 101574 333978
rect 101642 333922 101698 333978
rect 101766 333922 101822 333978
rect 124518 328294 124574 328350
rect 124642 328294 124698 328350
rect 124518 328170 124574 328226
rect 124642 328170 124698 328226
rect 124518 328046 124574 328102
rect 124642 328046 124698 328102
rect 124518 327922 124574 327978
rect 124642 327922 124698 327978
rect 128394 328294 128450 328350
rect 128518 328294 128574 328350
rect 128642 328294 128698 328350
rect 128766 328294 128822 328350
rect 128394 328170 128450 328226
rect 128518 328170 128574 328226
rect 128642 328170 128698 328226
rect 128766 328170 128822 328226
rect 128394 328046 128450 328102
rect 128518 328046 128574 328102
rect 128642 328046 128698 328102
rect 128766 328046 128822 328102
rect 128394 327922 128450 327978
rect 128518 327922 128574 327978
rect 128642 327922 128698 327978
rect 128766 327922 128822 327978
rect 101394 316294 101450 316350
rect 101518 316294 101574 316350
rect 101642 316294 101698 316350
rect 101766 316294 101822 316350
rect 101394 316170 101450 316226
rect 101518 316170 101574 316226
rect 101642 316170 101698 316226
rect 101766 316170 101822 316226
rect 101394 316046 101450 316102
rect 101518 316046 101574 316102
rect 101642 316046 101698 316102
rect 101766 316046 101822 316102
rect 101394 315922 101450 315978
rect 101518 315922 101574 315978
rect 101642 315922 101698 315978
rect 101766 315922 101822 315978
rect 101394 298294 101450 298350
rect 101518 298294 101574 298350
rect 101642 298294 101698 298350
rect 101766 298294 101822 298350
rect 101394 298170 101450 298226
rect 101518 298170 101574 298226
rect 101642 298170 101698 298226
rect 101766 298170 101822 298226
rect 101394 298046 101450 298102
rect 101518 298046 101574 298102
rect 101642 298046 101698 298102
rect 101766 298046 101822 298102
rect 101394 297922 101450 297978
rect 101518 297922 101574 297978
rect 101642 297922 101698 297978
rect 101766 297922 101822 297978
rect 128394 310294 128450 310350
rect 128518 310294 128574 310350
rect 128642 310294 128698 310350
rect 128766 310294 128822 310350
rect 128394 310170 128450 310226
rect 128518 310170 128574 310226
rect 128642 310170 128698 310226
rect 128766 310170 128822 310226
rect 128394 310046 128450 310102
rect 128518 310046 128574 310102
rect 128642 310046 128698 310102
rect 128766 310046 128822 310102
rect 128394 309922 128450 309978
rect 128518 309922 128574 309978
rect 128642 309922 128698 309978
rect 128766 309922 128822 309978
rect 128394 292294 128450 292350
rect 128518 292294 128574 292350
rect 128642 292294 128698 292350
rect 128766 292294 128822 292350
rect 128394 292170 128450 292226
rect 128518 292170 128574 292226
rect 128642 292170 128698 292226
rect 128766 292170 128822 292226
rect 128394 292046 128450 292102
rect 128518 292046 128574 292102
rect 128642 292046 128698 292102
rect 128766 292046 128822 292102
rect 128394 291922 128450 291978
rect 128518 291922 128574 291978
rect 128642 291922 128698 291978
rect 128766 291922 128822 291978
rect 101394 280294 101450 280350
rect 101518 280294 101574 280350
rect 101642 280294 101698 280350
rect 101766 280294 101822 280350
rect 101394 280170 101450 280226
rect 101518 280170 101574 280226
rect 101642 280170 101698 280226
rect 101766 280170 101822 280226
rect 101394 280046 101450 280102
rect 101518 280046 101574 280102
rect 101642 280046 101698 280102
rect 101766 280046 101822 280102
rect 101394 279922 101450 279978
rect 101518 279922 101574 279978
rect 101642 279922 101698 279978
rect 101766 279922 101822 279978
rect 101394 262294 101450 262350
rect 101518 262294 101574 262350
rect 101642 262294 101698 262350
rect 101766 262294 101822 262350
rect 101394 262170 101450 262226
rect 101518 262170 101574 262226
rect 101642 262170 101698 262226
rect 101766 262170 101822 262226
rect 101394 262046 101450 262102
rect 101518 262046 101574 262102
rect 101642 262046 101698 262102
rect 101766 262046 101822 262102
rect 101394 261922 101450 261978
rect 101518 261922 101574 261978
rect 101642 261922 101698 261978
rect 101766 261922 101822 261978
rect 101394 244294 101450 244350
rect 101518 244294 101574 244350
rect 101642 244294 101698 244350
rect 101766 244294 101822 244350
rect 101394 244170 101450 244226
rect 101518 244170 101574 244226
rect 101642 244170 101698 244226
rect 101766 244170 101822 244226
rect 101394 244046 101450 244102
rect 101518 244046 101574 244102
rect 101642 244046 101698 244102
rect 101766 244046 101822 244102
rect 101394 243922 101450 243978
rect 101518 243922 101574 243978
rect 101642 243922 101698 243978
rect 101766 243922 101822 243978
rect 97674 220294 97730 220350
rect 97798 220294 97854 220350
rect 97922 220294 97978 220350
rect 98046 220294 98102 220350
rect 97674 220170 97730 220226
rect 97798 220170 97854 220226
rect 97922 220170 97978 220226
rect 98046 220170 98102 220226
rect 97674 220046 97730 220102
rect 97798 220046 97854 220102
rect 97922 220046 97978 220102
rect 98046 220046 98102 220102
rect 97674 219922 97730 219978
rect 97798 219922 97854 219978
rect 97922 219922 97978 219978
rect 98046 219922 98102 219978
rect 101394 226294 101450 226350
rect 101518 226294 101574 226350
rect 101642 226294 101698 226350
rect 101766 226294 101822 226350
rect 101394 226170 101450 226226
rect 101518 226170 101574 226226
rect 101642 226170 101698 226226
rect 101766 226170 101822 226226
rect 101394 226046 101450 226102
rect 101518 226046 101574 226102
rect 101642 226046 101698 226102
rect 101766 226046 101822 226102
rect 101394 225922 101450 225978
rect 101518 225922 101574 225978
rect 101642 225922 101698 225978
rect 101766 225922 101822 225978
rect 128394 274294 128450 274350
rect 128518 274294 128574 274350
rect 128642 274294 128698 274350
rect 128766 274294 128822 274350
rect 128394 274170 128450 274226
rect 128518 274170 128574 274226
rect 128642 274170 128698 274226
rect 128766 274170 128822 274226
rect 128394 274046 128450 274102
rect 128518 274046 128574 274102
rect 128642 274046 128698 274102
rect 128766 274046 128822 274102
rect 128394 273922 128450 273978
rect 128518 273922 128574 273978
rect 128642 273922 128698 273978
rect 128766 273922 128822 273978
rect 128394 256294 128450 256350
rect 128518 256294 128574 256350
rect 128642 256294 128698 256350
rect 128766 256294 128822 256350
rect 128394 256170 128450 256226
rect 128518 256170 128574 256226
rect 128642 256170 128698 256226
rect 128766 256170 128822 256226
rect 128394 256046 128450 256102
rect 128518 256046 128574 256102
rect 128642 256046 128698 256102
rect 128766 256046 128822 256102
rect 128394 255922 128450 255978
rect 128518 255922 128574 255978
rect 128642 255922 128698 255978
rect 128766 255922 128822 255978
rect 128394 238294 128450 238350
rect 128518 238294 128574 238350
rect 128642 238294 128698 238350
rect 128766 238294 128822 238350
rect 128394 238170 128450 238226
rect 128518 238170 128574 238226
rect 128642 238170 128698 238226
rect 128766 238170 128822 238226
rect 128394 238046 128450 238102
rect 128518 238046 128574 238102
rect 128642 238046 128698 238102
rect 128766 238046 128822 238102
rect 128394 237922 128450 237978
rect 128518 237922 128574 237978
rect 128642 237922 128698 237978
rect 128766 237922 128822 237978
rect 128394 220294 128450 220350
rect 128518 220294 128574 220350
rect 128642 220294 128698 220350
rect 128766 220294 128822 220350
rect 128394 220170 128450 220226
rect 128518 220170 128574 220226
rect 128642 220170 128698 220226
rect 128766 220170 128822 220226
rect 128394 220046 128450 220102
rect 128518 220046 128574 220102
rect 128642 220046 128698 220102
rect 128766 220046 128822 220102
rect 128394 219922 128450 219978
rect 128518 219922 128574 219978
rect 128642 219922 128698 219978
rect 128766 219922 128822 219978
rect 132114 478294 132170 478350
rect 132238 478294 132294 478350
rect 132362 478294 132418 478350
rect 132486 478294 132542 478350
rect 132114 478170 132170 478226
rect 132238 478170 132294 478226
rect 132362 478170 132418 478226
rect 132486 478170 132542 478226
rect 132114 478046 132170 478102
rect 132238 478046 132294 478102
rect 132362 478046 132418 478102
rect 132486 478046 132542 478102
rect 132114 477922 132170 477978
rect 132238 477922 132294 477978
rect 132362 477922 132418 477978
rect 132486 477922 132542 477978
rect 132114 460294 132170 460350
rect 132238 460294 132294 460350
rect 132362 460294 132418 460350
rect 132486 460294 132542 460350
rect 132114 460170 132170 460226
rect 132238 460170 132294 460226
rect 132362 460170 132418 460226
rect 132486 460170 132542 460226
rect 132114 460046 132170 460102
rect 132238 460046 132294 460102
rect 132362 460046 132418 460102
rect 132486 460046 132542 460102
rect 132114 459922 132170 459978
rect 132238 459922 132294 459978
rect 132362 459922 132418 459978
rect 132486 459922 132542 459978
rect 132114 442294 132170 442350
rect 132238 442294 132294 442350
rect 132362 442294 132418 442350
rect 132486 442294 132542 442350
rect 132114 442170 132170 442226
rect 132238 442170 132294 442226
rect 132362 442170 132418 442226
rect 132486 442170 132542 442226
rect 132114 442046 132170 442102
rect 132238 442046 132294 442102
rect 132362 442046 132418 442102
rect 132486 442046 132542 442102
rect 132114 441922 132170 441978
rect 132238 441922 132294 441978
rect 132362 441922 132418 441978
rect 132486 441922 132542 441978
rect 132114 424294 132170 424350
rect 132238 424294 132294 424350
rect 132362 424294 132418 424350
rect 132486 424294 132542 424350
rect 132114 424170 132170 424226
rect 132238 424170 132294 424226
rect 132362 424170 132418 424226
rect 132486 424170 132542 424226
rect 132114 424046 132170 424102
rect 132238 424046 132294 424102
rect 132362 424046 132418 424102
rect 132486 424046 132542 424102
rect 132114 423922 132170 423978
rect 132238 423922 132294 423978
rect 132362 423922 132418 423978
rect 132486 423922 132542 423978
rect 157052 409382 157108 409438
rect 159114 580294 159170 580350
rect 159238 580294 159294 580350
rect 159362 580294 159418 580350
rect 159486 580294 159542 580350
rect 159114 580170 159170 580226
rect 159238 580170 159294 580226
rect 159362 580170 159418 580226
rect 159486 580170 159542 580226
rect 159114 580046 159170 580102
rect 159238 580046 159294 580102
rect 159362 580046 159418 580102
rect 159486 580046 159542 580102
rect 159114 579922 159170 579978
rect 159238 579922 159294 579978
rect 159362 579922 159418 579978
rect 159486 579922 159542 579978
rect 159114 562294 159170 562350
rect 159238 562294 159294 562350
rect 159362 562294 159418 562350
rect 159486 562294 159542 562350
rect 159114 562170 159170 562226
rect 159238 562170 159294 562226
rect 159362 562170 159418 562226
rect 159486 562170 159542 562226
rect 159114 562046 159170 562102
rect 159238 562046 159294 562102
rect 159362 562046 159418 562102
rect 159486 562046 159542 562102
rect 159114 561922 159170 561978
rect 159238 561922 159294 561978
rect 159362 561922 159418 561978
rect 159486 561922 159542 561978
rect 159114 544294 159170 544350
rect 159238 544294 159294 544350
rect 159362 544294 159418 544350
rect 159486 544294 159542 544350
rect 159114 544170 159170 544226
rect 159238 544170 159294 544226
rect 159362 544170 159418 544226
rect 159486 544170 159542 544226
rect 159114 544046 159170 544102
rect 159238 544046 159294 544102
rect 159362 544046 159418 544102
rect 159486 544046 159542 544102
rect 159114 543922 159170 543978
rect 159238 543922 159294 543978
rect 159362 543922 159418 543978
rect 159486 543922 159542 543978
rect 159114 526294 159170 526350
rect 159238 526294 159294 526350
rect 159362 526294 159418 526350
rect 159486 526294 159542 526350
rect 159114 526170 159170 526226
rect 159238 526170 159294 526226
rect 159362 526170 159418 526226
rect 159486 526170 159542 526226
rect 159114 526046 159170 526102
rect 159238 526046 159294 526102
rect 159362 526046 159418 526102
rect 159486 526046 159542 526102
rect 159114 525922 159170 525978
rect 159238 525922 159294 525978
rect 159362 525922 159418 525978
rect 159486 525922 159542 525978
rect 159114 508294 159170 508350
rect 159238 508294 159294 508350
rect 159362 508294 159418 508350
rect 159486 508294 159542 508350
rect 159114 508170 159170 508226
rect 159238 508170 159294 508226
rect 159362 508170 159418 508226
rect 159486 508170 159542 508226
rect 159114 508046 159170 508102
rect 159238 508046 159294 508102
rect 159362 508046 159418 508102
rect 159486 508046 159542 508102
rect 159114 507922 159170 507978
rect 159238 507922 159294 507978
rect 159362 507922 159418 507978
rect 159486 507922 159542 507978
rect 159114 490294 159170 490350
rect 159238 490294 159294 490350
rect 159362 490294 159418 490350
rect 159486 490294 159542 490350
rect 159114 490170 159170 490226
rect 159238 490170 159294 490226
rect 159362 490170 159418 490226
rect 159486 490170 159542 490226
rect 159114 490046 159170 490102
rect 159238 490046 159294 490102
rect 159362 490046 159418 490102
rect 159486 490046 159542 490102
rect 159114 489922 159170 489978
rect 159238 489922 159294 489978
rect 159362 489922 159418 489978
rect 159486 489922 159542 489978
rect 159114 472294 159170 472350
rect 159238 472294 159294 472350
rect 159362 472294 159418 472350
rect 159486 472294 159542 472350
rect 159114 472170 159170 472226
rect 159238 472170 159294 472226
rect 159362 472170 159418 472226
rect 159486 472170 159542 472226
rect 159114 472046 159170 472102
rect 159238 472046 159294 472102
rect 159362 472046 159418 472102
rect 159486 472046 159542 472102
rect 159114 471922 159170 471978
rect 159238 471922 159294 471978
rect 159362 471922 159418 471978
rect 159486 471922 159542 471978
rect 159114 454294 159170 454350
rect 159238 454294 159294 454350
rect 159362 454294 159418 454350
rect 159486 454294 159542 454350
rect 159114 454170 159170 454226
rect 159238 454170 159294 454226
rect 159362 454170 159418 454226
rect 159486 454170 159542 454226
rect 159114 454046 159170 454102
rect 159238 454046 159294 454102
rect 159362 454046 159418 454102
rect 159486 454046 159542 454102
rect 159114 453922 159170 453978
rect 159238 453922 159294 453978
rect 159362 453922 159418 453978
rect 159486 453922 159542 453978
rect 159114 436294 159170 436350
rect 159238 436294 159294 436350
rect 159362 436294 159418 436350
rect 159486 436294 159542 436350
rect 159114 436170 159170 436226
rect 159238 436170 159294 436226
rect 159362 436170 159418 436226
rect 159486 436170 159542 436226
rect 159114 436046 159170 436102
rect 159238 436046 159294 436102
rect 159362 436046 159418 436102
rect 159486 436046 159542 436102
rect 159114 435922 159170 435978
rect 159238 435922 159294 435978
rect 159362 435922 159418 435978
rect 159486 435922 159542 435978
rect 159114 418294 159170 418350
rect 159238 418294 159294 418350
rect 159362 418294 159418 418350
rect 159486 418294 159542 418350
rect 159114 418170 159170 418226
rect 159238 418170 159294 418226
rect 159362 418170 159418 418226
rect 159486 418170 159542 418226
rect 159114 418046 159170 418102
rect 159238 418046 159294 418102
rect 159362 418046 159418 418102
rect 159486 418046 159542 418102
rect 159114 417922 159170 417978
rect 159238 417922 159294 417978
rect 159362 417922 159418 417978
rect 159486 417922 159542 417978
rect 150332 407942 150388 407998
rect 132114 406294 132170 406350
rect 132238 406294 132294 406350
rect 132362 406294 132418 406350
rect 132486 406294 132542 406350
rect 132114 406170 132170 406226
rect 132238 406170 132294 406226
rect 132362 406170 132418 406226
rect 132486 406170 132542 406226
rect 132114 406046 132170 406102
rect 132238 406046 132294 406102
rect 132362 406046 132418 406102
rect 132486 406046 132542 406102
rect 132114 405922 132170 405978
rect 132238 405922 132294 405978
rect 132362 405922 132418 405978
rect 132486 405922 132542 405978
rect 132114 388294 132170 388350
rect 132238 388294 132294 388350
rect 132362 388294 132418 388350
rect 132486 388294 132542 388350
rect 132114 388170 132170 388226
rect 132238 388170 132294 388226
rect 132362 388170 132418 388226
rect 132486 388170 132542 388226
rect 132114 388046 132170 388102
rect 132238 388046 132294 388102
rect 132362 388046 132418 388102
rect 132486 388046 132542 388102
rect 132114 387922 132170 387978
rect 132238 387922 132294 387978
rect 132362 387922 132418 387978
rect 132486 387922 132542 387978
rect 132114 370294 132170 370350
rect 132238 370294 132294 370350
rect 132362 370294 132418 370350
rect 132486 370294 132542 370350
rect 132114 370170 132170 370226
rect 132238 370170 132294 370226
rect 132362 370170 132418 370226
rect 132486 370170 132542 370226
rect 132114 370046 132170 370102
rect 132238 370046 132294 370102
rect 132362 370046 132418 370102
rect 132486 370046 132542 370102
rect 132114 369922 132170 369978
rect 132238 369922 132294 369978
rect 132362 369922 132418 369978
rect 132486 369922 132542 369978
rect 159114 400294 159170 400350
rect 159238 400294 159294 400350
rect 159362 400294 159418 400350
rect 159486 400294 159542 400350
rect 159114 400170 159170 400226
rect 159238 400170 159294 400226
rect 159362 400170 159418 400226
rect 159486 400170 159542 400226
rect 159114 400046 159170 400102
rect 159238 400046 159294 400102
rect 159362 400046 159418 400102
rect 159486 400046 159542 400102
rect 159114 399922 159170 399978
rect 159238 399922 159294 399978
rect 159362 399922 159418 399978
rect 159486 399922 159542 399978
rect 159114 382294 159170 382350
rect 159238 382294 159294 382350
rect 159362 382294 159418 382350
rect 159486 382294 159542 382350
rect 159114 382170 159170 382226
rect 159238 382170 159294 382226
rect 159362 382170 159418 382226
rect 159486 382170 159542 382226
rect 159114 382046 159170 382102
rect 159238 382046 159294 382102
rect 159362 382046 159418 382102
rect 159486 382046 159542 382102
rect 159114 381922 159170 381978
rect 159238 381922 159294 381978
rect 159362 381922 159418 381978
rect 159486 381922 159542 381978
rect 159114 364294 159170 364350
rect 159238 364294 159294 364350
rect 159362 364294 159418 364350
rect 159486 364294 159542 364350
rect 159114 364170 159170 364226
rect 159238 364170 159294 364226
rect 159362 364170 159418 364226
rect 159486 364170 159542 364226
rect 159114 364046 159170 364102
rect 159238 364046 159294 364102
rect 159362 364046 159418 364102
rect 159486 364046 159542 364102
rect 159114 363922 159170 363978
rect 159238 363922 159294 363978
rect 159362 363922 159418 363978
rect 159486 363922 159542 363978
rect 132114 352294 132170 352350
rect 132238 352294 132294 352350
rect 132362 352294 132418 352350
rect 132486 352294 132542 352350
rect 132114 352170 132170 352226
rect 132238 352170 132294 352226
rect 132362 352170 132418 352226
rect 132486 352170 132542 352226
rect 132114 352046 132170 352102
rect 132238 352046 132294 352102
rect 132362 352046 132418 352102
rect 132486 352046 132542 352102
rect 132114 351922 132170 351978
rect 132238 351922 132294 351978
rect 132362 351922 132418 351978
rect 132486 351922 132542 351978
rect 139878 352294 139934 352350
rect 140002 352294 140058 352350
rect 139878 352170 139934 352226
rect 140002 352170 140058 352226
rect 139878 352046 139934 352102
rect 140002 352046 140058 352102
rect 139878 351922 139934 351978
rect 140002 351922 140058 351978
rect 155238 346294 155294 346350
rect 155362 346294 155418 346350
rect 155238 346170 155294 346226
rect 155362 346170 155418 346226
rect 155238 346046 155294 346102
rect 155362 346046 155418 346102
rect 155238 345922 155294 345978
rect 155362 345922 155418 345978
rect 159114 346294 159170 346350
rect 159238 346294 159294 346350
rect 159362 346294 159418 346350
rect 159486 346294 159542 346350
rect 159114 346170 159170 346226
rect 159238 346170 159294 346226
rect 159362 346170 159418 346226
rect 159486 346170 159542 346226
rect 159114 346046 159170 346102
rect 159238 346046 159294 346102
rect 159362 346046 159418 346102
rect 159486 346046 159542 346102
rect 159114 345922 159170 345978
rect 159238 345922 159294 345978
rect 159362 345922 159418 345978
rect 159486 345922 159542 345978
rect 132114 334294 132170 334350
rect 132238 334294 132294 334350
rect 132362 334294 132418 334350
rect 132486 334294 132542 334350
rect 132114 334170 132170 334226
rect 132238 334170 132294 334226
rect 132362 334170 132418 334226
rect 132486 334170 132542 334226
rect 132114 334046 132170 334102
rect 132238 334046 132294 334102
rect 132362 334046 132418 334102
rect 132486 334046 132542 334102
rect 132114 333922 132170 333978
rect 132238 333922 132294 333978
rect 132362 333922 132418 333978
rect 132486 333922 132542 333978
rect 139878 334294 139934 334350
rect 140002 334294 140058 334350
rect 139878 334170 139934 334226
rect 140002 334170 140058 334226
rect 139878 334046 139934 334102
rect 140002 334046 140058 334102
rect 139878 333922 139934 333978
rect 140002 333922 140058 333978
rect 155238 328294 155294 328350
rect 155362 328294 155418 328350
rect 155238 328170 155294 328226
rect 155362 328170 155418 328226
rect 155238 328046 155294 328102
rect 155362 328046 155418 328102
rect 155238 327922 155294 327978
rect 155362 327922 155418 327978
rect 159114 328294 159170 328350
rect 159238 328294 159294 328350
rect 159362 328294 159418 328350
rect 159486 328294 159542 328350
rect 159114 328170 159170 328226
rect 159238 328170 159294 328226
rect 159362 328170 159418 328226
rect 159486 328170 159542 328226
rect 159114 328046 159170 328102
rect 159238 328046 159294 328102
rect 159362 328046 159418 328102
rect 159486 328046 159542 328102
rect 159114 327922 159170 327978
rect 159238 327922 159294 327978
rect 159362 327922 159418 327978
rect 159486 327922 159542 327978
rect 132114 316294 132170 316350
rect 132238 316294 132294 316350
rect 132362 316294 132418 316350
rect 132486 316294 132542 316350
rect 132114 316170 132170 316226
rect 132238 316170 132294 316226
rect 132362 316170 132418 316226
rect 132486 316170 132542 316226
rect 132114 316046 132170 316102
rect 132238 316046 132294 316102
rect 132362 316046 132418 316102
rect 132486 316046 132542 316102
rect 132114 315922 132170 315978
rect 132238 315922 132294 315978
rect 132362 315922 132418 315978
rect 132486 315922 132542 315978
rect 132114 298294 132170 298350
rect 132238 298294 132294 298350
rect 132362 298294 132418 298350
rect 132486 298294 132542 298350
rect 132114 298170 132170 298226
rect 132238 298170 132294 298226
rect 132362 298170 132418 298226
rect 132486 298170 132542 298226
rect 132114 298046 132170 298102
rect 132238 298046 132294 298102
rect 132362 298046 132418 298102
rect 132486 298046 132542 298102
rect 132114 297922 132170 297978
rect 132238 297922 132294 297978
rect 132362 297922 132418 297978
rect 132486 297922 132542 297978
rect 159114 310294 159170 310350
rect 159238 310294 159294 310350
rect 159362 310294 159418 310350
rect 159486 310294 159542 310350
rect 159114 310170 159170 310226
rect 159238 310170 159294 310226
rect 159362 310170 159418 310226
rect 159486 310170 159542 310226
rect 159114 310046 159170 310102
rect 159238 310046 159294 310102
rect 159362 310046 159418 310102
rect 159486 310046 159542 310102
rect 159114 309922 159170 309978
rect 159238 309922 159294 309978
rect 159362 309922 159418 309978
rect 159486 309922 159542 309978
rect 159114 292294 159170 292350
rect 159238 292294 159294 292350
rect 159362 292294 159418 292350
rect 159486 292294 159542 292350
rect 159114 292170 159170 292226
rect 159238 292170 159294 292226
rect 159362 292170 159418 292226
rect 159486 292170 159542 292226
rect 159114 292046 159170 292102
rect 159238 292046 159294 292102
rect 159362 292046 159418 292102
rect 159486 292046 159542 292102
rect 159114 291922 159170 291978
rect 159238 291922 159294 291978
rect 159362 291922 159418 291978
rect 159486 291922 159542 291978
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 162834 568294 162890 568350
rect 162958 568294 163014 568350
rect 163082 568294 163138 568350
rect 163206 568294 163262 568350
rect 162834 568170 162890 568226
rect 162958 568170 163014 568226
rect 163082 568170 163138 568226
rect 163206 568170 163262 568226
rect 162834 568046 162890 568102
rect 162958 568046 163014 568102
rect 163082 568046 163138 568102
rect 163206 568046 163262 568102
rect 162834 567922 162890 567978
rect 162958 567922 163014 567978
rect 163082 567922 163138 567978
rect 163206 567922 163262 567978
rect 162834 550294 162890 550350
rect 162958 550294 163014 550350
rect 163082 550294 163138 550350
rect 163206 550294 163262 550350
rect 162834 550170 162890 550226
rect 162958 550170 163014 550226
rect 163082 550170 163138 550226
rect 163206 550170 163262 550226
rect 162834 550046 162890 550102
rect 162958 550046 163014 550102
rect 163082 550046 163138 550102
rect 163206 550046 163262 550102
rect 162834 549922 162890 549978
rect 162958 549922 163014 549978
rect 163082 549922 163138 549978
rect 163206 549922 163262 549978
rect 162834 532294 162890 532350
rect 162958 532294 163014 532350
rect 163082 532294 163138 532350
rect 163206 532294 163262 532350
rect 162834 532170 162890 532226
rect 162958 532170 163014 532226
rect 163082 532170 163138 532226
rect 163206 532170 163262 532226
rect 162834 532046 162890 532102
rect 162958 532046 163014 532102
rect 163082 532046 163138 532102
rect 163206 532046 163262 532102
rect 162834 531922 162890 531978
rect 162958 531922 163014 531978
rect 163082 531922 163138 531978
rect 163206 531922 163262 531978
rect 162834 514294 162890 514350
rect 162958 514294 163014 514350
rect 163082 514294 163138 514350
rect 163206 514294 163262 514350
rect 162834 514170 162890 514226
rect 162958 514170 163014 514226
rect 163082 514170 163138 514226
rect 163206 514170 163262 514226
rect 162834 514046 162890 514102
rect 162958 514046 163014 514102
rect 163082 514046 163138 514102
rect 163206 514046 163262 514102
rect 162834 513922 162890 513978
rect 162958 513922 163014 513978
rect 163082 513922 163138 513978
rect 163206 513922 163262 513978
rect 162834 496294 162890 496350
rect 162958 496294 163014 496350
rect 163082 496294 163138 496350
rect 163206 496294 163262 496350
rect 162834 496170 162890 496226
rect 162958 496170 163014 496226
rect 163082 496170 163138 496226
rect 163206 496170 163262 496226
rect 162834 496046 162890 496102
rect 162958 496046 163014 496102
rect 163082 496046 163138 496102
rect 163206 496046 163262 496102
rect 162834 495922 162890 495978
rect 162958 495922 163014 495978
rect 163082 495922 163138 495978
rect 163206 495922 163262 495978
rect 162834 478294 162890 478350
rect 162958 478294 163014 478350
rect 163082 478294 163138 478350
rect 163206 478294 163262 478350
rect 162834 478170 162890 478226
rect 162958 478170 163014 478226
rect 163082 478170 163138 478226
rect 163206 478170 163262 478226
rect 162834 478046 162890 478102
rect 162958 478046 163014 478102
rect 163082 478046 163138 478102
rect 163206 478046 163262 478102
rect 162834 477922 162890 477978
rect 162958 477922 163014 477978
rect 163082 477922 163138 477978
rect 163206 477922 163262 477978
rect 162834 460294 162890 460350
rect 162958 460294 163014 460350
rect 163082 460294 163138 460350
rect 163206 460294 163262 460350
rect 162834 460170 162890 460226
rect 162958 460170 163014 460226
rect 163082 460170 163138 460226
rect 163206 460170 163262 460226
rect 162834 460046 162890 460102
rect 162958 460046 163014 460102
rect 163082 460046 163138 460102
rect 163206 460046 163262 460102
rect 162834 459922 162890 459978
rect 162958 459922 163014 459978
rect 163082 459922 163138 459978
rect 163206 459922 163262 459978
rect 162834 442294 162890 442350
rect 162958 442294 163014 442350
rect 163082 442294 163138 442350
rect 163206 442294 163262 442350
rect 162834 442170 162890 442226
rect 162958 442170 163014 442226
rect 163082 442170 163138 442226
rect 163206 442170 163262 442226
rect 162834 442046 162890 442102
rect 162958 442046 163014 442102
rect 163082 442046 163138 442102
rect 163206 442046 163262 442102
rect 162834 441922 162890 441978
rect 162958 441922 163014 441978
rect 163082 441922 163138 441978
rect 163206 441922 163262 441978
rect 162834 424294 162890 424350
rect 162958 424294 163014 424350
rect 163082 424294 163138 424350
rect 163206 424294 163262 424350
rect 162834 424170 162890 424226
rect 162958 424170 163014 424226
rect 163082 424170 163138 424226
rect 163206 424170 163262 424226
rect 162834 424046 162890 424102
rect 162958 424046 163014 424102
rect 163082 424046 163138 424102
rect 163206 424046 163262 424102
rect 162834 423922 162890 423978
rect 162958 423922 163014 423978
rect 163082 423922 163138 423978
rect 163206 423922 163262 423978
rect 162834 406294 162890 406350
rect 162958 406294 163014 406350
rect 163082 406294 163138 406350
rect 163206 406294 163262 406350
rect 162834 406170 162890 406226
rect 162958 406170 163014 406226
rect 163082 406170 163138 406226
rect 163206 406170 163262 406226
rect 162834 406046 162890 406102
rect 162958 406046 163014 406102
rect 163082 406046 163138 406102
rect 163206 406046 163262 406102
rect 162834 405922 162890 405978
rect 162958 405922 163014 405978
rect 163082 405922 163138 405978
rect 163206 405922 163262 405978
rect 162834 388294 162890 388350
rect 162958 388294 163014 388350
rect 163082 388294 163138 388350
rect 163206 388294 163262 388350
rect 162834 388170 162890 388226
rect 162958 388170 163014 388226
rect 163082 388170 163138 388226
rect 163206 388170 163262 388226
rect 162834 388046 162890 388102
rect 162958 388046 163014 388102
rect 163082 388046 163138 388102
rect 163206 388046 163262 388102
rect 162834 387922 162890 387978
rect 162958 387922 163014 387978
rect 163082 387922 163138 387978
rect 163206 387922 163262 387978
rect 162834 370294 162890 370350
rect 162958 370294 163014 370350
rect 163082 370294 163138 370350
rect 163206 370294 163262 370350
rect 162834 370170 162890 370226
rect 162958 370170 163014 370226
rect 163082 370170 163138 370226
rect 163206 370170 163262 370226
rect 162834 370046 162890 370102
rect 162958 370046 163014 370102
rect 163082 370046 163138 370102
rect 163206 370046 163262 370102
rect 162834 369922 162890 369978
rect 162958 369922 163014 369978
rect 163082 369922 163138 369978
rect 163206 369922 163262 369978
rect 162834 352294 162890 352350
rect 162958 352294 163014 352350
rect 163082 352294 163138 352350
rect 163206 352294 163262 352350
rect 162834 352170 162890 352226
rect 162958 352170 163014 352226
rect 163082 352170 163138 352226
rect 163206 352170 163262 352226
rect 162834 352046 162890 352102
rect 162958 352046 163014 352102
rect 163082 352046 163138 352102
rect 163206 352046 163262 352102
rect 162834 351922 162890 351978
rect 162958 351922 163014 351978
rect 163082 351922 163138 351978
rect 163206 351922 163262 351978
rect 162834 334294 162890 334350
rect 162958 334294 163014 334350
rect 163082 334294 163138 334350
rect 163206 334294 163262 334350
rect 162834 334170 162890 334226
rect 162958 334170 163014 334226
rect 163082 334170 163138 334226
rect 163206 334170 163262 334226
rect 162834 334046 162890 334102
rect 162958 334046 163014 334102
rect 163082 334046 163138 334102
rect 163206 334046 163262 334102
rect 162834 333922 162890 333978
rect 162958 333922 163014 333978
rect 163082 333922 163138 333978
rect 163206 333922 163262 333978
rect 162834 316294 162890 316350
rect 162958 316294 163014 316350
rect 163082 316294 163138 316350
rect 163206 316294 163262 316350
rect 162834 316170 162890 316226
rect 162958 316170 163014 316226
rect 163082 316170 163138 316226
rect 163206 316170 163262 316226
rect 162834 316046 162890 316102
rect 162958 316046 163014 316102
rect 163082 316046 163138 316102
rect 163206 316046 163262 316102
rect 162834 315922 162890 315978
rect 162958 315922 163014 315978
rect 163082 315922 163138 315978
rect 163206 315922 163262 315978
rect 162834 298294 162890 298350
rect 162958 298294 163014 298350
rect 163082 298294 163138 298350
rect 163206 298294 163262 298350
rect 162834 298170 162890 298226
rect 162958 298170 163014 298226
rect 163082 298170 163138 298226
rect 163206 298170 163262 298226
rect 162834 298046 162890 298102
rect 162958 298046 163014 298102
rect 163082 298046 163138 298102
rect 163206 298046 163262 298102
rect 162834 297922 162890 297978
rect 162958 297922 163014 297978
rect 163082 297922 163138 297978
rect 163206 297922 163262 297978
rect 132114 280294 132170 280350
rect 132238 280294 132294 280350
rect 132362 280294 132418 280350
rect 132486 280294 132542 280350
rect 132114 280170 132170 280226
rect 132238 280170 132294 280226
rect 132362 280170 132418 280226
rect 132486 280170 132542 280226
rect 132114 280046 132170 280102
rect 132238 280046 132294 280102
rect 132362 280046 132418 280102
rect 132486 280046 132542 280102
rect 132114 279922 132170 279978
rect 132238 279922 132294 279978
rect 132362 279922 132418 279978
rect 132486 279922 132542 279978
rect 147078 280294 147134 280350
rect 147202 280294 147258 280350
rect 147078 280170 147134 280226
rect 147202 280170 147258 280226
rect 147078 280046 147134 280102
rect 147202 280046 147258 280102
rect 147078 279922 147134 279978
rect 147202 279922 147258 279978
rect 152902 280294 152958 280350
rect 153026 280294 153082 280350
rect 152902 280170 152958 280226
rect 153026 280170 153082 280226
rect 152902 280046 152958 280102
rect 153026 280046 153082 280102
rect 152902 279922 152958 279978
rect 153026 279922 153082 279978
rect 158726 280294 158782 280350
rect 158850 280294 158906 280350
rect 158726 280170 158782 280226
rect 158850 280170 158906 280226
rect 158726 280046 158782 280102
rect 158850 280046 158906 280102
rect 158726 279922 158782 279978
rect 158850 279922 158906 279978
rect 164550 280294 164606 280350
rect 164674 280294 164730 280350
rect 164550 280170 164606 280226
rect 164674 280170 164730 280226
rect 164550 280046 164606 280102
rect 164674 280046 164730 280102
rect 164550 279922 164606 279978
rect 164674 279922 164730 279978
rect 153692 275642 153748 275698
rect 144166 274294 144222 274350
rect 144290 274294 144346 274350
rect 144166 274170 144222 274226
rect 144290 274170 144346 274226
rect 144166 274046 144222 274102
rect 144290 274046 144346 274102
rect 144166 273922 144222 273978
rect 144290 273922 144346 273978
rect 149990 274294 150046 274350
rect 150114 274294 150170 274350
rect 149990 274170 150046 274226
rect 150114 274170 150170 274226
rect 149990 274046 150046 274102
rect 150114 274046 150170 274102
rect 149990 273922 150046 273978
rect 150114 273922 150170 273978
rect 155814 274294 155870 274350
rect 155938 274294 155994 274350
rect 155814 274170 155870 274226
rect 155938 274170 155994 274226
rect 155814 274046 155870 274102
rect 155938 274046 155994 274102
rect 155814 273922 155870 273978
rect 155938 273922 155994 273978
rect 161638 274294 161694 274350
rect 161762 274294 161818 274350
rect 161638 274170 161694 274226
rect 161762 274170 161818 274226
rect 161638 274046 161694 274102
rect 161762 274046 161818 274102
rect 161638 273922 161694 273978
rect 161762 273922 161818 273978
rect 153692 267002 153748 267058
rect 153804 270602 153860 270658
rect 168028 340082 168084 340138
rect 168028 322442 168084 322498
rect 168364 320822 168420 320878
rect 168252 320642 168308 320698
rect 168140 320462 168196 320518
rect 153804 265382 153860 265438
rect 132114 262294 132170 262350
rect 132238 262294 132294 262350
rect 132362 262294 132418 262350
rect 132486 262294 132542 262350
rect 132114 262170 132170 262226
rect 132238 262170 132294 262226
rect 132362 262170 132418 262226
rect 132486 262170 132542 262226
rect 132114 262046 132170 262102
rect 132238 262046 132294 262102
rect 132362 262046 132418 262102
rect 132486 262046 132542 262102
rect 132114 261922 132170 261978
rect 132238 261922 132294 261978
rect 132362 261922 132418 261978
rect 132486 261922 132542 261978
rect 168812 267002 168868 267058
rect 162834 262294 162890 262350
rect 162958 262294 163014 262350
rect 163082 262294 163138 262350
rect 163206 262294 163262 262350
rect 162834 262170 162890 262226
rect 162958 262170 163014 262226
rect 163082 262170 163138 262226
rect 163206 262170 163262 262226
rect 162834 262046 162890 262102
rect 162958 262046 163014 262102
rect 163082 262046 163138 262102
rect 163206 262046 163262 262102
rect 162834 261922 162890 261978
rect 162958 261922 163014 261978
rect 163082 261922 163138 261978
rect 163206 261922 163262 261978
rect 132114 244294 132170 244350
rect 132238 244294 132294 244350
rect 132362 244294 132418 244350
rect 132486 244294 132542 244350
rect 132114 244170 132170 244226
rect 132238 244170 132294 244226
rect 132362 244170 132418 244226
rect 132486 244170 132542 244226
rect 132114 244046 132170 244102
rect 132238 244046 132294 244102
rect 132362 244046 132418 244102
rect 132486 244046 132542 244102
rect 132114 243922 132170 243978
rect 132238 243922 132294 243978
rect 132362 243922 132418 243978
rect 132486 243922 132542 243978
rect 132114 226294 132170 226350
rect 132238 226294 132294 226350
rect 132362 226294 132418 226350
rect 132486 226294 132542 226350
rect 132114 226170 132170 226226
rect 132238 226170 132294 226226
rect 132362 226170 132418 226226
rect 132486 226170 132542 226226
rect 132114 226046 132170 226102
rect 132238 226046 132294 226102
rect 132362 226046 132418 226102
rect 132486 226046 132542 226102
rect 132114 225922 132170 225978
rect 132238 225922 132294 225978
rect 132362 225922 132418 225978
rect 132486 225922 132542 225978
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 170492 237662 170548 237718
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 177996 270602 178052 270658
rect 174636 251162 174692 251218
rect 182924 402362 182980 402418
rect 184604 403982 184660 404038
rect 184716 403262 184772 403318
rect 186284 402542 186340 402598
rect 186396 381302 186452 381358
rect 184492 210842 184548 210898
rect 187068 288782 187124 288838
rect 187068 285722 187124 285778
rect 187852 407762 187908 407818
rect 187740 407582 187796 407638
rect 189834 562294 189890 562350
rect 189958 562294 190014 562350
rect 190082 562294 190138 562350
rect 190206 562294 190262 562350
rect 189834 562170 189890 562226
rect 189958 562170 190014 562226
rect 190082 562170 190138 562226
rect 190206 562170 190262 562226
rect 189834 562046 189890 562102
rect 189958 562046 190014 562102
rect 190082 562046 190138 562102
rect 190206 562046 190262 562102
rect 189834 561922 189890 561978
rect 189958 561922 190014 561978
rect 190082 561922 190138 561978
rect 190206 561922 190262 561978
rect 189834 544294 189890 544350
rect 189958 544294 190014 544350
rect 190082 544294 190138 544350
rect 190206 544294 190262 544350
rect 189834 544170 189890 544226
rect 189958 544170 190014 544226
rect 190082 544170 190138 544226
rect 190206 544170 190262 544226
rect 189834 544046 189890 544102
rect 189958 544046 190014 544102
rect 190082 544046 190138 544102
rect 190206 544046 190262 544102
rect 189834 543922 189890 543978
rect 189958 543922 190014 543978
rect 190082 543922 190138 543978
rect 190206 543922 190262 543978
rect 189834 526294 189890 526350
rect 189958 526294 190014 526350
rect 190082 526294 190138 526350
rect 190206 526294 190262 526350
rect 189834 526170 189890 526226
rect 189958 526170 190014 526226
rect 190082 526170 190138 526226
rect 190206 526170 190262 526226
rect 189834 526046 189890 526102
rect 189958 526046 190014 526102
rect 190082 526046 190138 526102
rect 190206 526046 190262 526102
rect 189834 525922 189890 525978
rect 189958 525922 190014 525978
rect 190082 525922 190138 525978
rect 190206 525922 190262 525978
rect 187964 397322 188020 397378
rect 189532 390662 189588 390718
rect 189834 508294 189890 508350
rect 189958 508294 190014 508350
rect 190082 508294 190138 508350
rect 190206 508294 190262 508350
rect 189834 508170 189890 508226
rect 189958 508170 190014 508226
rect 190082 508170 190138 508226
rect 190206 508170 190262 508226
rect 189834 508046 189890 508102
rect 189958 508046 190014 508102
rect 190082 508046 190138 508102
rect 190206 508046 190262 508102
rect 189834 507922 189890 507978
rect 189958 507922 190014 507978
rect 190082 507922 190138 507978
rect 190206 507922 190262 507978
rect 189834 490294 189890 490350
rect 189958 490294 190014 490350
rect 190082 490294 190138 490350
rect 190206 490294 190262 490350
rect 189834 490170 189890 490226
rect 189958 490170 190014 490226
rect 190082 490170 190138 490226
rect 190206 490170 190262 490226
rect 189834 490046 189890 490102
rect 189958 490046 190014 490102
rect 190082 490046 190138 490102
rect 190206 490046 190262 490102
rect 189834 489922 189890 489978
rect 189958 489922 190014 489978
rect 190082 489922 190138 489978
rect 190206 489922 190262 489978
rect 189834 472294 189890 472350
rect 189958 472294 190014 472350
rect 190082 472294 190138 472350
rect 190206 472294 190262 472350
rect 189834 472170 189890 472226
rect 189958 472170 190014 472226
rect 190082 472170 190138 472226
rect 190206 472170 190262 472226
rect 189834 472046 189890 472102
rect 189958 472046 190014 472102
rect 190082 472046 190138 472102
rect 190206 472046 190262 472102
rect 189834 471922 189890 471978
rect 189958 471922 190014 471978
rect 190082 471922 190138 471978
rect 190206 471922 190262 471978
rect 189834 454294 189890 454350
rect 189958 454294 190014 454350
rect 190082 454294 190138 454350
rect 190206 454294 190262 454350
rect 189834 454170 189890 454226
rect 189958 454170 190014 454226
rect 190082 454170 190138 454226
rect 190206 454170 190262 454226
rect 189834 454046 189890 454102
rect 189958 454046 190014 454102
rect 190082 454046 190138 454102
rect 190206 454046 190262 454102
rect 189834 453922 189890 453978
rect 189958 453922 190014 453978
rect 190082 453922 190138 453978
rect 190206 453922 190262 453978
rect 189834 436294 189890 436350
rect 189958 436294 190014 436350
rect 190082 436294 190138 436350
rect 190206 436294 190262 436350
rect 189834 436170 189890 436226
rect 189958 436170 190014 436226
rect 190082 436170 190138 436226
rect 190206 436170 190262 436226
rect 189834 436046 189890 436102
rect 189958 436046 190014 436102
rect 190082 436046 190138 436102
rect 190206 436046 190262 436102
rect 189834 435922 189890 435978
rect 189958 435922 190014 435978
rect 190082 435922 190138 435978
rect 190206 435922 190262 435978
rect 189834 418294 189890 418350
rect 189958 418294 190014 418350
rect 190082 418294 190138 418350
rect 190206 418294 190262 418350
rect 189834 418170 189890 418226
rect 189958 418170 190014 418226
rect 190082 418170 190138 418226
rect 190206 418170 190262 418226
rect 189834 418046 189890 418102
rect 189958 418046 190014 418102
rect 190082 418046 190138 418102
rect 190206 418046 190262 418102
rect 189834 417922 189890 417978
rect 189958 417922 190014 417978
rect 190082 417922 190138 417978
rect 190206 417922 190262 417978
rect 189834 400294 189890 400350
rect 189958 400294 190014 400350
rect 190082 400294 190138 400350
rect 190206 400294 190262 400350
rect 189834 400170 189890 400226
rect 189958 400170 190014 400226
rect 190082 400170 190138 400226
rect 190206 400170 190262 400226
rect 189834 400046 189890 400102
rect 189958 400046 190014 400102
rect 190082 400046 190138 400102
rect 190206 400046 190262 400102
rect 189834 399922 189890 399978
rect 189958 399922 190014 399978
rect 190082 399922 190138 399978
rect 190206 399922 190262 399978
rect 189834 382294 189890 382350
rect 189958 382294 190014 382350
rect 190082 382294 190138 382350
rect 190206 382294 190262 382350
rect 189834 382170 189890 382226
rect 189958 382170 190014 382226
rect 190082 382170 190138 382226
rect 190206 382170 190262 382226
rect 189834 382046 189890 382102
rect 189958 382046 190014 382102
rect 190082 382046 190138 382102
rect 190206 382046 190262 382102
rect 189834 381922 189890 381978
rect 189958 381922 190014 381978
rect 190082 381922 190138 381978
rect 190206 381922 190262 381978
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 193554 568294 193610 568350
rect 193678 568294 193734 568350
rect 193802 568294 193858 568350
rect 193926 568294 193982 568350
rect 193554 568170 193610 568226
rect 193678 568170 193734 568226
rect 193802 568170 193858 568226
rect 193926 568170 193982 568226
rect 193554 568046 193610 568102
rect 193678 568046 193734 568102
rect 193802 568046 193858 568102
rect 193926 568046 193982 568102
rect 193554 567922 193610 567978
rect 193678 567922 193734 567978
rect 193802 567922 193858 567978
rect 193926 567922 193982 567978
rect 194518 562294 194574 562350
rect 194642 562294 194698 562350
rect 194518 562170 194574 562226
rect 194642 562170 194698 562226
rect 194518 562046 194574 562102
rect 194642 562046 194698 562102
rect 194518 561922 194574 561978
rect 194642 561922 194698 561978
rect 193554 550294 193610 550350
rect 193678 550294 193734 550350
rect 193802 550294 193858 550350
rect 193926 550294 193982 550350
rect 193554 550170 193610 550226
rect 193678 550170 193734 550226
rect 193802 550170 193858 550226
rect 193926 550170 193982 550226
rect 193554 550046 193610 550102
rect 193678 550046 193734 550102
rect 193802 550046 193858 550102
rect 193926 550046 193982 550102
rect 193554 549922 193610 549978
rect 193678 549922 193734 549978
rect 193802 549922 193858 549978
rect 193926 549922 193982 549978
rect 194518 544294 194574 544350
rect 194642 544294 194698 544350
rect 194518 544170 194574 544226
rect 194642 544170 194698 544226
rect 194518 544046 194574 544102
rect 194642 544046 194698 544102
rect 194518 543922 194574 543978
rect 194642 543922 194698 543978
rect 193554 532294 193610 532350
rect 193678 532294 193734 532350
rect 193802 532294 193858 532350
rect 193926 532294 193982 532350
rect 193554 532170 193610 532226
rect 193678 532170 193734 532226
rect 193802 532170 193858 532226
rect 193926 532170 193982 532226
rect 193554 532046 193610 532102
rect 193678 532046 193734 532102
rect 193802 532046 193858 532102
rect 193926 532046 193982 532102
rect 193554 531922 193610 531978
rect 193678 531922 193734 531978
rect 193802 531922 193858 531978
rect 193926 531922 193982 531978
rect 194518 526294 194574 526350
rect 194642 526294 194698 526350
rect 194518 526170 194574 526226
rect 194642 526170 194698 526226
rect 194518 526046 194574 526102
rect 194642 526046 194698 526102
rect 194518 525922 194574 525978
rect 194642 525922 194698 525978
rect 193554 514294 193610 514350
rect 193678 514294 193734 514350
rect 193802 514294 193858 514350
rect 193926 514294 193982 514350
rect 193554 514170 193610 514226
rect 193678 514170 193734 514226
rect 193802 514170 193858 514226
rect 193926 514170 193982 514226
rect 193554 514046 193610 514102
rect 193678 514046 193734 514102
rect 193802 514046 193858 514102
rect 193926 514046 193982 514102
rect 193554 513922 193610 513978
rect 193678 513922 193734 513978
rect 193802 513922 193858 513978
rect 193926 513922 193982 513978
rect 194518 508294 194574 508350
rect 194642 508294 194698 508350
rect 194518 508170 194574 508226
rect 194642 508170 194698 508226
rect 194518 508046 194574 508102
rect 194642 508046 194698 508102
rect 194518 507922 194574 507978
rect 194642 507922 194698 507978
rect 193554 496294 193610 496350
rect 193678 496294 193734 496350
rect 193802 496294 193858 496350
rect 193926 496294 193982 496350
rect 193554 496170 193610 496226
rect 193678 496170 193734 496226
rect 193802 496170 193858 496226
rect 193926 496170 193982 496226
rect 193554 496046 193610 496102
rect 193678 496046 193734 496102
rect 193802 496046 193858 496102
rect 193926 496046 193982 496102
rect 193554 495922 193610 495978
rect 193678 495922 193734 495978
rect 193802 495922 193858 495978
rect 193926 495922 193982 495978
rect 194518 490294 194574 490350
rect 194642 490294 194698 490350
rect 194518 490170 194574 490226
rect 194642 490170 194698 490226
rect 194518 490046 194574 490102
rect 194642 490046 194698 490102
rect 194518 489922 194574 489978
rect 194642 489922 194698 489978
rect 193554 478294 193610 478350
rect 193678 478294 193734 478350
rect 193802 478294 193858 478350
rect 193926 478294 193982 478350
rect 193554 478170 193610 478226
rect 193678 478170 193734 478226
rect 193802 478170 193858 478226
rect 193926 478170 193982 478226
rect 193554 478046 193610 478102
rect 193678 478046 193734 478102
rect 193802 478046 193858 478102
rect 193926 478046 193982 478102
rect 193554 477922 193610 477978
rect 193678 477922 193734 477978
rect 193802 477922 193858 477978
rect 193926 477922 193982 477978
rect 194518 472294 194574 472350
rect 194642 472294 194698 472350
rect 194518 472170 194574 472226
rect 194642 472170 194698 472226
rect 194518 472046 194574 472102
rect 194642 472046 194698 472102
rect 194518 471922 194574 471978
rect 194642 471922 194698 471978
rect 193554 460294 193610 460350
rect 193678 460294 193734 460350
rect 193802 460294 193858 460350
rect 193926 460294 193982 460350
rect 193554 460170 193610 460226
rect 193678 460170 193734 460226
rect 193802 460170 193858 460226
rect 193926 460170 193982 460226
rect 193554 460046 193610 460102
rect 193678 460046 193734 460102
rect 193802 460046 193858 460102
rect 193926 460046 193982 460102
rect 193554 459922 193610 459978
rect 193678 459922 193734 459978
rect 193802 459922 193858 459978
rect 193926 459922 193982 459978
rect 194518 454294 194574 454350
rect 194642 454294 194698 454350
rect 194518 454170 194574 454226
rect 194642 454170 194698 454226
rect 194518 454046 194574 454102
rect 194642 454046 194698 454102
rect 194518 453922 194574 453978
rect 194642 453922 194698 453978
rect 193554 442294 193610 442350
rect 193678 442294 193734 442350
rect 193802 442294 193858 442350
rect 193926 442294 193982 442350
rect 193554 442170 193610 442226
rect 193678 442170 193734 442226
rect 193802 442170 193858 442226
rect 193926 442170 193982 442226
rect 193554 442046 193610 442102
rect 193678 442046 193734 442102
rect 193802 442046 193858 442102
rect 193926 442046 193982 442102
rect 193554 441922 193610 441978
rect 193678 441922 193734 441978
rect 193802 441922 193858 441978
rect 193926 441922 193982 441978
rect 194518 436294 194574 436350
rect 194642 436294 194698 436350
rect 194518 436170 194574 436226
rect 194642 436170 194698 436226
rect 194518 436046 194574 436102
rect 194642 436046 194698 436102
rect 194518 435922 194574 435978
rect 194642 435922 194698 435978
rect 193554 424294 193610 424350
rect 193678 424294 193734 424350
rect 193802 424294 193858 424350
rect 193926 424294 193982 424350
rect 193554 424170 193610 424226
rect 193678 424170 193734 424226
rect 193802 424170 193858 424226
rect 193926 424170 193982 424226
rect 193554 424046 193610 424102
rect 193678 424046 193734 424102
rect 193802 424046 193858 424102
rect 193926 424046 193982 424102
rect 193554 423922 193610 423978
rect 193678 423922 193734 423978
rect 193802 423922 193858 423978
rect 193926 423922 193982 423978
rect 194518 418294 194574 418350
rect 194642 418294 194698 418350
rect 194518 418170 194574 418226
rect 194642 418170 194698 418226
rect 194518 418046 194574 418102
rect 194642 418046 194698 418102
rect 194518 417922 194574 417978
rect 194642 417922 194698 417978
rect 193554 406294 193610 406350
rect 193678 406294 193734 406350
rect 193802 406294 193858 406350
rect 193926 406294 193982 406350
rect 193554 406170 193610 406226
rect 193678 406170 193734 406226
rect 193802 406170 193858 406226
rect 193926 406170 193982 406226
rect 193554 406046 193610 406102
rect 193678 406046 193734 406102
rect 193802 406046 193858 406102
rect 193926 406046 193982 406102
rect 193554 405922 193610 405978
rect 193678 405922 193734 405978
rect 193802 405922 193858 405978
rect 193926 405922 193982 405978
rect 193554 388294 193610 388350
rect 193678 388294 193734 388350
rect 193802 388294 193858 388350
rect 193926 388294 193982 388350
rect 193554 388170 193610 388226
rect 193678 388170 193734 388226
rect 193802 388170 193858 388226
rect 193926 388170 193982 388226
rect 193554 388046 193610 388102
rect 193678 388046 193734 388102
rect 193802 388046 193858 388102
rect 193926 388046 193982 388102
rect 193554 387922 193610 387978
rect 193678 387922 193734 387978
rect 193802 387922 193858 387978
rect 193926 387922 193982 387978
rect 201404 401642 201460 401698
rect 203196 393722 203252 393778
rect 203084 393362 203140 393418
rect 204764 393902 204820 393958
rect 204876 393182 204932 393238
rect 206444 398222 206500 398278
rect 206556 393542 206612 393598
rect 193554 370294 193610 370350
rect 193678 370294 193734 370350
rect 193802 370294 193858 370350
rect 193926 370294 193982 370350
rect 193554 370170 193610 370226
rect 193678 370170 193734 370226
rect 193802 370170 193858 370226
rect 193926 370170 193982 370226
rect 193554 370046 193610 370102
rect 193678 370046 193734 370102
rect 193802 370046 193858 370102
rect 193926 370046 193982 370102
rect 193554 369922 193610 369978
rect 193678 369922 193734 369978
rect 193802 369922 193858 369978
rect 193926 369922 193982 369978
rect 190652 367982 190708 368038
rect 190652 366542 190708 366598
rect 190652 366380 190708 366418
rect 190652 366362 190708 366380
rect 190652 364588 190708 364618
rect 190652 364562 190708 364588
rect 189834 364294 189890 364350
rect 189958 364294 190014 364350
rect 190082 364294 190138 364350
rect 190206 364294 190262 364350
rect 189834 364170 189890 364226
rect 189958 364170 190014 364226
rect 190082 364170 190138 364226
rect 190206 364170 190262 364226
rect 189834 364046 189890 364102
rect 189958 364046 190014 364102
rect 190082 364046 190138 364102
rect 190206 364046 190262 364102
rect 189834 363922 189890 363978
rect 189958 363922 190014 363978
rect 190082 363922 190138 363978
rect 190206 363922 190262 363978
rect 189834 346294 189890 346350
rect 189958 346294 190014 346350
rect 190082 346294 190138 346350
rect 190206 346294 190262 346350
rect 189834 346170 189890 346226
rect 189958 346170 190014 346226
rect 190082 346170 190138 346226
rect 190206 346170 190262 346226
rect 189834 346046 189890 346102
rect 189958 346046 190014 346102
rect 190082 346046 190138 346102
rect 190206 346046 190262 346102
rect 189834 345922 189890 345978
rect 189958 345922 190014 345978
rect 190082 345922 190138 345978
rect 190206 345922 190262 345978
rect 189834 328294 189890 328350
rect 189958 328294 190014 328350
rect 190082 328294 190138 328350
rect 190206 328294 190262 328350
rect 189834 328170 189890 328226
rect 189958 328170 190014 328226
rect 190082 328170 190138 328226
rect 190206 328170 190262 328226
rect 189834 328046 189890 328102
rect 189958 328046 190014 328102
rect 190082 328046 190138 328102
rect 190206 328046 190262 328102
rect 189834 327922 189890 327978
rect 189958 327922 190014 327978
rect 190082 327922 190138 327978
rect 190206 327922 190262 327978
rect 194518 364294 194574 364350
rect 194642 364294 194698 364350
rect 194518 364170 194574 364226
rect 194642 364170 194698 364226
rect 194518 364046 194574 364102
rect 194642 364046 194698 364102
rect 194518 363922 194574 363978
rect 194642 363922 194698 363978
rect 193554 352294 193610 352350
rect 193678 352294 193734 352350
rect 193802 352294 193858 352350
rect 193926 352294 193982 352350
rect 193554 352170 193610 352226
rect 193678 352170 193734 352226
rect 193802 352170 193858 352226
rect 193926 352170 193982 352226
rect 193554 352046 193610 352102
rect 193678 352046 193734 352102
rect 193802 352046 193858 352102
rect 193926 352046 193982 352102
rect 193554 351922 193610 351978
rect 193678 351922 193734 351978
rect 193802 351922 193858 351978
rect 193926 351922 193982 351978
rect 194518 346294 194574 346350
rect 194642 346294 194698 346350
rect 194518 346170 194574 346226
rect 194642 346170 194698 346226
rect 194518 346046 194574 346102
rect 194642 346046 194698 346102
rect 194518 345922 194574 345978
rect 194642 345922 194698 345978
rect 193554 334294 193610 334350
rect 193678 334294 193734 334350
rect 193802 334294 193858 334350
rect 193926 334294 193982 334350
rect 193554 334170 193610 334226
rect 193678 334170 193734 334226
rect 193802 334170 193858 334226
rect 193926 334170 193982 334226
rect 193554 334046 193610 334102
rect 193678 334046 193734 334102
rect 193802 334046 193858 334102
rect 193926 334046 193982 334102
rect 193554 333922 193610 333978
rect 193678 333922 193734 333978
rect 193802 333922 193858 333978
rect 193926 333922 193982 333978
rect 190652 319202 190708 319258
rect 194518 328294 194574 328350
rect 194642 328294 194698 328350
rect 194518 328170 194574 328226
rect 194642 328170 194698 328226
rect 194518 328046 194574 328102
rect 194642 328046 194698 328102
rect 194518 327922 194574 327978
rect 194642 327922 194698 327978
rect 193554 316294 193610 316350
rect 193678 316294 193734 316350
rect 193802 316294 193858 316350
rect 193926 316294 193982 316350
rect 193554 316170 193610 316226
rect 193678 316170 193734 316226
rect 193802 316170 193858 316226
rect 193926 316170 193982 316226
rect 193554 316046 193610 316102
rect 193678 316046 193734 316102
rect 193802 316046 193858 316102
rect 193926 316046 193982 316102
rect 193554 315922 193610 315978
rect 193678 315922 193734 315978
rect 193802 315922 193858 315978
rect 193926 315922 193982 315978
rect 189834 310294 189890 310350
rect 189958 310294 190014 310350
rect 190082 310294 190138 310350
rect 190206 310294 190262 310350
rect 189834 310170 189890 310226
rect 189958 310170 190014 310226
rect 190082 310170 190138 310226
rect 190206 310170 190262 310226
rect 189834 310046 189890 310102
rect 189958 310046 190014 310102
rect 190082 310046 190138 310102
rect 190206 310046 190262 310102
rect 189834 309922 189890 309978
rect 189958 309922 190014 309978
rect 190082 309922 190138 309978
rect 190206 309922 190262 309978
rect 188076 288962 188132 289018
rect 188076 287342 188132 287398
rect 188076 285902 188132 285958
rect 188076 283922 188132 283978
rect 188076 270602 188132 270658
rect 189834 292294 189890 292350
rect 189958 292294 190014 292350
rect 190082 292294 190138 292350
rect 190206 292294 190262 292350
rect 189834 292170 189890 292226
rect 189958 292170 190014 292226
rect 190082 292170 190138 292226
rect 190206 292170 190262 292226
rect 189834 292046 189890 292102
rect 189958 292046 190014 292102
rect 190082 292046 190138 292102
rect 190206 292046 190262 292102
rect 189834 291922 189890 291978
rect 189958 291922 190014 291978
rect 190082 291922 190138 291978
rect 190206 291922 190262 291978
rect 189834 274294 189890 274350
rect 189958 274294 190014 274350
rect 190082 274294 190138 274350
rect 190206 274294 190262 274350
rect 189834 274170 189890 274226
rect 189958 274170 190014 274226
rect 190082 274170 190138 274226
rect 190206 274170 190262 274226
rect 189834 274046 189890 274102
rect 189958 274046 190014 274102
rect 190082 274046 190138 274102
rect 190206 274046 190262 274102
rect 189834 273922 189890 273978
rect 189958 273922 190014 273978
rect 190082 273922 190138 273978
rect 190206 273922 190262 273978
rect 189834 256294 189890 256350
rect 189958 256294 190014 256350
rect 190082 256294 190138 256350
rect 190206 256294 190262 256350
rect 189834 256170 189890 256226
rect 189958 256170 190014 256226
rect 190082 256170 190138 256226
rect 190206 256170 190262 256226
rect 189834 256046 189890 256102
rect 189958 256046 190014 256102
rect 190082 256046 190138 256102
rect 190206 256046 190262 256102
rect 189834 255922 189890 255978
rect 189958 255922 190014 255978
rect 190082 255922 190138 255978
rect 190206 255922 190262 255978
rect 189834 238294 189890 238350
rect 189958 238294 190014 238350
rect 190082 238294 190138 238350
rect 190206 238294 190262 238350
rect 189834 238170 189890 238226
rect 189958 238170 190014 238226
rect 190082 238170 190138 238226
rect 190206 238170 190262 238226
rect 189834 238046 189890 238102
rect 189958 238046 190014 238102
rect 190082 238046 190138 238102
rect 190206 238046 190262 238102
rect 189834 237922 189890 237978
rect 189958 237922 190014 237978
rect 190082 237922 190138 237978
rect 190206 237922 190262 237978
rect 194518 310294 194574 310350
rect 194642 310294 194698 310350
rect 194518 310170 194574 310226
rect 194642 310170 194698 310226
rect 194518 310046 194574 310102
rect 194642 310046 194698 310102
rect 194518 309922 194574 309978
rect 194642 309922 194698 309978
rect 193554 298294 193610 298350
rect 193678 298294 193734 298350
rect 193802 298294 193858 298350
rect 193926 298294 193982 298350
rect 193554 298170 193610 298226
rect 193678 298170 193734 298226
rect 193802 298170 193858 298226
rect 193926 298170 193982 298226
rect 193554 298046 193610 298102
rect 193678 298046 193734 298102
rect 193802 298046 193858 298102
rect 193926 298046 193982 298102
rect 193554 297922 193610 297978
rect 193678 297922 193734 297978
rect 193802 297922 193858 297978
rect 193926 297922 193982 297978
rect 190652 292562 190708 292618
rect 194518 292294 194574 292350
rect 194642 292294 194698 292350
rect 194518 292170 194574 292226
rect 194642 292170 194698 292226
rect 194518 292046 194574 292102
rect 194642 292046 194698 292102
rect 194518 291922 194574 291978
rect 194642 291922 194698 291978
rect 193554 280294 193610 280350
rect 193678 280294 193734 280350
rect 193802 280294 193858 280350
rect 193926 280294 193982 280350
rect 193554 280170 193610 280226
rect 193678 280170 193734 280226
rect 193802 280170 193858 280226
rect 193926 280170 193982 280226
rect 193554 280046 193610 280102
rect 193678 280046 193734 280102
rect 193802 280046 193858 280102
rect 193926 280046 193982 280102
rect 193554 279922 193610 279978
rect 193678 279922 193734 279978
rect 193802 279922 193858 279978
rect 193926 279922 193982 279978
rect 194518 274294 194574 274350
rect 194642 274294 194698 274350
rect 194518 274170 194574 274226
rect 194642 274170 194698 274226
rect 194518 274046 194574 274102
rect 194642 274046 194698 274102
rect 194518 273922 194574 273978
rect 194642 273922 194698 273978
rect 193554 262294 193610 262350
rect 193678 262294 193734 262350
rect 193802 262294 193858 262350
rect 193926 262294 193982 262350
rect 193554 262170 193610 262226
rect 193678 262170 193734 262226
rect 193802 262170 193858 262226
rect 193926 262170 193982 262226
rect 193554 262046 193610 262102
rect 193678 262046 193734 262102
rect 193802 262046 193858 262102
rect 193926 262046 193982 262102
rect 193554 261922 193610 261978
rect 193678 261922 193734 261978
rect 193802 261922 193858 261978
rect 193926 261922 193982 261978
rect 190652 260342 190708 260398
rect 190652 255482 190708 255538
rect 190652 252062 190708 252118
rect 194518 256294 194574 256350
rect 194642 256294 194698 256350
rect 194518 256170 194574 256226
rect 194642 256170 194698 256226
rect 194518 256046 194574 256102
rect 194642 256046 194698 256102
rect 194518 255922 194574 255978
rect 194642 255922 194698 255978
rect 193554 244294 193610 244350
rect 193678 244294 193734 244350
rect 193802 244294 193858 244350
rect 193926 244294 193982 244350
rect 193554 244170 193610 244226
rect 193678 244170 193734 244226
rect 193802 244170 193858 244226
rect 193926 244170 193982 244226
rect 193554 244046 193610 244102
rect 193678 244046 193734 244102
rect 193802 244046 193858 244102
rect 193926 244046 193982 244102
rect 193554 243922 193610 243978
rect 193678 243922 193734 243978
rect 193802 243922 193858 243978
rect 193926 243922 193982 243978
rect 193554 226294 193610 226350
rect 193678 226294 193734 226350
rect 193802 226294 193858 226350
rect 193926 226294 193982 226350
rect 193554 226170 193610 226226
rect 193678 226170 193734 226226
rect 193802 226170 193858 226226
rect 193926 226170 193982 226226
rect 193554 226046 193610 226102
rect 193678 226046 193734 226102
rect 193802 226046 193858 226102
rect 193926 226046 193982 226102
rect 193554 225922 193610 225978
rect 193678 225922 193734 225978
rect 193802 225922 193858 225978
rect 193926 225922 193982 225978
rect 189834 220294 189890 220350
rect 189958 220294 190014 220350
rect 190082 220294 190138 220350
rect 190206 220294 190262 220350
rect 189834 220170 189890 220226
rect 189958 220170 190014 220226
rect 190082 220170 190138 220226
rect 190206 220170 190262 220226
rect 189834 220046 189890 220102
rect 189958 220046 190014 220102
rect 190082 220046 190138 220102
rect 190206 220046 190262 220102
rect 189834 219922 189890 219978
rect 189958 219922 190014 219978
rect 190082 219922 190138 219978
rect 190206 219922 190262 219978
rect 208124 404162 208180 404218
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 224274 568294 224330 568350
rect 224398 568294 224454 568350
rect 224522 568294 224578 568350
rect 224646 568294 224702 568350
rect 224274 568170 224330 568226
rect 224398 568170 224454 568226
rect 224522 568170 224578 568226
rect 224646 568170 224702 568226
rect 224274 568046 224330 568102
rect 224398 568046 224454 568102
rect 224522 568046 224578 568102
rect 224646 568046 224702 568102
rect 224274 567922 224330 567978
rect 224398 567922 224454 567978
rect 224522 567922 224578 567978
rect 224646 567922 224702 567978
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 254994 568294 255050 568350
rect 255118 568294 255174 568350
rect 255242 568294 255298 568350
rect 255366 568294 255422 568350
rect 254994 568170 255050 568226
rect 255118 568170 255174 568226
rect 255242 568170 255298 568226
rect 255366 568170 255422 568226
rect 254994 568046 255050 568102
rect 255118 568046 255174 568102
rect 255242 568046 255298 568102
rect 255366 568046 255422 568102
rect 254994 567922 255050 567978
rect 255118 567922 255174 567978
rect 255242 567922 255298 567978
rect 255366 567922 255422 567978
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 285714 568294 285770 568350
rect 285838 568294 285894 568350
rect 285962 568294 286018 568350
rect 286086 568294 286142 568350
rect 285714 568170 285770 568226
rect 285838 568170 285894 568226
rect 285962 568170 286018 568226
rect 286086 568170 286142 568226
rect 285714 568046 285770 568102
rect 285838 568046 285894 568102
rect 285962 568046 286018 568102
rect 286086 568046 286142 568102
rect 285714 567922 285770 567978
rect 285838 567922 285894 567978
rect 285962 567922 286018 567978
rect 286086 567922 286142 567978
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 316434 568294 316490 568350
rect 316558 568294 316614 568350
rect 316682 568294 316738 568350
rect 316806 568294 316862 568350
rect 316434 568170 316490 568226
rect 316558 568170 316614 568226
rect 316682 568170 316738 568226
rect 316806 568170 316862 568226
rect 316434 568046 316490 568102
rect 316558 568046 316614 568102
rect 316682 568046 316738 568102
rect 316806 568046 316862 568102
rect 316434 567922 316490 567978
rect 316558 567922 316614 567978
rect 316682 567922 316738 567978
rect 316806 567922 316862 567978
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 347154 568294 347210 568350
rect 347278 568294 347334 568350
rect 347402 568294 347458 568350
rect 347526 568294 347582 568350
rect 347154 568170 347210 568226
rect 347278 568170 347334 568226
rect 347402 568170 347458 568226
rect 347526 568170 347582 568226
rect 347154 568046 347210 568102
rect 347278 568046 347334 568102
rect 347402 568046 347458 568102
rect 347526 568046 347582 568102
rect 347154 567922 347210 567978
rect 347278 567922 347334 567978
rect 347402 567922 347458 567978
rect 347526 567922 347582 567978
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 377874 568294 377930 568350
rect 377998 568294 378054 568350
rect 378122 568294 378178 568350
rect 378246 568294 378302 568350
rect 377874 568170 377930 568226
rect 377998 568170 378054 568226
rect 378122 568170 378178 568226
rect 378246 568170 378302 568226
rect 377874 568046 377930 568102
rect 377998 568046 378054 568102
rect 378122 568046 378178 568102
rect 378246 568046 378302 568102
rect 377874 567922 377930 567978
rect 377998 567922 378054 567978
rect 378122 567922 378178 567978
rect 378246 567922 378302 567978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 408594 568294 408650 568350
rect 408718 568294 408774 568350
rect 408842 568294 408898 568350
rect 408966 568294 409022 568350
rect 408594 568170 408650 568226
rect 408718 568170 408774 568226
rect 408842 568170 408898 568226
rect 408966 568170 409022 568226
rect 408594 568046 408650 568102
rect 408718 568046 408774 568102
rect 408842 568046 408898 568102
rect 408966 568046 409022 568102
rect 408594 567922 408650 567978
rect 408718 567922 408774 567978
rect 408842 567922 408898 567978
rect 408966 567922 409022 567978
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 439314 568294 439370 568350
rect 439438 568294 439494 568350
rect 439562 568294 439618 568350
rect 439686 568294 439742 568350
rect 439314 568170 439370 568226
rect 439438 568170 439494 568226
rect 439562 568170 439618 568226
rect 439686 568170 439742 568226
rect 439314 568046 439370 568102
rect 439438 568046 439494 568102
rect 439562 568046 439618 568102
rect 439686 568046 439742 568102
rect 439314 567922 439370 567978
rect 439438 567922 439494 567978
rect 439562 567922 439618 567978
rect 439686 567922 439742 567978
rect 225238 562294 225294 562350
rect 225362 562294 225418 562350
rect 225238 562170 225294 562226
rect 225362 562170 225418 562226
rect 225238 562046 225294 562102
rect 225362 562046 225418 562102
rect 225238 561922 225294 561978
rect 225362 561922 225418 561978
rect 255958 562294 256014 562350
rect 256082 562294 256138 562350
rect 255958 562170 256014 562226
rect 256082 562170 256138 562226
rect 255958 562046 256014 562102
rect 256082 562046 256138 562102
rect 255958 561922 256014 561978
rect 256082 561922 256138 561978
rect 286678 562294 286734 562350
rect 286802 562294 286858 562350
rect 286678 562170 286734 562226
rect 286802 562170 286858 562226
rect 286678 562046 286734 562102
rect 286802 562046 286858 562102
rect 286678 561922 286734 561978
rect 286802 561922 286858 561978
rect 317398 562294 317454 562350
rect 317522 562294 317578 562350
rect 317398 562170 317454 562226
rect 317522 562170 317578 562226
rect 317398 562046 317454 562102
rect 317522 562046 317578 562102
rect 317398 561922 317454 561978
rect 317522 561922 317578 561978
rect 348118 562294 348174 562350
rect 348242 562294 348298 562350
rect 348118 562170 348174 562226
rect 348242 562170 348298 562226
rect 348118 562046 348174 562102
rect 348242 562046 348298 562102
rect 348118 561922 348174 561978
rect 348242 561922 348298 561978
rect 378838 562294 378894 562350
rect 378962 562294 379018 562350
rect 378838 562170 378894 562226
rect 378962 562170 379018 562226
rect 378838 562046 378894 562102
rect 378962 562046 379018 562102
rect 378838 561922 378894 561978
rect 378962 561922 379018 561978
rect 409558 562294 409614 562350
rect 409682 562294 409738 562350
rect 409558 562170 409614 562226
rect 409682 562170 409738 562226
rect 409558 562046 409614 562102
rect 409682 562046 409738 562102
rect 409558 561922 409614 561978
rect 409682 561922 409738 561978
rect 440278 562294 440334 562350
rect 440402 562294 440458 562350
rect 440278 562170 440334 562226
rect 440402 562170 440458 562226
rect 440278 562046 440334 562102
rect 440402 562046 440458 562102
rect 440278 561922 440334 561978
rect 440402 561922 440458 561978
rect 209878 550294 209934 550350
rect 210002 550294 210058 550350
rect 209878 550170 209934 550226
rect 210002 550170 210058 550226
rect 209878 550046 209934 550102
rect 210002 550046 210058 550102
rect 209878 549922 209934 549978
rect 210002 549922 210058 549978
rect 240598 550294 240654 550350
rect 240722 550294 240778 550350
rect 240598 550170 240654 550226
rect 240722 550170 240778 550226
rect 240598 550046 240654 550102
rect 240722 550046 240778 550102
rect 240598 549922 240654 549978
rect 240722 549922 240778 549978
rect 271318 550294 271374 550350
rect 271442 550294 271498 550350
rect 271318 550170 271374 550226
rect 271442 550170 271498 550226
rect 271318 550046 271374 550102
rect 271442 550046 271498 550102
rect 271318 549922 271374 549978
rect 271442 549922 271498 549978
rect 302038 550294 302094 550350
rect 302162 550294 302218 550350
rect 302038 550170 302094 550226
rect 302162 550170 302218 550226
rect 302038 550046 302094 550102
rect 302162 550046 302218 550102
rect 302038 549922 302094 549978
rect 302162 549922 302218 549978
rect 332758 550294 332814 550350
rect 332882 550294 332938 550350
rect 332758 550170 332814 550226
rect 332882 550170 332938 550226
rect 332758 550046 332814 550102
rect 332882 550046 332938 550102
rect 332758 549922 332814 549978
rect 332882 549922 332938 549978
rect 363478 550294 363534 550350
rect 363602 550294 363658 550350
rect 363478 550170 363534 550226
rect 363602 550170 363658 550226
rect 363478 550046 363534 550102
rect 363602 550046 363658 550102
rect 363478 549922 363534 549978
rect 363602 549922 363658 549978
rect 394198 550294 394254 550350
rect 394322 550294 394378 550350
rect 394198 550170 394254 550226
rect 394322 550170 394378 550226
rect 394198 550046 394254 550102
rect 394322 550046 394378 550102
rect 394198 549922 394254 549978
rect 394322 549922 394378 549978
rect 424918 550294 424974 550350
rect 425042 550294 425098 550350
rect 424918 550170 424974 550226
rect 425042 550170 425098 550226
rect 424918 550046 424974 550102
rect 425042 550046 425098 550102
rect 424918 549922 424974 549978
rect 425042 549922 425098 549978
rect 225238 544294 225294 544350
rect 225362 544294 225418 544350
rect 225238 544170 225294 544226
rect 225362 544170 225418 544226
rect 225238 544046 225294 544102
rect 225362 544046 225418 544102
rect 225238 543922 225294 543978
rect 225362 543922 225418 543978
rect 255958 544294 256014 544350
rect 256082 544294 256138 544350
rect 255958 544170 256014 544226
rect 256082 544170 256138 544226
rect 255958 544046 256014 544102
rect 256082 544046 256138 544102
rect 255958 543922 256014 543978
rect 256082 543922 256138 543978
rect 286678 544294 286734 544350
rect 286802 544294 286858 544350
rect 286678 544170 286734 544226
rect 286802 544170 286858 544226
rect 286678 544046 286734 544102
rect 286802 544046 286858 544102
rect 286678 543922 286734 543978
rect 286802 543922 286858 543978
rect 317398 544294 317454 544350
rect 317522 544294 317578 544350
rect 317398 544170 317454 544226
rect 317522 544170 317578 544226
rect 317398 544046 317454 544102
rect 317522 544046 317578 544102
rect 317398 543922 317454 543978
rect 317522 543922 317578 543978
rect 348118 544294 348174 544350
rect 348242 544294 348298 544350
rect 348118 544170 348174 544226
rect 348242 544170 348298 544226
rect 348118 544046 348174 544102
rect 348242 544046 348298 544102
rect 348118 543922 348174 543978
rect 348242 543922 348298 543978
rect 378838 544294 378894 544350
rect 378962 544294 379018 544350
rect 378838 544170 378894 544226
rect 378962 544170 379018 544226
rect 378838 544046 378894 544102
rect 378962 544046 379018 544102
rect 378838 543922 378894 543978
rect 378962 543922 379018 543978
rect 409558 544294 409614 544350
rect 409682 544294 409738 544350
rect 409558 544170 409614 544226
rect 409682 544170 409738 544226
rect 409558 544046 409614 544102
rect 409682 544046 409738 544102
rect 409558 543922 409614 543978
rect 409682 543922 409738 543978
rect 440278 544294 440334 544350
rect 440402 544294 440458 544350
rect 440278 544170 440334 544226
rect 440402 544170 440458 544226
rect 440278 544046 440334 544102
rect 440402 544046 440458 544102
rect 440278 543922 440334 543978
rect 440402 543922 440458 543978
rect 209878 532294 209934 532350
rect 210002 532294 210058 532350
rect 209878 532170 209934 532226
rect 210002 532170 210058 532226
rect 209878 532046 209934 532102
rect 210002 532046 210058 532102
rect 209878 531922 209934 531978
rect 210002 531922 210058 531978
rect 240598 532294 240654 532350
rect 240722 532294 240778 532350
rect 240598 532170 240654 532226
rect 240722 532170 240778 532226
rect 240598 532046 240654 532102
rect 240722 532046 240778 532102
rect 240598 531922 240654 531978
rect 240722 531922 240778 531978
rect 271318 532294 271374 532350
rect 271442 532294 271498 532350
rect 271318 532170 271374 532226
rect 271442 532170 271498 532226
rect 271318 532046 271374 532102
rect 271442 532046 271498 532102
rect 271318 531922 271374 531978
rect 271442 531922 271498 531978
rect 302038 532294 302094 532350
rect 302162 532294 302218 532350
rect 302038 532170 302094 532226
rect 302162 532170 302218 532226
rect 302038 532046 302094 532102
rect 302162 532046 302218 532102
rect 302038 531922 302094 531978
rect 302162 531922 302218 531978
rect 332758 532294 332814 532350
rect 332882 532294 332938 532350
rect 332758 532170 332814 532226
rect 332882 532170 332938 532226
rect 332758 532046 332814 532102
rect 332882 532046 332938 532102
rect 332758 531922 332814 531978
rect 332882 531922 332938 531978
rect 363478 532294 363534 532350
rect 363602 532294 363658 532350
rect 363478 532170 363534 532226
rect 363602 532170 363658 532226
rect 363478 532046 363534 532102
rect 363602 532046 363658 532102
rect 363478 531922 363534 531978
rect 363602 531922 363658 531978
rect 394198 532294 394254 532350
rect 394322 532294 394378 532350
rect 394198 532170 394254 532226
rect 394322 532170 394378 532226
rect 394198 532046 394254 532102
rect 394322 532046 394378 532102
rect 394198 531922 394254 531978
rect 394322 531922 394378 531978
rect 424918 532294 424974 532350
rect 425042 532294 425098 532350
rect 424918 532170 424974 532226
rect 425042 532170 425098 532226
rect 424918 532046 424974 532102
rect 425042 532046 425098 532102
rect 424918 531922 424974 531978
rect 425042 531922 425098 531978
rect 225238 526294 225294 526350
rect 225362 526294 225418 526350
rect 225238 526170 225294 526226
rect 225362 526170 225418 526226
rect 225238 526046 225294 526102
rect 225362 526046 225418 526102
rect 225238 525922 225294 525978
rect 225362 525922 225418 525978
rect 255958 526294 256014 526350
rect 256082 526294 256138 526350
rect 255958 526170 256014 526226
rect 256082 526170 256138 526226
rect 255958 526046 256014 526102
rect 256082 526046 256138 526102
rect 255958 525922 256014 525978
rect 256082 525922 256138 525978
rect 286678 526294 286734 526350
rect 286802 526294 286858 526350
rect 286678 526170 286734 526226
rect 286802 526170 286858 526226
rect 286678 526046 286734 526102
rect 286802 526046 286858 526102
rect 286678 525922 286734 525978
rect 286802 525922 286858 525978
rect 317398 526294 317454 526350
rect 317522 526294 317578 526350
rect 317398 526170 317454 526226
rect 317522 526170 317578 526226
rect 317398 526046 317454 526102
rect 317522 526046 317578 526102
rect 317398 525922 317454 525978
rect 317522 525922 317578 525978
rect 348118 526294 348174 526350
rect 348242 526294 348298 526350
rect 348118 526170 348174 526226
rect 348242 526170 348298 526226
rect 348118 526046 348174 526102
rect 348242 526046 348298 526102
rect 348118 525922 348174 525978
rect 348242 525922 348298 525978
rect 378838 526294 378894 526350
rect 378962 526294 379018 526350
rect 378838 526170 378894 526226
rect 378962 526170 379018 526226
rect 378838 526046 378894 526102
rect 378962 526046 379018 526102
rect 378838 525922 378894 525978
rect 378962 525922 379018 525978
rect 409558 526294 409614 526350
rect 409682 526294 409738 526350
rect 409558 526170 409614 526226
rect 409682 526170 409738 526226
rect 409558 526046 409614 526102
rect 409682 526046 409738 526102
rect 409558 525922 409614 525978
rect 409682 525922 409738 525978
rect 440278 526294 440334 526350
rect 440402 526294 440458 526350
rect 440278 526170 440334 526226
rect 440402 526170 440458 526226
rect 440278 526046 440334 526102
rect 440402 526046 440458 526102
rect 440278 525922 440334 525978
rect 440402 525922 440458 525978
rect 209878 514294 209934 514350
rect 210002 514294 210058 514350
rect 209878 514170 209934 514226
rect 210002 514170 210058 514226
rect 209878 514046 209934 514102
rect 210002 514046 210058 514102
rect 209878 513922 209934 513978
rect 210002 513922 210058 513978
rect 240598 514294 240654 514350
rect 240722 514294 240778 514350
rect 240598 514170 240654 514226
rect 240722 514170 240778 514226
rect 240598 514046 240654 514102
rect 240722 514046 240778 514102
rect 240598 513922 240654 513978
rect 240722 513922 240778 513978
rect 271318 514294 271374 514350
rect 271442 514294 271498 514350
rect 271318 514170 271374 514226
rect 271442 514170 271498 514226
rect 271318 514046 271374 514102
rect 271442 514046 271498 514102
rect 271318 513922 271374 513978
rect 271442 513922 271498 513978
rect 302038 514294 302094 514350
rect 302162 514294 302218 514350
rect 302038 514170 302094 514226
rect 302162 514170 302218 514226
rect 302038 514046 302094 514102
rect 302162 514046 302218 514102
rect 302038 513922 302094 513978
rect 302162 513922 302218 513978
rect 332758 514294 332814 514350
rect 332882 514294 332938 514350
rect 332758 514170 332814 514226
rect 332882 514170 332938 514226
rect 332758 514046 332814 514102
rect 332882 514046 332938 514102
rect 332758 513922 332814 513978
rect 332882 513922 332938 513978
rect 363478 514294 363534 514350
rect 363602 514294 363658 514350
rect 363478 514170 363534 514226
rect 363602 514170 363658 514226
rect 363478 514046 363534 514102
rect 363602 514046 363658 514102
rect 363478 513922 363534 513978
rect 363602 513922 363658 513978
rect 394198 514294 394254 514350
rect 394322 514294 394378 514350
rect 394198 514170 394254 514226
rect 394322 514170 394378 514226
rect 394198 514046 394254 514102
rect 394322 514046 394378 514102
rect 394198 513922 394254 513978
rect 394322 513922 394378 513978
rect 424918 514294 424974 514350
rect 425042 514294 425098 514350
rect 424918 514170 424974 514226
rect 425042 514170 425098 514226
rect 424918 514046 424974 514102
rect 425042 514046 425098 514102
rect 424918 513922 424974 513978
rect 425042 513922 425098 513978
rect 225238 508294 225294 508350
rect 225362 508294 225418 508350
rect 225238 508170 225294 508226
rect 225362 508170 225418 508226
rect 225238 508046 225294 508102
rect 225362 508046 225418 508102
rect 225238 507922 225294 507978
rect 225362 507922 225418 507978
rect 255958 508294 256014 508350
rect 256082 508294 256138 508350
rect 255958 508170 256014 508226
rect 256082 508170 256138 508226
rect 255958 508046 256014 508102
rect 256082 508046 256138 508102
rect 255958 507922 256014 507978
rect 256082 507922 256138 507978
rect 286678 508294 286734 508350
rect 286802 508294 286858 508350
rect 286678 508170 286734 508226
rect 286802 508170 286858 508226
rect 286678 508046 286734 508102
rect 286802 508046 286858 508102
rect 286678 507922 286734 507978
rect 286802 507922 286858 507978
rect 317398 508294 317454 508350
rect 317522 508294 317578 508350
rect 317398 508170 317454 508226
rect 317522 508170 317578 508226
rect 317398 508046 317454 508102
rect 317522 508046 317578 508102
rect 317398 507922 317454 507978
rect 317522 507922 317578 507978
rect 348118 508294 348174 508350
rect 348242 508294 348298 508350
rect 348118 508170 348174 508226
rect 348242 508170 348298 508226
rect 348118 508046 348174 508102
rect 348242 508046 348298 508102
rect 348118 507922 348174 507978
rect 348242 507922 348298 507978
rect 378838 508294 378894 508350
rect 378962 508294 379018 508350
rect 378838 508170 378894 508226
rect 378962 508170 379018 508226
rect 378838 508046 378894 508102
rect 378962 508046 379018 508102
rect 378838 507922 378894 507978
rect 378962 507922 379018 507978
rect 409558 508294 409614 508350
rect 409682 508294 409738 508350
rect 409558 508170 409614 508226
rect 409682 508170 409738 508226
rect 409558 508046 409614 508102
rect 409682 508046 409738 508102
rect 409558 507922 409614 507978
rect 409682 507922 409738 507978
rect 440278 508294 440334 508350
rect 440402 508294 440458 508350
rect 440278 508170 440334 508226
rect 440402 508170 440458 508226
rect 440278 508046 440334 508102
rect 440402 508046 440458 508102
rect 440278 507922 440334 507978
rect 440402 507922 440458 507978
rect 209878 496294 209934 496350
rect 210002 496294 210058 496350
rect 209878 496170 209934 496226
rect 210002 496170 210058 496226
rect 209878 496046 209934 496102
rect 210002 496046 210058 496102
rect 209878 495922 209934 495978
rect 210002 495922 210058 495978
rect 240598 496294 240654 496350
rect 240722 496294 240778 496350
rect 240598 496170 240654 496226
rect 240722 496170 240778 496226
rect 240598 496046 240654 496102
rect 240722 496046 240778 496102
rect 240598 495922 240654 495978
rect 240722 495922 240778 495978
rect 271318 496294 271374 496350
rect 271442 496294 271498 496350
rect 271318 496170 271374 496226
rect 271442 496170 271498 496226
rect 271318 496046 271374 496102
rect 271442 496046 271498 496102
rect 271318 495922 271374 495978
rect 271442 495922 271498 495978
rect 302038 496294 302094 496350
rect 302162 496294 302218 496350
rect 302038 496170 302094 496226
rect 302162 496170 302218 496226
rect 302038 496046 302094 496102
rect 302162 496046 302218 496102
rect 302038 495922 302094 495978
rect 302162 495922 302218 495978
rect 332758 496294 332814 496350
rect 332882 496294 332938 496350
rect 332758 496170 332814 496226
rect 332882 496170 332938 496226
rect 332758 496046 332814 496102
rect 332882 496046 332938 496102
rect 332758 495922 332814 495978
rect 332882 495922 332938 495978
rect 363478 496294 363534 496350
rect 363602 496294 363658 496350
rect 363478 496170 363534 496226
rect 363602 496170 363658 496226
rect 363478 496046 363534 496102
rect 363602 496046 363658 496102
rect 363478 495922 363534 495978
rect 363602 495922 363658 495978
rect 394198 496294 394254 496350
rect 394322 496294 394378 496350
rect 394198 496170 394254 496226
rect 394322 496170 394378 496226
rect 394198 496046 394254 496102
rect 394322 496046 394378 496102
rect 394198 495922 394254 495978
rect 394322 495922 394378 495978
rect 424918 496294 424974 496350
rect 425042 496294 425098 496350
rect 424918 496170 424974 496226
rect 425042 496170 425098 496226
rect 424918 496046 424974 496102
rect 425042 496046 425098 496102
rect 424918 495922 424974 495978
rect 425042 495922 425098 495978
rect 225238 490294 225294 490350
rect 225362 490294 225418 490350
rect 225238 490170 225294 490226
rect 225362 490170 225418 490226
rect 225238 490046 225294 490102
rect 225362 490046 225418 490102
rect 225238 489922 225294 489978
rect 225362 489922 225418 489978
rect 255958 490294 256014 490350
rect 256082 490294 256138 490350
rect 255958 490170 256014 490226
rect 256082 490170 256138 490226
rect 255958 490046 256014 490102
rect 256082 490046 256138 490102
rect 255958 489922 256014 489978
rect 256082 489922 256138 489978
rect 286678 490294 286734 490350
rect 286802 490294 286858 490350
rect 286678 490170 286734 490226
rect 286802 490170 286858 490226
rect 286678 490046 286734 490102
rect 286802 490046 286858 490102
rect 286678 489922 286734 489978
rect 286802 489922 286858 489978
rect 317398 490294 317454 490350
rect 317522 490294 317578 490350
rect 317398 490170 317454 490226
rect 317522 490170 317578 490226
rect 317398 490046 317454 490102
rect 317522 490046 317578 490102
rect 317398 489922 317454 489978
rect 317522 489922 317578 489978
rect 348118 490294 348174 490350
rect 348242 490294 348298 490350
rect 348118 490170 348174 490226
rect 348242 490170 348298 490226
rect 348118 490046 348174 490102
rect 348242 490046 348298 490102
rect 348118 489922 348174 489978
rect 348242 489922 348298 489978
rect 378838 490294 378894 490350
rect 378962 490294 379018 490350
rect 378838 490170 378894 490226
rect 378962 490170 379018 490226
rect 378838 490046 378894 490102
rect 378962 490046 379018 490102
rect 378838 489922 378894 489978
rect 378962 489922 379018 489978
rect 409558 490294 409614 490350
rect 409682 490294 409738 490350
rect 409558 490170 409614 490226
rect 409682 490170 409738 490226
rect 409558 490046 409614 490102
rect 409682 490046 409738 490102
rect 409558 489922 409614 489978
rect 409682 489922 409738 489978
rect 440278 490294 440334 490350
rect 440402 490294 440458 490350
rect 440278 490170 440334 490226
rect 440402 490170 440458 490226
rect 440278 490046 440334 490102
rect 440402 490046 440458 490102
rect 440278 489922 440334 489978
rect 440402 489922 440458 489978
rect 209878 478294 209934 478350
rect 210002 478294 210058 478350
rect 209878 478170 209934 478226
rect 210002 478170 210058 478226
rect 209878 478046 209934 478102
rect 210002 478046 210058 478102
rect 209878 477922 209934 477978
rect 210002 477922 210058 477978
rect 240598 478294 240654 478350
rect 240722 478294 240778 478350
rect 240598 478170 240654 478226
rect 240722 478170 240778 478226
rect 240598 478046 240654 478102
rect 240722 478046 240778 478102
rect 240598 477922 240654 477978
rect 240722 477922 240778 477978
rect 271318 478294 271374 478350
rect 271442 478294 271498 478350
rect 271318 478170 271374 478226
rect 271442 478170 271498 478226
rect 271318 478046 271374 478102
rect 271442 478046 271498 478102
rect 271318 477922 271374 477978
rect 271442 477922 271498 477978
rect 302038 478294 302094 478350
rect 302162 478294 302218 478350
rect 302038 478170 302094 478226
rect 302162 478170 302218 478226
rect 302038 478046 302094 478102
rect 302162 478046 302218 478102
rect 302038 477922 302094 477978
rect 302162 477922 302218 477978
rect 332758 478294 332814 478350
rect 332882 478294 332938 478350
rect 332758 478170 332814 478226
rect 332882 478170 332938 478226
rect 332758 478046 332814 478102
rect 332882 478046 332938 478102
rect 332758 477922 332814 477978
rect 332882 477922 332938 477978
rect 363478 478294 363534 478350
rect 363602 478294 363658 478350
rect 363478 478170 363534 478226
rect 363602 478170 363658 478226
rect 363478 478046 363534 478102
rect 363602 478046 363658 478102
rect 363478 477922 363534 477978
rect 363602 477922 363658 477978
rect 394198 478294 394254 478350
rect 394322 478294 394378 478350
rect 394198 478170 394254 478226
rect 394322 478170 394378 478226
rect 394198 478046 394254 478102
rect 394322 478046 394378 478102
rect 394198 477922 394254 477978
rect 394322 477922 394378 477978
rect 424918 478294 424974 478350
rect 425042 478294 425098 478350
rect 424918 478170 424974 478226
rect 425042 478170 425098 478226
rect 424918 478046 424974 478102
rect 425042 478046 425098 478102
rect 424918 477922 424974 477978
rect 425042 477922 425098 477978
rect 225238 472294 225294 472350
rect 225362 472294 225418 472350
rect 225238 472170 225294 472226
rect 225362 472170 225418 472226
rect 225238 472046 225294 472102
rect 225362 472046 225418 472102
rect 225238 471922 225294 471978
rect 225362 471922 225418 471978
rect 255958 472294 256014 472350
rect 256082 472294 256138 472350
rect 255958 472170 256014 472226
rect 256082 472170 256138 472226
rect 255958 472046 256014 472102
rect 256082 472046 256138 472102
rect 255958 471922 256014 471978
rect 256082 471922 256138 471978
rect 286678 472294 286734 472350
rect 286802 472294 286858 472350
rect 286678 472170 286734 472226
rect 286802 472170 286858 472226
rect 286678 472046 286734 472102
rect 286802 472046 286858 472102
rect 286678 471922 286734 471978
rect 286802 471922 286858 471978
rect 317398 472294 317454 472350
rect 317522 472294 317578 472350
rect 317398 472170 317454 472226
rect 317522 472170 317578 472226
rect 317398 472046 317454 472102
rect 317522 472046 317578 472102
rect 317398 471922 317454 471978
rect 317522 471922 317578 471978
rect 348118 472294 348174 472350
rect 348242 472294 348298 472350
rect 348118 472170 348174 472226
rect 348242 472170 348298 472226
rect 348118 472046 348174 472102
rect 348242 472046 348298 472102
rect 348118 471922 348174 471978
rect 348242 471922 348298 471978
rect 378838 472294 378894 472350
rect 378962 472294 379018 472350
rect 378838 472170 378894 472226
rect 378962 472170 379018 472226
rect 378838 472046 378894 472102
rect 378962 472046 379018 472102
rect 378838 471922 378894 471978
rect 378962 471922 379018 471978
rect 409558 472294 409614 472350
rect 409682 472294 409738 472350
rect 409558 472170 409614 472226
rect 409682 472170 409738 472226
rect 409558 472046 409614 472102
rect 409682 472046 409738 472102
rect 409558 471922 409614 471978
rect 409682 471922 409738 471978
rect 440278 472294 440334 472350
rect 440402 472294 440458 472350
rect 440278 472170 440334 472226
rect 440402 472170 440458 472226
rect 440278 472046 440334 472102
rect 440402 472046 440458 472102
rect 440278 471922 440334 471978
rect 440402 471922 440458 471978
rect 209878 460294 209934 460350
rect 210002 460294 210058 460350
rect 209878 460170 209934 460226
rect 210002 460170 210058 460226
rect 209878 460046 209934 460102
rect 210002 460046 210058 460102
rect 209878 459922 209934 459978
rect 210002 459922 210058 459978
rect 240598 460294 240654 460350
rect 240722 460294 240778 460350
rect 240598 460170 240654 460226
rect 240722 460170 240778 460226
rect 240598 460046 240654 460102
rect 240722 460046 240778 460102
rect 240598 459922 240654 459978
rect 240722 459922 240778 459978
rect 271318 460294 271374 460350
rect 271442 460294 271498 460350
rect 271318 460170 271374 460226
rect 271442 460170 271498 460226
rect 271318 460046 271374 460102
rect 271442 460046 271498 460102
rect 271318 459922 271374 459978
rect 271442 459922 271498 459978
rect 302038 460294 302094 460350
rect 302162 460294 302218 460350
rect 302038 460170 302094 460226
rect 302162 460170 302218 460226
rect 302038 460046 302094 460102
rect 302162 460046 302218 460102
rect 302038 459922 302094 459978
rect 302162 459922 302218 459978
rect 332758 460294 332814 460350
rect 332882 460294 332938 460350
rect 332758 460170 332814 460226
rect 332882 460170 332938 460226
rect 332758 460046 332814 460102
rect 332882 460046 332938 460102
rect 332758 459922 332814 459978
rect 332882 459922 332938 459978
rect 363478 460294 363534 460350
rect 363602 460294 363658 460350
rect 363478 460170 363534 460226
rect 363602 460170 363658 460226
rect 363478 460046 363534 460102
rect 363602 460046 363658 460102
rect 363478 459922 363534 459978
rect 363602 459922 363658 459978
rect 394198 460294 394254 460350
rect 394322 460294 394378 460350
rect 394198 460170 394254 460226
rect 394322 460170 394378 460226
rect 394198 460046 394254 460102
rect 394322 460046 394378 460102
rect 394198 459922 394254 459978
rect 394322 459922 394378 459978
rect 424918 460294 424974 460350
rect 425042 460294 425098 460350
rect 424918 460170 424974 460226
rect 425042 460170 425098 460226
rect 424918 460046 424974 460102
rect 425042 460046 425098 460102
rect 424918 459922 424974 459978
rect 425042 459922 425098 459978
rect 225238 454294 225294 454350
rect 225362 454294 225418 454350
rect 225238 454170 225294 454226
rect 225362 454170 225418 454226
rect 225238 454046 225294 454102
rect 225362 454046 225418 454102
rect 225238 453922 225294 453978
rect 225362 453922 225418 453978
rect 255958 454294 256014 454350
rect 256082 454294 256138 454350
rect 255958 454170 256014 454226
rect 256082 454170 256138 454226
rect 255958 454046 256014 454102
rect 256082 454046 256138 454102
rect 255958 453922 256014 453978
rect 256082 453922 256138 453978
rect 286678 454294 286734 454350
rect 286802 454294 286858 454350
rect 286678 454170 286734 454226
rect 286802 454170 286858 454226
rect 286678 454046 286734 454102
rect 286802 454046 286858 454102
rect 286678 453922 286734 453978
rect 286802 453922 286858 453978
rect 317398 454294 317454 454350
rect 317522 454294 317578 454350
rect 317398 454170 317454 454226
rect 317522 454170 317578 454226
rect 317398 454046 317454 454102
rect 317522 454046 317578 454102
rect 317398 453922 317454 453978
rect 317522 453922 317578 453978
rect 348118 454294 348174 454350
rect 348242 454294 348298 454350
rect 348118 454170 348174 454226
rect 348242 454170 348298 454226
rect 348118 454046 348174 454102
rect 348242 454046 348298 454102
rect 348118 453922 348174 453978
rect 348242 453922 348298 453978
rect 378838 454294 378894 454350
rect 378962 454294 379018 454350
rect 378838 454170 378894 454226
rect 378962 454170 379018 454226
rect 378838 454046 378894 454102
rect 378962 454046 379018 454102
rect 378838 453922 378894 453978
rect 378962 453922 379018 453978
rect 409558 454294 409614 454350
rect 409682 454294 409738 454350
rect 409558 454170 409614 454226
rect 409682 454170 409738 454226
rect 409558 454046 409614 454102
rect 409682 454046 409738 454102
rect 409558 453922 409614 453978
rect 409682 453922 409738 453978
rect 440278 454294 440334 454350
rect 440402 454294 440458 454350
rect 440278 454170 440334 454226
rect 440402 454170 440458 454226
rect 440278 454046 440334 454102
rect 440402 454046 440458 454102
rect 440278 453922 440334 453978
rect 440402 453922 440458 453978
rect 209878 442294 209934 442350
rect 210002 442294 210058 442350
rect 209878 442170 209934 442226
rect 210002 442170 210058 442226
rect 209878 442046 209934 442102
rect 210002 442046 210058 442102
rect 209878 441922 209934 441978
rect 210002 441922 210058 441978
rect 240598 442294 240654 442350
rect 240722 442294 240778 442350
rect 240598 442170 240654 442226
rect 240722 442170 240778 442226
rect 240598 442046 240654 442102
rect 240722 442046 240778 442102
rect 240598 441922 240654 441978
rect 240722 441922 240778 441978
rect 271318 442294 271374 442350
rect 271442 442294 271498 442350
rect 271318 442170 271374 442226
rect 271442 442170 271498 442226
rect 271318 442046 271374 442102
rect 271442 442046 271498 442102
rect 271318 441922 271374 441978
rect 271442 441922 271498 441978
rect 302038 442294 302094 442350
rect 302162 442294 302218 442350
rect 302038 442170 302094 442226
rect 302162 442170 302218 442226
rect 302038 442046 302094 442102
rect 302162 442046 302218 442102
rect 302038 441922 302094 441978
rect 302162 441922 302218 441978
rect 332758 442294 332814 442350
rect 332882 442294 332938 442350
rect 332758 442170 332814 442226
rect 332882 442170 332938 442226
rect 332758 442046 332814 442102
rect 332882 442046 332938 442102
rect 332758 441922 332814 441978
rect 332882 441922 332938 441978
rect 363478 442294 363534 442350
rect 363602 442294 363658 442350
rect 363478 442170 363534 442226
rect 363602 442170 363658 442226
rect 363478 442046 363534 442102
rect 363602 442046 363658 442102
rect 363478 441922 363534 441978
rect 363602 441922 363658 441978
rect 394198 442294 394254 442350
rect 394322 442294 394378 442350
rect 394198 442170 394254 442226
rect 394322 442170 394378 442226
rect 394198 442046 394254 442102
rect 394322 442046 394378 442102
rect 394198 441922 394254 441978
rect 394322 441922 394378 441978
rect 424918 442294 424974 442350
rect 425042 442294 425098 442350
rect 424918 442170 424974 442226
rect 425042 442170 425098 442226
rect 424918 442046 424974 442102
rect 425042 442046 425098 442102
rect 424918 441922 424974 441978
rect 425042 441922 425098 441978
rect 225238 436294 225294 436350
rect 225362 436294 225418 436350
rect 225238 436170 225294 436226
rect 225362 436170 225418 436226
rect 225238 436046 225294 436102
rect 225362 436046 225418 436102
rect 225238 435922 225294 435978
rect 225362 435922 225418 435978
rect 255958 436294 256014 436350
rect 256082 436294 256138 436350
rect 255958 436170 256014 436226
rect 256082 436170 256138 436226
rect 255958 436046 256014 436102
rect 256082 436046 256138 436102
rect 255958 435922 256014 435978
rect 256082 435922 256138 435978
rect 286678 436294 286734 436350
rect 286802 436294 286858 436350
rect 286678 436170 286734 436226
rect 286802 436170 286858 436226
rect 286678 436046 286734 436102
rect 286802 436046 286858 436102
rect 286678 435922 286734 435978
rect 286802 435922 286858 435978
rect 317398 436294 317454 436350
rect 317522 436294 317578 436350
rect 317398 436170 317454 436226
rect 317522 436170 317578 436226
rect 317398 436046 317454 436102
rect 317522 436046 317578 436102
rect 317398 435922 317454 435978
rect 317522 435922 317578 435978
rect 348118 436294 348174 436350
rect 348242 436294 348298 436350
rect 348118 436170 348174 436226
rect 348242 436170 348298 436226
rect 348118 436046 348174 436102
rect 348242 436046 348298 436102
rect 348118 435922 348174 435978
rect 348242 435922 348298 435978
rect 378838 436294 378894 436350
rect 378962 436294 379018 436350
rect 378838 436170 378894 436226
rect 378962 436170 379018 436226
rect 378838 436046 378894 436102
rect 378962 436046 379018 436102
rect 378838 435922 378894 435978
rect 378962 435922 379018 435978
rect 409558 436294 409614 436350
rect 409682 436294 409738 436350
rect 409558 436170 409614 436226
rect 409682 436170 409738 436226
rect 409558 436046 409614 436102
rect 409682 436046 409738 436102
rect 409558 435922 409614 435978
rect 409682 435922 409738 435978
rect 440278 436294 440334 436350
rect 440402 436294 440458 436350
rect 440278 436170 440334 436226
rect 440402 436170 440458 436226
rect 440278 436046 440334 436102
rect 440402 436046 440458 436102
rect 440278 435922 440334 435978
rect 440402 435922 440458 435978
rect 209878 424294 209934 424350
rect 210002 424294 210058 424350
rect 209878 424170 209934 424226
rect 210002 424170 210058 424226
rect 209878 424046 209934 424102
rect 210002 424046 210058 424102
rect 209878 423922 209934 423978
rect 210002 423922 210058 423978
rect 240598 424294 240654 424350
rect 240722 424294 240778 424350
rect 240598 424170 240654 424226
rect 240722 424170 240778 424226
rect 240598 424046 240654 424102
rect 240722 424046 240778 424102
rect 240598 423922 240654 423978
rect 240722 423922 240778 423978
rect 271318 424294 271374 424350
rect 271442 424294 271498 424350
rect 271318 424170 271374 424226
rect 271442 424170 271498 424226
rect 271318 424046 271374 424102
rect 271442 424046 271498 424102
rect 271318 423922 271374 423978
rect 271442 423922 271498 423978
rect 302038 424294 302094 424350
rect 302162 424294 302218 424350
rect 302038 424170 302094 424226
rect 302162 424170 302218 424226
rect 302038 424046 302094 424102
rect 302162 424046 302218 424102
rect 302038 423922 302094 423978
rect 302162 423922 302218 423978
rect 332758 424294 332814 424350
rect 332882 424294 332938 424350
rect 332758 424170 332814 424226
rect 332882 424170 332938 424226
rect 332758 424046 332814 424102
rect 332882 424046 332938 424102
rect 332758 423922 332814 423978
rect 332882 423922 332938 423978
rect 363478 424294 363534 424350
rect 363602 424294 363658 424350
rect 363478 424170 363534 424226
rect 363602 424170 363658 424226
rect 363478 424046 363534 424102
rect 363602 424046 363658 424102
rect 363478 423922 363534 423978
rect 363602 423922 363658 423978
rect 394198 424294 394254 424350
rect 394322 424294 394378 424350
rect 394198 424170 394254 424226
rect 394322 424170 394378 424226
rect 394198 424046 394254 424102
rect 394322 424046 394378 424102
rect 394198 423922 394254 423978
rect 394322 423922 394378 423978
rect 424918 424294 424974 424350
rect 425042 424294 425098 424350
rect 424918 424170 424974 424226
rect 425042 424170 425098 424226
rect 424918 424046 424974 424102
rect 425042 424046 425098 424102
rect 424918 423922 424974 423978
rect 425042 423922 425098 423978
rect 225238 418294 225294 418350
rect 225362 418294 225418 418350
rect 225238 418170 225294 418226
rect 225362 418170 225418 418226
rect 225238 418046 225294 418102
rect 225362 418046 225418 418102
rect 225238 417922 225294 417978
rect 225362 417922 225418 417978
rect 255958 418294 256014 418350
rect 256082 418294 256138 418350
rect 255958 418170 256014 418226
rect 256082 418170 256138 418226
rect 255958 418046 256014 418102
rect 256082 418046 256138 418102
rect 255958 417922 256014 417978
rect 256082 417922 256138 417978
rect 286678 418294 286734 418350
rect 286802 418294 286858 418350
rect 286678 418170 286734 418226
rect 286802 418170 286858 418226
rect 286678 418046 286734 418102
rect 286802 418046 286858 418102
rect 286678 417922 286734 417978
rect 286802 417922 286858 417978
rect 317398 418294 317454 418350
rect 317522 418294 317578 418350
rect 317398 418170 317454 418226
rect 317522 418170 317578 418226
rect 317398 418046 317454 418102
rect 317522 418046 317578 418102
rect 317398 417922 317454 417978
rect 317522 417922 317578 417978
rect 348118 418294 348174 418350
rect 348242 418294 348298 418350
rect 348118 418170 348174 418226
rect 348242 418170 348298 418226
rect 348118 418046 348174 418102
rect 348242 418046 348298 418102
rect 348118 417922 348174 417978
rect 348242 417922 348298 417978
rect 378838 418294 378894 418350
rect 378962 418294 379018 418350
rect 378838 418170 378894 418226
rect 378962 418170 379018 418226
rect 378838 418046 378894 418102
rect 378962 418046 379018 418102
rect 378838 417922 378894 417978
rect 378962 417922 379018 417978
rect 409558 418294 409614 418350
rect 409682 418294 409738 418350
rect 409558 418170 409614 418226
rect 409682 418170 409738 418226
rect 409558 418046 409614 418102
rect 409682 418046 409738 418102
rect 409558 417922 409614 417978
rect 409682 417922 409738 417978
rect 440278 418294 440334 418350
rect 440402 418294 440458 418350
rect 440278 418170 440334 418226
rect 440402 418170 440458 418226
rect 440278 418046 440334 418102
rect 440402 418046 440458 418102
rect 440278 417922 440334 417978
rect 440402 417922 440458 417978
rect 354396 409742 354452 409798
rect 289772 409382 289828 409438
rect 288876 409202 288932 409258
rect 209916 404342 209972 404398
rect 209804 402722 209860 402778
rect 220554 400294 220610 400350
rect 220678 400294 220734 400350
rect 220802 400294 220858 400350
rect 220926 400294 220982 400350
rect 220554 400170 220610 400226
rect 220678 400170 220734 400226
rect 220802 400170 220858 400226
rect 220926 400170 220982 400226
rect 220554 400046 220610 400102
rect 220678 400046 220734 400102
rect 220802 400046 220858 400102
rect 220926 400046 220982 400102
rect 220554 399922 220610 399978
rect 220678 399922 220734 399978
rect 220802 399922 220858 399978
rect 220926 399922 220982 399978
rect 220554 382294 220610 382350
rect 220678 382294 220734 382350
rect 220802 382294 220858 382350
rect 220926 382294 220982 382350
rect 220554 382170 220610 382226
rect 220678 382170 220734 382226
rect 220802 382170 220858 382226
rect 220926 382170 220982 382226
rect 220554 382046 220610 382102
rect 220678 382046 220734 382102
rect 220802 382046 220858 382102
rect 220926 382046 220982 382102
rect 220554 381922 220610 381978
rect 220678 381922 220734 381978
rect 220802 381922 220858 381978
rect 220926 381922 220982 381978
rect 209878 370294 209934 370350
rect 210002 370294 210058 370350
rect 209878 370170 209934 370226
rect 210002 370170 210058 370226
rect 209878 370046 209934 370102
rect 210002 370046 210058 370102
rect 209878 369922 209934 369978
rect 210002 369922 210058 369978
rect 210812 367982 210868 368038
rect 209878 352294 209934 352350
rect 210002 352294 210058 352350
rect 209878 352170 209934 352226
rect 210002 352170 210058 352226
rect 209878 352046 209934 352102
rect 210002 352046 210058 352102
rect 209878 351922 209934 351978
rect 210002 351922 210058 351978
rect 206668 340082 206724 340138
rect 209878 334294 209934 334350
rect 210002 334294 210058 334350
rect 209878 334170 209934 334226
rect 210002 334170 210058 334226
rect 209878 334046 209934 334102
rect 210002 334046 210058 334102
rect 209878 333922 209934 333978
rect 210002 333922 210058 333978
rect 209878 316294 209934 316350
rect 210002 316294 210058 316350
rect 209878 316170 209934 316226
rect 210002 316170 210058 316226
rect 209878 316046 209934 316102
rect 210002 316046 210058 316102
rect 209878 315922 209934 315978
rect 210002 315922 210058 315978
rect 209878 298294 209934 298350
rect 210002 298294 210058 298350
rect 209878 298170 209934 298226
rect 210002 298170 210058 298226
rect 209878 298046 209934 298102
rect 210002 298046 210058 298102
rect 209878 297922 209934 297978
rect 210002 297922 210058 297978
rect 209878 280294 209934 280350
rect 210002 280294 210058 280350
rect 209878 280170 209934 280226
rect 210002 280170 210058 280226
rect 209878 280046 209934 280102
rect 210002 280046 210058 280102
rect 209878 279922 209934 279978
rect 210002 279922 210058 279978
rect 209878 262294 209934 262350
rect 210002 262294 210058 262350
rect 209878 262170 209934 262226
rect 210002 262170 210058 262226
rect 209878 262046 209934 262102
rect 210002 262046 210058 262102
rect 209878 261922 209934 261978
rect 210002 261922 210058 261978
rect 209878 244294 209934 244350
rect 210002 244294 210058 244350
rect 209878 244170 209934 244226
rect 210002 244170 210058 244226
rect 209878 244046 209934 244102
rect 210002 244046 210058 244102
rect 209878 243922 209934 243978
rect 210002 243922 210058 243978
rect 209916 231002 209972 231058
rect 214172 366542 214228 366598
rect 217532 366362 217588 366418
rect 214284 364562 214340 364618
rect 224274 406294 224330 406350
rect 224398 406294 224454 406350
rect 224522 406294 224578 406350
rect 224646 406294 224702 406350
rect 224274 406170 224330 406226
rect 224398 406170 224454 406226
rect 224522 406170 224578 406226
rect 224646 406170 224702 406226
rect 224274 406046 224330 406102
rect 224398 406046 224454 406102
rect 224522 406046 224578 406102
rect 224646 406046 224702 406102
rect 224274 405922 224330 405978
rect 224398 405922 224454 405978
rect 224522 405922 224578 405978
rect 224646 405922 224702 405978
rect 224274 388294 224330 388350
rect 224398 388294 224454 388350
rect 224522 388294 224578 388350
rect 224646 388294 224702 388350
rect 224274 388170 224330 388226
rect 224398 388170 224454 388226
rect 224522 388170 224578 388226
rect 224646 388170 224702 388226
rect 224274 388046 224330 388102
rect 224398 388046 224454 388102
rect 224522 388046 224578 388102
rect 224646 388046 224702 388102
rect 224274 387922 224330 387978
rect 224398 387922 224454 387978
rect 224522 387922 224578 387978
rect 224646 387922 224702 387978
rect 224028 378782 224084 378838
rect 222012 372122 222068 372178
rect 220554 364294 220610 364350
rect 220678 364294 220734 364350
rect 220802 364294 220858 364350
rect 220926 364294 220982 364350
rect 220554 364170 220610 364226
rect 220678 364170 220734 364226
rect 220802 364170 220858 364226
rect 220926 364170 220982 364226
rect 220554 364046 220610 364102
rect 220678 364046 220734 364102
rect 220802 364046 220858 364102
rect 220926 364046 220982 364102
rect 220554 363922 220610 363978
rect 220678 363922 220734 363978
rect 220802 363922 220858 363978
rect 220926 363922 220982 363978
rect 220554 346294 220610 346350
rect 220678 346294 220734 346350
rect 220802 346294 220858 346350
rect 220926 346294 220982 346350
rect 220554 346170 220610 346226
rect 220678 346170 220734 346226
rect 220802 346170 220858 346226
rect 220926 346170 220982 346226
rect 220554 346046 220610 346102
rect 220678 346046 220734 346102
rect 220802 346046 220858 346102
rect 220926 346046 220982 346102
rect 220554 345922 220610 345978
rect 220678 345922 220734 345978
rect 220802 345922 220858 345978
rect 220926 345922 220982 345978
rect 220554 328294 220610 328350
rect 220678 328294 220734 328350
rect 220802 328294 220858 328350
rect 220926 328294 220982 328350
rect 220554 328170 220610 328226
rect 220678 328170 220734 328226
rect 220802 328170 220858 328226
rect 220926 328170 220982 328226
rect 220554 328046 220610 328102
rect 220678 328046 220734 328102
rect 220802 328046 220858 328102
rect 220926 328046 220982 328102
rect 220554 327922 220610 327978
rect 220678 327922 220734 327978
rect 220802 327922 220858 327978
rect 220926 327922 220982 327978
rect 217644 319202 217700 319258
rect 220554 310294 220610 310350
rect 220678 310294 220734 310350
rect 220802 310294 220858 310350
rect 220926 310294 220982 310350
rect 220554 310170 220610 310226
rect 220678 310170 220734 310226
rect 220802 310170 220858 310226
rect 220926 310170 220982 310226
rect 220554 310046 220610 310102
rect 220678 310046 220734 310102
rect 220802 310046 220858 310102
rect 220926 310046 220982 310102
rect 220554 309922 220610 309978
rect 220678 309922 220734 309978
rect 220802 309922 220858 309978
rect 220926 309922 220982 309978
rect 220554 292294 220610 292350
rect 220678 292294 220734 292350
rect 220802 292294 220858 292350
rect 220926 292294 220982 292350
rect 220554 292170 220610 292226
rect 220678 292170 220734 292226
rect 220802 292170 220858 292226
rect 220926 292170 220982 292226
rect 220554 292046 220610 292102
rect 220678 292046 220734 292102
rect 220802 292046 220858 292102
rect 220926 292046 220982 292102
rect 220554 291922 220610 291978
rect 220678 291922 220734 291978
rect 220802 291922 220858 291978
rect 220926 291922 220982 291978
rect 220554 274294 220610 274350
rect 220678 274294 220734 274350
rect 220802 274294 220858 274350
rect 220926 274294 220982 274350
rect 220554 274170 220610 274226
rect 220678 274170 220734 274226
rect 220802 274170 220858 274226
rect 220926 274170 220982 274226
rect 220554 274046 220610 274102
rect 220678 274046 220734 274102
rect 220802 274046 220858 274102
rect 220926 274046 220982 274102
rect 220554 273922 220610 273978
rect 220678 273922 220734 273978
rect 220802 273922 220858 273978
rect 220926 273922 220982 273978
rect 220554 256294 220610 256350
rect 220678 256294 220734 256350
rect 220802 256294 220858 256350
rect 220926 256294 220982 256350
rect 220554 256170 220610 256226
rect 220678 256170 220734 256226
rect 220802 256170 220858 256226
rect 220926 256170 220982 256226
rect 220554 256046 220610 256102
rect 220678 256046 220734 256102
rect 220802 256046 220858 256102
rect 220926 256046 220982 256102
rect 220554 255922 220610 255978
rect 220678 255922 220734 255978
rect 220802 255922 220858 255978
rect 220926 255922 220982 255978
rect 220554 238294 220610 238350
rect 220678 238294 220734 238350
rect 220802 238294 220858 238350
rect 220926 238294 220982 238350
rect 220554 238170 220610 238226
rect 220678 238170 220734 238226
rect 220802 238170 220858 238226
rect 220926 238170 220982 238226
rect 220554 238046 220610 238102
rect 220678 238046 220734 238102
rect 220802 238046 220858 238102
rect 220926 238046 220982 238102
rect 220554 237922 220610 237978
rect 220678 237922 220734 237978
rect 220802 237922 220858 237978
rect 220926 237922 220982 237978
rect 220554 220294 220610 220350
rect 220678 220294 220734 220350
rect 220802 220294 220858 220350
rect 220926 220294 220982 220350
rect 220554 220170 220610 220226
rect 220678 220170 220734 220226
rect 220802 220170 220858 220226
rect 220926 220170 220982 220226
rect 220554 220046 220610 220102
rect 220678 220046 220734 220102
rect 220802 220046 220858 220102
rect 220926 220046 220982 220102
rect 220554 219922 220610 219978
rect 220678 219922 220734 219978
rect 220802 219922 220858 219978
rect 220926 219922 220982 219978
rect 226716 394802 226772 394858
rect 225148 377342 225204 377398
rect 225820 377162 225876 377218
rect 224274 370294 224330 370350
rect 224398 370294 224454 370350
rect 224522 370294 224578 370350
rect 224646 370294 224702 370350
rect 224274 370170 224330 370226
rect 224398 370170 224454 370226
rect 224522 370170 224578 370226
rect 224646 370170 224702 370226
rect 224274 370046 224330 370102
rect 224398 370046 224454 370102
rect 224522 370046 224578 370102
rect 224646 370046 224702 370102
rect 224274 369922 224330 369978
rect 224398 369922 224454 369978
rect 224522 369922 224578 369978
rect 224646 369922 224702 369978
rect 225238 364294 225294 364350
rect 225362 364294 225418 364350
rect 225238 364170 225294 364226
rect 225362 364170 225418 364226
rect 225238 364046 225294 364102
rect 225362 364046 225418 364102
rect 225238 363922 225294 363978
rect 225362 363922 225418 363978
rect 224274 352294 224330 352350
rect 224398 352294 224454 352350
rect 224522 352294 224578 352350
rect 224646 352294 224702 352350
rect 224274 352170 224330 352226
rect 224398 352170 224454 352226
rect 224522 352170 224578 352226
rect 224646 352170 224702 352226
rect 224274 352046 224330 352102
rect 224398 352046 224454 352102
rect 224522 352046 224578 352102
rect 224646 352046 224702 352102
rect 224274 351922 224330 351978
rect 224398 351922 224454 351978
rect 224522 351922 224578 351978
rect 224646 351922 224702 351978
rect 225238 346294 225294 346350
rect 225362 346294 225418 346350
rect 225238 346170 225294 346226
rect 225362 346170 225418 346226
rect 225238 346046 225294 346102
rect 225362 346046 225418 346102
rect 225238 345922 225294 345978
rect 225362 345922 225418 345978
rect 224274 334294 224330 334350
rect 224398 334294 224454 334350
rect 224522 334294 224578 334350
rect 224646 334294 224702 334350
rect 224274 334170 224330 334226
rect 224398 334170 224454 334226
rect 224522 334170 224578 334226
rect 224646 334170 224702 334226
rect 224274 334046 224330 334102
rect 224398 334046 224454 334102
rect 224522 334046 224578 334102
rect 224646 334046 224702 334102
rect 224274 333922 224330 333978
rect 224398 333922 224454 333978
rect 224522 333922 224578 333978
rect 224646 333922 224702 333978
rect 225238 328294 225294 328350
rect 225362 328294 225418 328350
rect 225238 328170 225294 328226
rect 225362 328170 225418 328226
rect 225238 328046 225294 328102
rect 225362 328046 225418 328102
rect 225238 327922 225294 327978
rect 225362 327922 225418 327978
rect 224274 316294 224330 316350
rect 224398 316294 224454 316350
rect 224522 316294 224578 316350
rect 224646 316294 224702 316350
rect 224274 316170 224330 316226
rect 224398 316170 224454 316226
rect 224522 316170 224578 316226
rect 224646 316170 224702 316226
rect 224274 316046 224330 316102
rect 224398 316046 224454 316102
rect 224522 316046 224578 316102
rect 224646 316046 224702 316102
rect 224274 315922 224330 315978
rect 224398 315922 224454 315978
rect 224522 315922 224578 315978
rect 224646 315922 224702 315978
rect 225238 310294 225294 310350
rect 225362 310294 225418 310350
rect 225238 310170 225294 310226
rect 225362 310170 225418 310226
rect 225238 310046 225294 310102
rect 225362 310046 225418 310102
rect 225238 309922 225294 309978
rect 225362 309922 225418 309978
rect 224274 298294 224330 298350
rect 224398 298294 224454 298350
rect 224522 298294 224578 298350
rect 224646 298294 224702 298350
rect 224274 298170 224330 298226
rect 224398 298170 224454 298226
rect 224522 298170 224578 298226
rect 224646 298170 224702 298226
rect 224274 298046 224330 298102
rect 224398 298046 224454 298102
rect 224522 298046 224578 298102
rect 224646 298046 224702 298102
rect 224274 297922 224330 297978
rect 224398 297922 224454 297978
rect 224522 297922 224578 297978
rect 224646 297922 224702 297978
rect 225238 292294 225294 292350
rect 225362 292294 225418 292350
rect 225238 292170 225294 292226
rect 225362 292170 225418 292226
rect 225238 292046 225294 292102
rect 225362 292046 225418 292102
rect 225238 291922 225294 291978
rect 225362 291922 225418 291978
rect 224274 280294 224330 280350
rect 224398 280294 224454 280350
rect 224522 280294 224578 280350
rect 224646 280294 224702 280350
rect 224274 280170 224330 280226
rect 224398 280170 224454 280226
rect 224522 280170 224578 280226
rect 224646 280170 224702 280226
rect 224274 280046 224330 280102
rect 224398 280046 224454 280102
rect 224522 280046 224578 280102
rect 224646 280046 224702 280102
rect 224274 279922 224330 279978
rect 224398 279922 224454 279978
rect 224522 279922 224578 279978
rect 224646 279922 224702 279978
rect 225238 274294 225294 274350
rect 225362 274294 225418 274350
rect 225238 274170 225294 274226
rect 225362 274170 225418 274226
rect 225238 274046 225294 274102
rect 225362 274046 225418 274102
rect 225238 273922 225294 273978
rect 225362 273922 225418 273978
rect 224274 262294 224330 262350
rect 224398 262294 224454 262350
rect 224522 262294 224578 262350
rect 224646 262294 224702 262350
rect 224274 262170 224330 262226
rect 224398 262170 224454 262226
rect 224522 262170 224578 262226
rect 224646 262170 224702 262226
rect 224274 262046 224330 262102
rect 224398 262046 224454 262102
rect 224522 262046 224578 262102
rect 224646 262046 224702 262102
rect 224274 261922 224330 261978
rect 224398 261922 224454 261978
rect 224522 261922 224578 261978
rect 224646 261922 224702 261978
rect 225238 256294 225294 256350
rect 225362 256294 225418 256350
rect 225238 256170 225294 256226
rect 225362 256170 225418 256226
rect 225238 256046 225294 256102
rect 225362 256046 225418 256102
rect 225238 255922 225294 255978
rect 225362 255922 225418 255978
rect 224274 244294 224330 244350
rect 224398 244294 224454 244350
rect 224522 244294 224578 244350
rect 224646 244294 224702 244350
rect 224274 244170 224330 244226
rect 224398 244170 224454 244226
rect 224522 244170 224578 244226
rect 224646 244170 224702 244226
rect 224274 244046 224330 244102
rect 224398 244046 224454 244102
rect 224522 244046 224578 244102
rect 224646 244046 224702 244102
rect 224274 243922 224330 243978
rect 224398 243922 224454 243978
rect 224522 243922 224578 243978
rect 224646 243922 224702 243978
rect 224274 226294 224330 226350
rect 224398 226294 224454 226350
rect 224522 226294 224578 226350
rect 224646 226294 224702 226350
rect 224274 226170 224330 226226
rect 224398 226170 224454 226226
rect 224522 226170 224578 226226
rect 224646 226170 224702 226226
rect 224274 226046 224330 226102
rect 224398 226046 224454 226102
rect 224522 226046 224578 226102
rect 224646 226046 224702 226102
rect 224274 225922 224330 225978
rect 224398 225922 224454 225978
rect 224522 225922 224578 225978
rect 224646 225922 224702 225978
rect 225148 224162 225204 224218
rect 251274 400294 251330 400350
rect 251398 400294 251454 400350
rect 251522 400294 251578 400350
rect 251646 400294 251702 400350
rect 251274 400170 251330 400226
rect 251398 400170 251454 400226
rect 251522 400170 251578 400226
rect 251646 400170 251702 400226
rect 251274 400046 251330 400102
rect 251398 400046 251454 400102
rect 251522 400046 251578 400102
rect 251646 400046 251702 400102
rect 251274 399922 251330 399978
rect 251398 399922 251454 399978
rect 251522 399922 251578 399978
rect 251646 399922 251702 399978
rect 239484 398402 239540 398458
rect 239372 392642 239428 392698
rect 229964 272042 230020 272098
rect 232540 373742 232596 373798
rect 230972 272042 231028 272098
rect 230972 265382 231028 265438
rect 235116 293822 235172 293878
rect 237804 311642 237860 311698
rect 238364 294722 238420 294778
rect 236796 294002 236852 294058
rect 236012 287342 236068 287398
rect 236236 285902 236292 285958
rect 236124 283922 236180 283978
rect 236348 270602 236404 270658
rect 236348 241622 236404 241678
rect 238588 376262 238644 376318
rect 250236 392282 250292 392338
rect 239708 294722 239764 294778
rect 239484 288782 239540 288838
rect 239596 292562 239652 292618
rect 239372 260342 239428 260398
rect 239484 285722 239540 285778
rect 239372 252062 239428 252118
rect 236684 231362 236740 231418
rect 236796 231182 236852 231238
rect 238476 227582 238532 227638
rect 233436 224162 233492 224218
rect 239820 293822 239876 293878
rect 239820 234602 239876 234658
rect 239932 288962 239988 289018
rect 240598 370294 240654 370350
rect 240722 370294 240778 370350
rect 240598 370170 240654 370226
rect 240722 370170 240778 370226
rect 240598 370046 240654 370102
rect 240722 370046 240778 370102
rect 240598 369922 240654 369978
rect 240722 369922 240778 369978
rect 240598 352294 240654 352350
rect 240722 352294 240778 352350
rect 240598 352170 240654 352226
rect 240722 352170 240778 352226
rect 240598 352046 240654 352102
rect 240722 352046 240778 352102
rect 240598 351922 240654 351978
rect 240722 351922 240778 351978
rect 240598 334294 240654 334350
rect 240722 334294 240778 334350
rect 240598 334170 240654 334226
rect 240722 334170 240778 334226
rect 240598 334046 240654 334102
rect 240722 334046 240778 334102
rect 240598 333922 240654 333978
rect 240722 333922 240778 333978
rect 240598 316294 240654 316350
rect 240722 316294 240778 316350
rect 240598 316170 240654 316226
rect 240722 316170 240778 316226
rect 240598 316046 240654 316102
rect 240722 316046 240778 316102
rect 240598 315922 240654 315978
rect 240722 315922 240778 315978
rect 240598 298294 240654 298350
rect 240722 298294 240778 298350
rect 240598 298170 240654 298226
rect 240722 298170 240778 298226
rect 240598 298046 240654 298102
rect 240722 298046 240778 298102
rect 240598 297922 240654 297978
rect 240722 297922 240778 297978
rect 240598 280294 240654 280350
rect 240722 280294 240778 280350
rect 240598 280170 240654 280226
rect 240722 280170 240778 280226
rect 240598 280046 240654 280102
rect 240722 280046 240778 280102
rect 240598 279922 240654 279978
rect 240722 279922 240778 279978
rect 240598 262294 240654 262350
rect 240722 262294 240778 262350
rect 240598 262170 240654 262226
rect 240722 262170 240778 262226
rect 240598 262046 240654 262102
rect 240722 262046 240778 262102
rect 240598 261922 240654 261978
rect 240722 261922 240778 261978
rect 241052 255482 241108 255538
rect 240598 244294 240654 244350
rect 240722 244294 240778 244350
rect 240598 244170 240654 244226
rect 240722 244170 240778 244226
rect 240598 244046 240654 244102
rect 240722 244046 240778 244102
rect 240598 243922 240654 243978
rect 240722 243922 240778 243978
rect 240044 227762 240100 227818
rect 239596 211382 239652 211438
rect 240156 211202 240212 211258
rect 241164 251162 241220 251218
rect 241164 241802 241220 241858
rect 251274 382294 251330 382350
rect 251398 382294 251454 382350
rect 251522 382294 251578 382350
rect 251646 382294 251702 382350
rect 251274 382170 251330 382226
rect 251398 382170 251454 382226
rect 251522 382170 251578 382226
rect 251646 382170 251702 382226
rect 251274 382046 251330 382102
rect 251398 382046 251454 382102
rect 251522 382046 251578 382102
rect 251646 382046 251702 382102
rect 251274 381922 251330 381978
rect 251398 381922 251454 381978
rect 251522 381922 251578 381978
rect 251646 381922 251702 381978
rect 254994 406294 255050 406350
rect 255118 406294 255174 406350
rect 255242 406294 255298 406350
rect 255366 406294 255422 406350
rect 254994 406170 255050 406226
rect 255118 406170 255174 406226
rect 255242 406170 255298 406226
rect 255366 406170 255422 406226
rect 254994 406046 255050 406102
rect 255118 406046 255174 406102
rect 255242 406046 255298 406102
rect 255366 406046 255422 406102
rect 254994 405922 255050 405978
rect 255118 405922 255174 405978
rect 255242 405922 255298 405978
rect 255366 405922 255422 405978
rect 267036 398942 267092 398998
rect 254994 388294 255050 388350
rect 255118 388294 255174 388350
rect 255242 388294 255298 388350
rect 255366 388294 255422 388350
rect 254994 388170 255050 388226
rect 255118 388170 255174 388226
rect 255242 388170 255298 388226
rect 255366 388170 255422 388226
rect 254994 388046 255050 388102
rect 255118 388046 255174 388102
rect 255242 388046 255298 388102
rect 255366 388046 255422 388102
rect 254994 387922 255050 387978
rect 255118 387922 255174 387978
rect 255242 387922 255298 387978
rect 255366 387922 255422 387978
rect 260316 392462 260372 392518
rect 281994 400294 282050 400350
rect 282118 400294 282174 400350
rect 282242 400294 282298 400350
rect 282366 400294 282422 400350
rect 281994 400170 282050 400226
rect 282118 400170 282174 400226
rect 282242 400170 282298 400226
rect 282366 400170 282422 400226
rect 281994 400046 282050 400102
rect 282118 400046 282174 400102
rect 282242 400046 282298 400102
rect 282366 400046 282422 400102
rect 281994 399922 282050 399978
rect 282118 399922 282174 399978
rect 282242 399922 282298 399978
rect 282366 399922 282422 399978
rect 281708 395522 281764 395578
rect 281994 382294 282050 382350
rect 282118 382294 282174 382350
rect 282242 382294 282298 382350
rect 282366 382294 282422 382350
rect 281994 382170 282050 382226
rect 282118 382170 282174 382226
rect 282242 382170 282298 382226
rect 282366 382170 282422 382226
rect 281994 382046 282050 382102
rect 282118 382046 282174 382102
rect 282242 382046 282298 382102
rect 282366 382046 282422 382102
rect 281994 381922 282050 381978
rect 282118 381922 282174 381978
rect 282242 381922 282298 381978
rect 282366 381922 282422 381978
rect 285714 406294 285770 406350
rect 285838 406294 285894 406350
rect 285962 406294 286018 406350
rect 286086 406294 286142 406350
rect 285714 406170 285770 406226
rect 285838 406170 285894 406226
rect 285962 406170 286018 406226
rect 286086 406170 286142 406226
rect 285714 406046 285770 406102
rect 285838 406046 285894 406102
rect 285962 406046 286018 406102
rect 286086 406046 286142 406102
rect 285714 405922 285770 405978
rect 285838 405922 285894 405978
rect 285962 405922 286018 405978
rect 286086 405922 286142 405978
rect 285714 388294 285770 388350
rect 285838 388294 285894 388350
rect 285962 388294 286018 388350
rect 286086 388294 286142 388350
rect 285714 388170 285770 388226
rect 285838 388170 285894 388226
rect 285962 388170 286018 388226
rect 286086 388170 286142 388226
rect 285714 388046 285770 388102
rect 285838 388046 285894 388102
rect 285962 388046 286018 388102
rect 286086 388046 286142 388102
rect 285714 387922 285770 387978
rect 285838 387922 285894 387978
rect 285962 387922 286018 387978
rect 286086 387922 286142 387978
rect 288092 407402 288148 407458
rect 291452 409382 291508 409438
rect 290556 405602 290612 405658
rect 295596 409022 295652 409078
rect 299852 407942 299908 407998
rect 293916 390842 293972 390898
rect 300636 407942 300692 407998
rect 301532 405422 301588 405478
rect 312714 400294 312770 400350
rect 312838 400294 312894 400350
rect 312962 400294 313018 400350
rect 313086 400294 313142 400350
rect 312714 400170 312770 400226
rect 312838 400170 312894 400226
rect 312962 400170 313018 400226
rect 313086 400170 313142 400226
rect 312714 400046 312770 400102
rect 312838 400046 312894 400102
rect 312962 400046 313018 400102
rect 313086 400046 313142 400102
rect 312714 399922 312770 399978
rect 312838 399922 312894 399978
rect 312962 399922 313018 399978
rect 313086 399922 313142 399978
rect 312396 396782 312452 396838
rect 316434 406294 316490 406350
rect 316558 406294 316614 406350
rect 316682 406294 316738 406350
rect 316806 406294 316862 406350
rect 316434 406170 316490 406226
rect 316558 406170 316614 406226
rect 316682 406170 316738 406226
rect 316806 406170 316862 406226
rect 316434 406046 316490 406102
rect 316558 406046 316614 406102
rect 316682 406046 316738 406102
rect 316806 406046 316862 406102
rect 316434 405922 316490 405978
rect 316558 405922 316614 405978
rect 316682 405922 316738 405978
rect 316806 405922 316862 405978
rect 312714 382294 312770 382350
rect 312838 382294 312894 382350
rect 312962 382294 313018 382350
rect 313086 382294 313142 382350
rect 312714 382170 312770 382226
rect 312838 382170 312894 382226
rect 312962 382170 313018 382226
rect 313086 382170 313142 382226
rect 312714 382046 312770 382102
rect 312838 382046 312894 382102
rect 312962 382046 313018 382102
rect 313086 382046 313142 382102
rect 299852 380762 299908 380818
rect 312714 381922 312770 381978
rect 312838 381922 312894 381978
rect 312962 381922 313018 381978
rect 313086 381922 313142 381978
rect 314076 396602 314132 396658
rect 315756 391022 315812 391078
rect 339612 407762 339668 407818
rect 316434 388294 316490 388350
rect 316558 388294 316614 388350
rect 316682 388294 316738 388350
rect 316806 388294 316862 388350
rect 316434 388170 316490 388226
rect 316558 388170 316614 388226
rect 316682 388170 316738 388226
rect 316806 388170 316862 388226
rect 316434 388046 316490 388102
rect 316558 388046 316614 388102
rect 316682 388046 316738 388102
rect 316806 388046 316862 388102
rect 316434 387922 316490 387978
rect 316558 387922 316614 387978
rect 316682 387922 316738 387978
rect 316806 387922 316862 387978
rect 315756 381302 315812 381358
rect 295596 380582 295652 380638
rect 280476 380402 280532 380458
rect 322588 390482 322644 390538
rect 338604 380582 338660 380638
rect 338492 380402 338548 380458
rect 271318 370294 271374 370350
rect 271442 370294 271498 370350
rect 271318 370170 271374 370226
rect 271442 370170 271498 370226
rect 271318 370046 271374 370102
rect 271442 370046 271498 370102
rect 271318 369922 271374 369978
rect 271442 369922 271498 369978
rect 302038 370294 302094 370350
rect 302162 370294 302218 370350
rect 302038 370170 302094 370226
rect 302162 370170 302218 370226
rect 302038 370046 302094 370102
rect 302162 370046 302218 370102
rect 302038 369922 302094 369978
rect 302162 369922 302218 369978
rect 332758 370294 332814 370350
rect 332882 370294 332938 370350
rect 332758 370170 332814 370226
rect 332882 370170 332938 370226
rect 332758 370046 332814 370102
rect 332882 370046 332938 370102
rect 332758 369922 332814 369978
rect 332882 369922 332938 369978
rect 255958 364294 256014 364350
rect 256082 364294 256138 364350
rect 255958 364170 256014 364226
rect 256082 364170 256138 364226
rect 255958 364046 256014 364102
rect 256082 364046 256138 364102
rect 255958 363922 256014 363978
rect 256082 363922 256138 363978
rect 286678 364294 286734 364350
rect 286802 364294 286858 364350
rect 286678 364170 286734 364226
rect 286802 364170 286858 364226
rect 286678 364046 286734 364102
rect 286802 364046 286858 364102
rect 286678 363922 286734 363978
rect 286802 363922 286858 363978
rect 317398 364294 317454 364350
rect 317522 364294 317578 364350
rect 317398 364170 317454 364226
rect 317522 364170 317578 364226
rect 317398 364046 317454 364102
rect 317522 364046 317578 364102
rect 317398 363922 317454 363978
rect 317522 363922 317578 363978
rect 271318 352294 271374 352350
rect 271442 352294 271498 352350
rect 271318 352170 271374 352226
rect 271442 352170 271498 352226
rect 271318 352046 271374 352102
rect 271442 352046 271498 352102
rect 271318 351922 271374 351978
rect 271442 351922 271498 351978
rect 302038 352294 302094 352350
rect 302162 352294 302218 352350
rect 302038 352170 302094 352226
rect 302162 352170 302218 352226
rect 302038 352046 302094 352102
rect 302162 352046 302218 352102
rect 302038 351922 302094 351978
rect 302162 351922 302218 351978
rect 332758 352294 332814 352350
rect 332882 352294 332938 352350
rect 332758 352170 332814 352226
rect 332882 352170 332938 352226
rect 332758 352046 332814 352102
rect 332882 352046 332938 352102
rect 332758 351922 332814 351978
rect 332882 351922 332938 351978
rect 255958 346294 256014 346350
rect 256082 346294 256138 346350
rect 255958 346170 256014 346226
rect 256082 346170 256138 346226
rect 255958 346046 256014 346102
rect 256082 346046 256138 346102
rect 255958 345922 256014 345978
rect 256082 345922 256138 345978
rect 286678 346294 286734 346350
rect 286802 346294 286858 346350
rect 286678 346170 286734 346226
rect 286802 346170 286858 346226
rect 286678 346046 286734 346102
rect 286802 346046 286858 346102
rect 286678 345922 286734 345978
rect 286802 345922 286858 345978
rect 317398 346294 317454 346350
rect 317522 346294 317578 346350
rect 317398 346170 317454 346226
rect 317522 346170 317578 346226
rect 317398 346046 317454 346102
rect 317522 346046 317578 346102
rect 317398 345922 317454 345978
rect 317522 345922 317578 345978
rect 338156 342422 338212 342478
rect 271318 334294 271374 334350
rect 271442 334294 271498 334350
rect 271318 334170 271374 334226
rect 271442 334170 271498 334226
rect 271318 334046 271374 334102
rect 271442 334046 271498 334102
rect 271318 333922 271374 333978
rect 271442 333922 271498 333978
rect 302038 334294 302094 334350
rect 302162 334294 302218 334350
rect 302038 334170 302094 334226
rect 302162 334170 302218 334226
rect 302038 334046 302094 334102
rect 302162 334046 302218 334102
rect 302038 333922 302094 333978
rect 302162 333922 302218 333978
rect 332758 334294 332814 334350
rect 332882 334294 332938 334350
rect 332758 334170 332814 334226
rect 332882 334170 332938 334226
rect 332758 334046 332814 334102
rect 332882 334046 332938 334102
rect 332758 333922 332814 333978
rect 332882 333922 332938 333978
rect 255958 328294 256014 328350
rect 256082 328294 256138 328350
rect 255958 328170 256014 328226
rect 256082 328170 256138 328226
rect 255958 328046 256014 328102
rect 256082 328046 256138 328102
rect 255958 327922 256014 327978
rect 256082 327922 256138 327978
rect 286678 328294 286734 328350
rect 286802 328294 286858 328350
rect 286678 328170 286734 328226
rect 286802 328170 286858 328226
rect 286678 328046 286734 328102
rect 286802 328046 286858 328102
rect 286678 327922 286734 327978
rect 286802 327922 286858 327978
rect 317398 328294 317454 328350
rect 317522 328294 317578 328350
rect 317398 328170 317454 328226
rect 317522 328170 317578 328226
rect 317398 328046 317454 328102
rect 317522 328046 317578 328102
rect 317398 327922 317454 327978
rect 317522 327922 317578 327978
rect 271318 316294 271374 316350
rect 271442 316294 271498 316350
rect 271318 316170 271374 316226
rect 271442 316170 271498 316226
rect 271318 316046 271374 316102
rect 271442 316046 271498 316102
rect 271318 315922 271374 315978
rect 271442 315922 271498 315978
rect 302038 316294 302094 316350
rect 302162 316294 302218 316350
rect 302038 316170 302094 316226
rect 302162 316170 302218 316226
rect 302038 316046 302094 316102
rect 302162 316046 302218 316102
rect 302038 315922 302094 315978
rect 302162 315922 302218 315978
rect 332758 316294 332814 316350
rect 332882 316294 332938 316350
rect 332758 316170 332814 316226
rect 332882 316170 332938 316226
rect 332758 316046 332814 316102
rect 332882 316046 332938 316102
rect 332758 315922 332814 315978
rect 332882 315922 332938 315978
rect 255958 310294 256014 310350
rect 256082 310294 256138 310350
rect 255958 310170 256014 310226
rect 256082 310170 256138 310226
rect 255958 310046 256014 310102
rect 256082 310046 256138 310102
rect 255958 309922 256014 309978
rect 256082 309922 256138 309978
rect 286678 310294 286734 310350
rect 286802 310294 286858 310350
rect 286678 310170 286734 310226
rect 286802 310170 286858 310226
rect 286678 310046 286734 310102
rect 286802 310046 286858 310102
rect 286678 309922 286734 309978
rect 286802 309922 286858 309978
rect 317398 310294 317454 310350
rect 317522 310294 317578 310350
rect 317398 310170 317454 310226
rect 317522 310170 317578 310226
rect 317398 310046 317454 310102
rect 317522 310046 317578 310102
rect 317398 309922 317454 309978
rect 317522 309922 317578 309978
rect 271318 298294 271374 298350
rect 271442 298294 271498 298350
rect 271318 298170 271374 298226
rect 271442 298170 271498 298226
rect 271318 298046 271374 298102
rect 271442 298046 271498 298102
rect 271318 297922 271374 297978
rect 271442 297922 271498 297978
rect 302038 298294 302094 298350
rect 302162 298294 302218 298350
rect 302038 298170 302094 298226
rect 302162 298170 302218 298226
rect 302038 298046 302094 298102
rect 302162 298046 302218 298102
rect 302038 297922 302094 297978
rect 302162 297922 302218 297978
rect 332758 298294 332814 298350
rect 332882 298294 332938 298350
rect 332758 298170 332814 298226
rect 332882 298170 332938 298226
rect 332758 298046 332814 298102
rect 332882 298046 332938 298102
rect 332758 297922 332814 297978
rect 332882 297922 332938 297978
rect 255958 292294 256014 292350
rect 256082 292294 256138 292350
rect 255958 292170 256014 292226
rect 256082 292170 256138 292226
rect 255958 292046 256014 292102
rect 256082 292046 256138 292102
rect 255958 291922 256014 291978
rect 256082 291922 256138 291978
rect 286678 292294 286734 292350
rect 286802 292294 286858 292350
rect 286678 292170 286734 292226
rect 286802 292170 286858 292226
rect 286678 292046 286734 292102
rect 286802 292046 286858 292102
rect 286678 291922 286734 291978
rect 286802 291922 286858 291978
rect 317398 292294 317454 292350
rect 317522 292294 317578 292350
rect 317398 292170 317454 292226
rect 317522 292170 317578 292226
rect 317398 292046 317454 292102
rect 317522 292046 317578 292102
rect 317398 291922 317454 291978
rect 317522 291922 317578 291978
rect 271318 280294 271374 280350
rect 271442 280294 271498 280350
rect 271318 280170 271374 280226
rect 271442 280170 271498 280226
rect 271318 280046 271374 280102
rect 271442 280046 271498 280102
rect 271318 279922 271374 279978
rect 271442 279922 271498 279978
rect 302038 280294 302094 280350
rect 302162 280294 302218 280350
rect 302038 280170 302094 280226
rect 302162 280170 302218 280226
rect 302038 280046 302094 280102
rect 302162 280046 302218 280102
rect 302038 279922 302094 279978
rect 302162 279922 302218 279978
rect 332758 280294 332814 280350
rect 332882 280294 332938 280350
rect 332758 280170 332814 280226
rect 332882 280170 332938 280226
rect 332758 280046 332814 280102
rect 332882 280046 332938 280102
rect 332758 279922 332814 279978
rect 332882 279922 332938 279978
rect 255958 274294 256014 274350
rect 256082 274294 256138 274350
rect 255958 274170 256014 274226
rect 256082 274170 256138 274226
rect 255958 274046 256014 274102
rect 256082 274046 256138 274102
rect 255958 273922 256014 273978
rect 256082 273922 256138 273978
rect 286678 274294 286734 274350
rect 286802 274294 286858 274350
rect 286678 274170 286734 274226
rect 286802 274170 286858 274226
rect 286678 274046 286734 274102
rect 286802 274046 286858 274102
rect 286678 273922 286734 273978
rect 286802 273922 286858 273978
rect 317398 274294 317454 274350
rect 317522 274294 317578 274350
rect 317398 274170 317454 274226
rect 317522 274170 317578 274226
rect 317398 274046 317454 274102
rect 317522 274046 317578 274102
rect 317398 273922 317454 273978
rect 317522 273922 317578 273978
rect 271318 262294 271374 262350
rect 271442 262294 271498 262350
rect 271318 262170 271374 262226
rect 271442 262170 271498 262226
rect 271318 262046 271374 262102
rect 271442 262046 271498 262102
rect 271318 261922 271374 261978
rect 271442 261922 271498 261978
rect 302038 262294 302094 262350
rect 302162 262294 302218 262350
rect 302038 262170 302094 262226
rect 302162 262170 302218 262226
rect 302038 262046 302094 262102
rect 302162 262046 302218 262102
rect 302038 261922 302094 261978
rect 302162 261922 302218 261978
rect 332758 262294 332814 262350
rect 332882 262294 332938 262350
rect 332758 262170 332814 262226
rect 332882 262170 332938 262226
rect 332758 262046 332814 262102
rect 332882 262046 332938 262102
rect 332758 261922 332814 261978
rect 332882 261922 332938 261978
rect 255958 256294 256014 256350
rect 256082 256294 256138 256350
rect 255958 256170 256014 256226
rect 256082 256170 256138 256226
rect 255958 256046 256014 256102
rect 256082 256046 256138 256102
rect 255958 255922 256014 255978
rect 256082 255922 256138 255978
rect 286678 256294 286734 256350
rect 286802 256294 286858 256350
rect 286678 256170 286734 256226
rect 286802 256170 286858 256226
rect 286678 256046 286734 256102
rect 286802 256046 286858 256102
rect 286678 255922 286734 255978
rect 286802 255922 286858 255978
rect 317398 256294 317454 256350
rect 317522 256294 317578 256350
rect 317398 256170 317454 256226
rect 317522 256170 317578 256226
rect 317398 256046 317454 256102
rect 317522 256046 317578 256102
rect 317398 255922 317454 255978
rect 317522 255922 317578 255978
rect 339276 342422 339332 342478
rect 338268 301922 338324 301978
rect 339388 301922 339444 301978
rect 338380 253682 338436 253738
rect 337932 244862 337988 244918
rect 338380 249902 338436 249958
rect 271318 244294 271374 244350
rect 271442 244294 271498 244350
rect 271318 244170 271374 244226
rect 271442 244170 271498 244226
rect 271318 244046 271374 244102
rect 271442 244046 271498 244102
rect 271318 243922 271374 243978
rect 271442 243922 271498 243978
rect 302038 244294 302094 244350
rect 302162 244294 302218 244350
rect 302038 244170 302094 244226
rect 302162 244170 302218 244226
rect 302038 244046 302094 244102
rect 302162 244046 302218 244102
rect 302038 243922 302094 243978
rect 302162 243922 302218 243978
rect 332758 244294 332814 244350
rect 332882 244294 332938 244350
rect 332758 244170 332814 244226
rect 332882 244170 332938 244226
rect 332758 244046 332814 244102
rect 332882 244046 332938 244102
rect 332758 243922 332814 243978
rect 332882 243922 332938 243978
rect 336924 241442 336980 241498
rect 289772 241082 289828 241138
rect 241836 227942 241892 227998
rect 245084 237122 245140 237178
rect 251274 238294 251330 238350
rect 251398 238294 251454 238350
rect 251522 238294 251578 238350
rect 251646 238294 251702 238350
rect 251274 238170 251330 238226
rect 251398 238170 251454 238226
rect 251522 238170 251578 238226
rect 251646 238170 251702 238226
rect 251274 238046 251330 238102
rect 251398 238046 251454 238102
rect 251522 238046 251578 238102
rect 251646 238046 251702 238102
rect 251274 237922 251330 237978
rect 251398 237922 251454 237978
rect 251522 237922 251578 237978
rect 251646 237922 251702 237978
rect 243404 224522 243460 224578
rect 244188 236942 244244 236998
rect 243516 224342 243572 224398
rect 241052 211022 241108 211078
rect 269836 237122 269892 237178
rect 251274 220294 251330 220350
rect 251398 220294 251454 220350
rect 251522 220294 251578 220350
rect 251646 220294 251702 220350
rect 251274 220170 251330 220226
rect 251398 220170 251454 220226
rect 251522 220170 251578 220226
rect 251646 220170 251702 220226
rect 251274 220046 251330 220102
rect 251398 220046 251454 220102
rect 251522 220046 251578 220102
rect 251646 220046 251702 220102
rect 251274 219922 251330 219978
rect 251398 219922 251454 219978
rect 251522 219922 251578 219978
rect 251646 219922 251702 219978
rect 44518 202294 44574 202350
rect 44642 202294 44698 202350
rect 44518 202170 44574 202226
rect 44642 202170 44698 202226
rect 44518 202046 44574 202102
rect 44642 202046 44698 202102
rect 44518 201922 44574 201978
rect 44642 201922 44698 201978
rect 75238 202294 75294 202350
rect 75362 202294 75418 202350
rect 75238 202170 75294 202226
rect 75362 202170 75418 202226
rect 75238 202046 75294 202102
rect 75362 202046 75418 202102
rect 75238 201922 75294 201978
rect 75362 201922 75418 201978
rect 105958 202294 106014 202350
rect 106082 202294 106138 202350
rect 105958 202170 106014 202226
rect 106082 202170 106138 202226
rect 105958 202046 106014 202102
rect 106082 202046 106138 202102
rect 105958 201922 106014 201978
rect 106082 201922 106138 201978
rect 136678 202294 136734 202350
rect 136802 202294 136858 202350
rect 136678 202170 136734 202226
rect 136802 202170 136858 202226
rect 136678 202046 136734 202102
rect 136802 202046 136858 202102
rect 136678 201922 136734 201978
rect 136802 201922 136858 201978
rect 167398 202294 167454 202350
rect 167522 202294 167578 202350
rect 167398 202170 167454 202226
rect 167522 202170 167578 202226
rect 167398 202046 167454 202102
rect 167522 202046 167578 202102
rect 167398 201922 167454 201978
rect 167522 201922 167578 201978
rect 198118 202294 198174 202350
rect 198242 202294 198298 202350
rect 198118 202170 198174 202226
rect 198242 202170 198298 202226
rect 198118 202046 198174 202102
rect 198242 202046 198298 202102
rect 198118 201922 198174 201978
rect 198242 201922 198298 201978
rect 228838 202294 228894 202350
rect 228962 202294 229018 202350
rect 228838 202170 228894 202226
rect 228962 202170 229018 202226
rect 228838 202046 228894 202102
rect 228962 202046 229018 202102
rect 228838 201922 228894 201978
rect 228962 201922 229018 201978
rect 259558 202294 259614 202350
rect 259682 202294 259738 202350
rect 259558 202170 259614 202226
rect 259682 202170 259738 202226
rect 259558 202046 259614 202102
rect 259682 202046 259738 202102
rect 259558 201922 259614 201978
rect 259682 201922 259738 201978
rect 59878 190294 59934 190350
rect 60002 190294 60058 190350
rect 59878 190170 59934 190226
rect 60002 190170 60058 190226
rect 59878 190046 59934 190102
rect 60002 190046 60058 190102
rect 59878 189922 59934 189978
rect 60002 189922 60058 189978
rect 90598 190294 90654 190350
rect 90722 190294 90778 190350
rect 90598 190170 90654 190226
rect 90722 190170 90778 190226
rect 90598 190046 90654 190102
rect 90722 190046 90778 190102
rect 90598 189922 90654 189978
rect 90722 189922 90778 189978
rect 121318 190294 121374 190350
rect 121442 190294 121498 190350
rect 121318 190170 121374 190226
rect 121442 190170 121498 190226
rect 121318 190046 121374 190102
rect 121442 190046 121498 190102
rect 121318 189922 121374 189978
rect 121442 189922 121498 189978
rect 152038 190294 152094 190350
rect 152162 190294 152218 190350
rect 152038 190170 152094 190226
rect 152162 190170 152218 190226
rect 152038 190046 152094 190102
rect 152162 190046 152218 190102
rect 152038 189922 152094 189978
rect 152162 189922 152218 189978
rect 182758 190294 182814 190350
rect 182882 190294 182938 190350
rect 182758 190170 182814 190226
rect 182882 190170 182938 190226
rect 182758 190046 182814 190102
rect 182882 190046 182938 190102
rect 182758 189922 182814 189978
rect 182882 189922 182938 189978
rect 213478 190294 213534 190350
rect 213602 190294 213658 190350
rect 213478 190170 213534 190226
rect 213602 190170 213658 190226
rect 213478 190046 213534 190102
rect 213602 190046 213658 190102
rect 213478 189922 213534 189978
rect 213602 189922 213658 189978
rect 244198 190294 244254 190350
rect 244322 190294 244378 190350
rect 244198 190170 244254 190226
rect 244322 190170 244378 190226
rect 244198 190046 244254 190102
rect 244322 190046 244378 190102
rect 244198 189922 244254 189978
rect 244322 189922 244378 189978
rect 44518 184294 44574 184350
rect 44642 184294 44698 184350
rect 44518 184170 44574 184226
rect 44642 184170 44698 184226
rect 44518 184046 44574 184102
rect 44642 184046 44698 184102
rect 44518 183922 44574 183978
rect 44642 183922 44698 183978
rect 75238 184294 75294 184350
rect 75362 184294 75418 184350
rect 75238 184170 75294 184226
rect 75362 184170 75418 184226
rect 75238 184046 75294 184102
rect 75362 184046 75418 184102
rect 75238 183922 75294 183978
rect 75362 183922 75418 183978
rect 105958 184294 106014 184350
rect 106082 184294 106138 184350
rect 105958 184170 106014 184226
rect 106082 184170 106138 184226
rect 105958 184046 106014 184102
rect 106082 184046 106138 184102
rect 105958 183922 106014 183978
rect 106082 183922 106138 183978
rect 136678 184294 136734 184350
rect 136802 184294 136858 184350
rect 136678 184170 136734 184226
rect 136802 184170 136858 184226
rect 136678 184046 136734 184102
rect 136802 184046 136858 184102
rect 136678 183922 136734 183978
rect 136802 183922 136858 183978
rect 167398 184294 167454 184350
rect 167522 184294 167578 184350
rect 167398 184170 167454 184226
rect 167522 184170 167578 184226
rect 167398 184046 167454 184102
rect 167522 184046 167578 184102
rect 167398 183922 167454 183978
rect 167522 183922 167578 183978
rect 198118 184294 198174 184350
rect 198242 184294 198298 184350
rect 198118 184170 198174 184226
rect 198242 184170 198298 184226
rect 198118 184046 198174 184102
rect 198242 184046 198298 184102
rect 198118 183922 198174 183978
rect 198242 183922 198298 183978
rect 228838 184294 228894 184350
rect 228962 184294 229018 184350
rect 228838 184170 228894 184226
rect 228962 184170 229018 184226
rect 228838 184046 228894 184102
rect 228962 184046 229018 184102
rect 228838 183922 228894 183978
rect 228962 183922 229018 183978
rect 259558 184294 259614 184350
rect 259682 184294 259738 184350
rect 259558 184170 259614 184226
rect 259682 184170 259738 184226
rect 259558 184046 259614 184102
rect 259682 184046 259738 184102
rect 259558 183922 259614 183978
rect 259682 183922 259738 183978
rect 59878 172294 59934 172350
rect 60002 172294 60058 172350
rect 59878 172170 59934 172226
rect 60002 172170 60058 172226
rect 59878 172046 59934 172102
rect 60002 172046 60058 172102
rect 59878 171922 59934 171978
rect 60002 171922 60058 171978
rect 90598 172294 90654 172350
rect 90722 172294 90778 172350
rect 90598 172170 90654 172226
rect 90722 172170 90778 172226
rect 90598 172046 90654 172102
rect 90722 172046 90778 172102
rect 90598 171922 90654 171978
rect 90722 171922 90778 171978
rect 121318 172294 121374 172350
rect 121442 172294 121498 172350
rect 121318 172170 121374 172226
rect 121442 172170 121498 172226
rect 121318 172046 121374 172102
rect 121442 172046 121498 172102
rect 121318 171922 121374 171978
rect 121442 171922 121498 171978
rect 152038 172294 152094 172350
rect 152162 172294 152218 172350
rect 152038 172170 152094 172226
rect 152162 172170 152218 172226
rect 152038 172046 152094 172102
rect 152162 172046 152218 172102
rect 152038 171922 152094 171978
rect 152162 171922 152218 171978
rect 182758 172294 182814 172350
rect 182882 172294 182938 172350
rect 182758 172170 182814 172226
rect 182882 172170 182938 172226
rect 182758 172046 182814 172102
rect 182882 172046 182938 172102
rect 182758 171922 182814 171978
rect 182882 171922 182938 171978
rect 213478 172294 213534 172350
rect 213602 172294 213658 172350
rect 213478 172170 213534 172226
rect 213602 172170 213658 172226
rect 213478 172046 213534 172102
rect 213602 172046 213658 172102
rect 213478 171922 213534 171978
rect 213602 171922 213658 171978
rect 244198 172294 244254 172350
rect 244322 172294 244378 172350
rect 244198 172170 244254 172226
rect 244322 172170 244378 172226
rect 244198 172046 244254 172102
rect 244322 172046 244378 172102
rect 244198 171922 244254 171978
rect 244322 171922 244378 171978
rect 44518 166294 44574 166350
rect 44642 166294 44698 166350
rect 44518 166170 44574 166226
rect 44642 166170 44698 166226
rect 44518 166046 44574 166102
rect 44642 166046 44698 166102
rect 44518 165922 44574 165978
rect 44642 165922 44698 165978
rect 75238 166294 75294 166350
rect 75362 166294 75418 166350
rect 75238 166170 75294 166226
rect 75362 166170 75418 166226
rect 75238 166046 75294 166102
rect 75362 166046 75418 166102
rect 75238 165922 75294 165978
rect 75362 165922 75418 165978
rect 105958 166294 106014 166350
rect 106082 166294 106138 166350
rect 105958 166170 106014 166226
rect 106082 166170 106138 166226
rect 105958 166046 106014 166102
rect 106082 166046 106138 166102
rect 105958 165922 106014 165978
rect 106082 165922 106138 165978
rect 136678 166294 136734 166350
rect 136802 166294 136858 166350
rect 136678 166170 136734 166226
rect 136802 166170 136858 166226
rect 136678 166046 136734 166102
rect 136802 166046 136858 166102
rect 136678 165922 136734 165978
rect 136802 165922 136858 165978
rect 167398 166294 167454 166350
rect 167522 166294 167578 166350
rect 167398 166170 167454 166226
rect 167522 166170 167578 166226
rect 167398 166046 167454 166102
rect 167522 166046 167578 166102
rect 167398 165922 167454 165978
rect 167522 165922 167578 165978
rect 198118 166294 198174 166350
rect 198242 166294 198298 166350
rect 198118 166170 198174 166226
rect 198242 166170 198298 166226
rect 198118 166046 198174 166102
rect 198242 166046 198298 166102
rect 198118 165922 198174 165978
rect 198242 165922 198298 165978
rect 228838 166294 228894 166350
rect 228962 166294 229018 166350
rect 228838 166170 228894 166226
rect 228962 166170 229018 166226
rect 228838 166046 228894 166102
rect 228962 166046 229018 166102
rect 228838 165922 228894 165978
rect 228962 165922 229018 165978
rect 259558 166294 259614 166350
rect 259682 166294 259738 166350
rect 259558 166170 259614 166226
rect 259682 166170 259738 166226
rect 259558 166046 259614 166102
rect 259682 166046 259738 166102
rect 259558 165922 259614 165978
rect 259682 165922 259738 165978
rect 59878 154294 59934 154350
rect 60002 154294 60058 154350
rect 59878 154170 59934 154226
rect 60002 154170 60058 154226
rect 59878 154046 59934 154102
rect 60002 154046 60058 154102
rect 59878 153922 59934 153978
rect 60002 153922 60058 153978
rect 90598 154294 90654 154350
rect 90722 154294 90778 154350
rect 90598 154170 90654 154226
rect 90722 154170 90778 154226
rect 90598 154046 90654 154102
rect 90722 154046 90778 154102
rect 90598 153922 90654 153978
rect 90722 153922 90778 153978
rect 121318 154294 121374 154350
rect 121442 154294 121498 154350
rect 121318 154170 121374 154226
rect 121442 154170 121498 154226
rect 121318 154046 121374 154102
rect 121442 154046 121498 154102
rect 121318 153922 121374 153978
rect 121442 153922 121498 153978
rect 152038 154294 152094 154350
rect 152162 154294 152218 154350
rect 152038 154170 152094 154226
rect 152162 154170 152218 154226
rect 152038 154046 152094 154102
rect 152162 154046 152218 154102
rect 152038 153922 152094 153978
rect 152162 153922 152218 153978
rect 182758 154294 182814 154350
rect 182882 154294 182938 154350
rect 182758 154170 182814 154226
rect 182882 154170 182938 154226
rect 182758 154046 182814 154102
rect 182882 154046 182938 154102
rect 182758 153922 182814 153978
rect 182882 153922 182938 153978
rect 213478 154294 213534 154350
rect 213602 154294 213658 154350
rect 213478 154170 213534 154226
rect 213602 154170 213658 154226
rect 213478 154046 213534 154102
rect 213602 154046 213658 154102
rect 213478 153922 213534 153978
rect 213602 153922 213658 153978
rect 244198 154294 244254 154350
rect 244322 154294 244378 154350
rect 244198 154170 244254 154226
rect 244322 154170 244378 154226
rect 244198 154046 244254 154102
rect 244322 154046 244378 154102
rect 244198 153922 244254 153978
rect 244322 153922 244378 153978
rect 44518 148294 44574 148350
rect 44642 148294 44698 148350
rect 44518 148170 44574 148226
rect 44642 148170 44698 148226
rect 44518 148046 44574 148102
rect 44642 148046 44698 148102
rect 44518 147922 44574 147978
rect 44642 147922 44698 147978
rect 75238 148294 75294 148350
rect 75362 148294 75418 148350
rect 75238 148170 75294 148226
rect 75362 148170 75418 148226
rect 75238 148046 75294 148102
rect 75362 148046 75418 148102
rect 75238 147922 75294 147978
rect 75362 147922 75418 147978
rect 105958 148294 106014 148350
rect 106082 148294 106138 148350
rect 105958 148170 106014 148226
rect 106082 148170 106138 148226
rect 105958 148046 106014 148102
rect 106082 148046 106138 148102
rect 105958 147922 106014 147978
rect 106082 147922 106138 147978
rect 136678 148294 136734 148350
rect 136802 148294 136858 148350
rect 136678 148170 136734 148226
rect 136802 148170 136858 148226
rect 136678 148046 136734 148102
rect 136802 148046 136858 148102
rect 136678 147922 136734 147978
rect 136802 147922 136858 147978
rect 167398 148294 167454 148350
rect 167522 148294 167578 148350
rect 167398 148170 167454 148226
rect 167522 148170 167578 148226
rect 167398 148046 167454 148102
rect 167522 148046 167578 148102
rect 167398 147922 167454 147978
rect 167522 147922 167578 147978
rect 198118 148294 198174 148350
rect 198242 148294 198298 148350
rect 198118 148170 198174 148226
rect 198242 148170 198298 148226
rect 198118 148046 198174 148102
rect 198242 148046 198298 148102
rect 198118 147922 198174 147978
rect 198242 147922 198298 147978
rect 228838 148294 228894 148350
rect 228962 148294 229018 148350
rect 228838 148170 228894 148226
rect 228962 148170 229018 148226
rect 228838 148046 228894 148102
rect 228962 148046 229018 148102
rect 228838 147922 228894 147978
rect 228962 147922 229018 147978
rect 259558 148294 259614 148350
rect 259682 148294 259738 148350
rect 259558 148170 259614 148226
rect 259682 148170 259738 148226
rect 259558 148046 259614 148102
rect 259682 148046 259738 148102
rect 259558 147922 259614 147978
rect 259682 147922 259738 147978
rect 59878 136294 59934 136350
rect 60002 136294 60058 136350
rect 59878 136170 59934 136226
rect 60002 136170 60058 136226
rect 59878 136046 59934 136102
rect 60002 136046 60058 136102
rect 59878 135922 59934 135978
rect 60002 135922 60058 135978
rect 90598 136294 90654 136350
rect 90722 136294 90778 136350
rect 90598 136170 90654 136226
rect 90722 136170 90778 136226
rect 90598 136046 90654 136102
rect 90722 136046 90778 136102
rect 90598 135922 90654 135978
rect 90722 135922 90778 135978
rect 121318 136294 121374 136350
rect 121442 136294 121498 136350
rect 121318 136170 121374 136226
rect 121442 136170 121498 136226
rect 121318 136046 121374 136102
rect 121442 136046 121498 136102
rect 121318 135922 121374 135978
rect 121442 135922 121498 135978
rect 152038 136294 152094 136350
rect 152162 136294 152218 136350
rect 152038 136170 152094 136226
rect 152162 136170 152218 136226
rect 152038 136046 152094 136102
rect 152162 136046 152218 136102
rect 152038 135922 152094 135978
rect 152162 135922 152218 135978
rect 182758 136294 182814 136350
rect 182882 136294 182938 136350
rect 182758 136170 182814 136226
rect 182882 136170 182938 136226
rect 182758 136046 182814 136102
rect 182882 136046 182938 136102
rect 182758 135922 182814 135978
rect 182882 135922 182938 135978
rect 213478 136294 213534 136350
rect 213602 136294 213658 136350
rect 213478 136170 213534 136226
rect 213602 136170 213658 136226
rect 213478 136046 213534 136102
rect 213602 136046 213658 136102
rect 213478 135922 213534 135978
rect 213602 135922 213658 135978
rect 244198 136294 244254 136350
rect 244322 136294 244378 136350
rect 244198 136170 244254 136226
rect 244322 136170 244378 136226
rect 244198 136046 244254 136102
rect 244322 136046 244378 136102
rect 244198 135922 244254 135978
rect 244322 135922 244378 135978
rect 44518 130294 44574 130350
rect 44642 130294 44698 130350
rect 44518 130170 44574 130226
rect 44642 130170 44698 130226
rect 44518 130046 44574 130102
rect 44642 130046 44698 130102
rect 44518 129922 44574 129978
rect 44642 129922 44698 129978
rect 75238 130294 75294 130350
rect 75362 130294 75418 130350
rect 75238 130170 75294 130226
rect 75362 130170 75418 130226
rect 75238 130046 75294 130102
rect 75362 130046 75418 130102
rect 75238 129922 75294 129978
rect 75362 129922 75418 129978
rect 105958 130294 106014 130350
rect 106082 130294 106138 130350
rect 105958 130170 106014 130226
rect 106082 130170 106138 130226
rect 105958 130046 106014 130102
rect 106082 130046 106138 130102
rect 105958 129922 106014 129978
rect 106082 129922 106138 129978
rect 136678 130294 136734 130350
rect 136802 130294 136858 130350
rect 136678 130170 136734 130226
rect 136802 130170 136858 130226
rect 136678 130046 136734 130102
rect 136802 130046 136858 130102
rect 136678 129922 136734 129978
rect 136802 129922 136858 129978
rect 167398 130294 167454 130350
rect 167522 130294 167578 130350
rect 167398 130170 167454 130226
rect 167522 130170 167578 130226
rect 167398 130046 167454 130102
rect 167522 130046 167578 130102
rect 167398 129922 167454 129978
rect 167522 129922 167578 129978
rect 198118 130294 198174 130350
rect 198242 130294 198298 130350
rect 198118 130170 198174 130226
rect 198242 130170 198298 130226
rect 198118 130046 198174 130102
rect 198242 130046 198298 130102
rect 198118 129922 198174 129978
rect 198242 129922 198298 129978
rect 228838 130294 228894 130350
rect 228962 130294 229018 130350
rect 228838 130170 228894 130226
rect 228962 130170 229018 130226
rect 228838 130046 228894 130102
rect 228962 130046 229018 130102
rect 228838 129922 228894 129978
rect 228962 129922 229018 129978
rect 259558 130294 259614 130350
rect 259682 130294 259738 130350
rect 259558 130170 259614 130226
rect 259682 130170 259738 130226
rect 259558 130046 259614 130102
rect 259682 130046 259738 130102
rect 259558 129922 259614 129978
rect 259682 129922 259738 129978
rect 59878 118294 59934 118350
rect 60002 118294 60058 118350
rect 59878 118170 59934 118226
rect 60002 118170 60058 118226
rect 59878 118046 59934 118102
rect 60002 118046 60058 118102
rect 59878 117922 59934 117978
rect 60002 117922 60058 117978
rect 90598 118294 90654 118350
rect 90722 118294 90778 118350
rect 90598 118170 90654 118226
rect 90722 118170 90778 118226
rect 90598 118046 90654 118102
rect 90722 118046 90778 118102
rect 90598 117922 90654 117978
rect 90722 117922 90778 117978
rect 121318 118294 121374 118350
rect 121442 118294 121498 118350
rect 121318 118170 121374 118226
rect 121442 118170 121498 118226
rect 121318 118046 121374 118102
rect 121442 118046 121498 118102
rect 121318 117922 121374 117978
rect 121442 117922 121498 117978
rect 152038 118294 152094 118350
rect 152162 118294 152218 118350
rect 152038 118170 152094 118226
rect 152162 118170 152218 118226
rect 152038 118046 152094 118102
rect 152162 118046 152218 118102
rect 152038 117922 152094 117978
rect 152162 117922 152218 117978
rect 182758 118294 182814 118350
rect 182882 118294 182938 118350
rect 182758 118170 182814 118226
rect 182882 118170 182938 118226
rect 182758 118046 182814 118102
rect 182882 118046 182938 118102
rect 182758 117922 182814 117978
rect 182882 117922 182938 117978
rect 213478 118294 213534 118350
rect 213602 118294 213658 118350
rect 213478 118170 213534 118226
rect 213602 118170 213658 118226
rect 213478 118046 213534 118102
rect 213602 118046 213658 118102
rect 213478 117922 213534 117978
rect 213602 117922 213658 117978
rect 244198 118294 244254 118350
rect 244322 118294 244378 118350
rect 244198 118170 244254 118226
rect 244322 118170 244378 118226
rect 244198 118046 244254 118102
rect 244322 118046 244378 118102
rect 244198 117922 244254 117978
rect 244322 117922 244378 117978
rect 44518 112294 44574 112350
rect 44642 112294 44698 112350
rect 44518 112170 44574 112226
rect 44642 112170 44698 112226
rect 44518 112046 44574 112102
rect 44642 112046 44698 112102
rect 44518 111922 44574 111978
rect 44642 111922 44698 111978
rect 75238 112294 75294 112350
rect 75362 112294 75418 112350
rect 75238 112170 75294 112226
rect 75362 112170 75418 112226
rect 75238 112046 75294 112102
rect 75362 112046 75418 112102
rect 75238 111922 75294 111978
rect 75362 111922 75418 111978
rect 105958 112294 106014 112350
rect 106082 112294 106138 112350
rect 105958 112170 106014 112226
rect 106082 112170 106138 112226
rect 105958 112046 106014 112102
rect 106082 112046 106138 112102
rect 105958 111922 106014 111978
rect 106082 111922 106138 111978
rect 136678 112294 136734 112350
rect 136802 112294 136858 112350
rect 136678 112170 136734 112226
rect 136802 112170 136858 112226
rect 136678 112046 136734 112102
rect 136802 112046 136858 112102
rect 136678 111922 136734 111978
rect 136802 111922 136858 111978
rect 167398 112294 167454 112350
rect 167522 112294 167578 112350
rect 167398 112170 167454 112226
rect 167522 112170 167578 112226
rect 167398 112046 167454 112102
rect 167522 112046 167578 112102
rect 167398 111922 167454 111978
rect 167522 111922 167578 111978
rect 198118 112294 198174 112350
rect 198242 112294 198298 112350
rect 198118 112170 198174 112226
rect 198242 112170 198298 112226
rect 198118 112046 198174 112102
rect 198242 112046 198298 112102
rect 198118 111922 198174 111978
rect 198242 111922 198298 111978
rect 228838 112294 228894 112350
rect 228962 112294 229018 112350
rect 228838 112170 228894 112226
rect 228962 112170 229018 112226
rect 228838 112046 228894 112102
rect 228962 112046 229018 112102
rect 228838 111922 228894 111978
rect 228962 111922 229018 111978
rect 259558 112294 259614 112350
rect 259682 112294 259738 112350
rect 259558 112170 259614 112226
rect 259682 112170 259738 112226
rect 259558 112046 259614 112102
rect 259682 112046 259738 112102
rect 259558 111922 259614 111978
rect 259682 111922 259738 111978
rect 59878 100294 59934 100350
rect 60002 100294 60058 100350
rect 59878 100170 59934 100226
rect 60002 100170 60058 100226
rect 59878 100046 59934 100102
rect 60002 100046 60058 100102
rect 59878 99922 59934 99978
rect 60002 99922 60058 99978
rect 90598 100294 90654 100350
rect 90722 100294 90778 100350
rect 90598 100170 90654 100226
rect 90722 100170 90778 100226
rect 90598 100046 90654 100102
rect 90722 100046 90778 100102
rect 90598 99922 90654 99978
rect 90722 99922 90778 99978
rect 121318 100294 121374 100350
rect 121442 100294 121498 100350
rect 121318 100170 121374 100226
rect 121442 100170 121498 100226
rect 121318 100046 121374 100102
rect 121442 100046 121498 100102
rect 121318 99922 121374 99978
rect 121442 99922 121498 99978
rect 152038 100294 152094 100350
rect 152162 100294 152218 100350
rect 152038 100170 152094 100226
rect 152162 100170 152218 100226
rect 152038 100046 152094 100102
rect 152162 100046 152218 100102
rect 152038 99922 152094 99978
rect 152162 99922 152218 99978
rect 182758 100294 182814 100350
rect 182882 100294 182938 100350
rect 182758 100170 182814 100226
rect 182882 100170 182938 100226
rect 182758 100046 182814 100102
rect 182882 100046 182938 100102
rect 182758 99922 182814 99978
rect 182882 99922 182938 99978
rect 213478 100294 213534 100350
rect 213602 100294 213658 100350
rect 213478 100170 213534 100226
rect 213602 100170 213658 100226
rect 213478 100046 213534 100102
rect 213602 100046 213658 100102
rect 213478 99922 213534 99978
rect 213602 99922 213658 99978
rect 244198 100294 244254 100350
rect 244322 100294 244378 100350
rect 244198 100170 244254 100226
rect 244322 100170 244378 100226
rect 244198 100046 244254 100102
rect 244322 100046 244378 100102
rect 244198 99922 244254 99978
rect 244322 99922 244378 99978
rect 44518 94294 44574 94350
rect 44642 94294 44698 94350
rect 44518 94170 44574 94226
rect 44642 94170 44698 94226
rect 44518 94046 44574 94102
rect 44642 94046 44698 94102
rect 44518 93922 44574 93978
rect 44642 93922 44698 93978
rect 75238 94294 75294 94350
rect 75362 94294 75418 94350
rect 75238 94170 75294 94226
rect 75362 94170 75418 94226
rect 75238 94046 75294 94102
rect 75362 94046 75418 94102
rect 75238 93922 75294 93978
rect 75362 93922 75418 93978
rect 105958 94294 106014 94350
rect 106082 94294 106138 94350
rect 105958 94170 106014 94226
rect 106082 94170 106138 94226
rect 105958 94046 106014 94102
rect 106082 94046 106138 94102
rect 105958 93922 106014 93978
rect 106082 93922 106138 93978
rect 136678 94294 136734 94350
rect 136802 94294 136858 94350
rect 136678 94170 136734 94226
rect 136802 94170 136858 94226
rect 136678 94046 136734 94102
rect 136802 94046 136858 94102
rect 136678 93922 136734 93978
rect 136802 93922 136858 93978
rect 167398 94294 167454 94350
rect 167522 94294 167578 94350
rect 167398 94170 167454 94226
rect 167522 94170 167578 94226
rect 167398 94046 167454 94102
rect 167522 94046 167578 94102
rect 167398 93922 167454 93978
rect 167522 93922 167578 93978
rect 198118 94294 198174 94350
rect 198242 94294 198298 94350
rect 198118 94170 198174 94226
rect 198242 94170 198298 94226
rect 198118 94046 198174 94102
rect 198242 94046 198298 94102
rect 198118 93922 198174 93978
rect 198242 93922 198298 93978
rect 228838 94294 228894 94350
rect 228962 94294 229018 94350
rect 228838 94170 228894 94226
rect 228962 94170 229018 94226
rect 228838 94046 228894 94102
rect 228962 94046 229018 94102
rect 228838 93922 228894 93978
rect 228962 93922 229018 93978
rect 259558 94294 259614 94350
rect 259682 94294 259738 94350
rect 259558 94170 259614 94226
rect 259682 94170 259738 94226
rect 259558 94046 259614 94102
rect 259682 94046 259738 94102
rect 259558 93922 259614 93978
rect 259682 93922 259738 93978
rect 59878 82294 59934 82350
rect 60002 82294 60058 82350
rect 59878 82170 59934 82226
rect 60002 82170 60058 82226
rect 59878 82046 59934 82102
rect 60002 82046 60058 82102
rect 59878 81922 59934 81978
rect 60002 81922 60058 81978
rect 90598 82294 90654 82350
rect 90722 82294 90778 82350
rect 90598 82170 90654 82226
rect 90722 82170 90778 82226
rect 90598 82046 90654 82102
rect 90722 82046 90778 82102
rect 90598 81922 90654 81978
rect 90722 81922 90778 81978
rect 121318 82294 121374 82350
rect 121442 82294 121498 82350
rect 121318 82170 121374 82226
rect 121442 82170 121498 82226
rect 121318 82046 121374 82102
rect 121442 82046 121498 82102
rect 121318 81922 121374 81978
rect 121442 81922 121498 81978
rect 152038 82294 152094 82350
rect 152162 82294 152218 82350
rect 152038 82170 152094 82226
rect 152162 82170 152218 82226
rect 152038 82046 152094 82102
rect 152162 82046 152218 82102
rect 152038 81922 152094 81978
rect 152162 81922 152218 81978
rect 182758 82294 182814 82350
rect 182882 82294 182938 82350
rect 182758 82170 182814 82226
rect 182882 82170 182938 82226
rect 182758 82046 182814 82102
rect 182882 82046 182938 82102
rect 182758 81922 182814 81978
rect 182882 81922 182938 81978
rect 213478 82294 213534 82350
rect 213602 82294 213658 82350
rect 213478 82170 213534 82226
rect 213602 82170 213658 82226
rect 213478 82046 213534 82102
rect 213602 82046 213658 82102
rect 213478 81922 213534 81978
rect 213602 81922 213658 81978
rect 244198 82294 244254 82350
rect 244322 82294 244378 82350
rect 244198 82170 244254 82226
rect 244322 82170 244378 82226
rect 244198 82046 244254 82102
rect 244322 82046 244378 82102
rect 244198 81922 244254 81978
rect 244322 81922 244378 81978
rect 44518 76294 44574 76350
rect 44642 76294 44698 76350
rect 44518 76170 44574 76226
rect 44642 76170 44698 76226
rect 44518 76046 44574 76102
rect 44642 76046 44698 76102
rect 44518 75922 44574 75978
rect 44642 75922 44698 75978
rect 75238 76294 75294 76350
rect 75362 76294 75418 76350
rect 75238 76170 75294 76226
rect 75362 76170 75418 76226
rect 75238 76046 75294 76102
rect 75362 76046 75418 76102
rect 75238 75922 75294 75978
rect 75362 75922 75418 75978
rect 105958 76294 106014 76350
rect 106082 76294 106138 76350
rect 105958 76170 106014 76226
rect 106082 76170 106138 76226
rect 105958 76046 106014 76102
rect 106082 76046 106138 76102
rect 105958 75922 106014 75978
rect 106082 75922 106138 75978
rect 136678 76294 136734 76350
rect 136802 76294 136858 76350
rect 136678 76170 136734 76226
rect 136802 76170 136858 76226
rect 136678 76046 136734 76102
rect 136802 76046 136858 76102
rect 136678 75922 136734 75978
rect 136802 75922 136858 75978
rect 167398 76294 167454 76350
rect 167522 76294 167578 76350
rect 167398 76170 167454 76226
rect 167522 76170 167578 76226
rect 167398 76046 167454 76102
rect 167522 76046 167578 76102
rect 167398 75922 167454 75978
rect 167522 75922 167578 75978
rect 198118 76294 198174 76350
rect 198242 76294 198298 76350
rect 198118 76170 198174 76226
rect 198242 76170 198298 76226
rect 198118 76046 198174 76102
rect 198242 76046 198298 76102
rect 198118 75922 198174 75978
rect 198242 75922 198298 75978
rect 228838 76294 228894 76350
rect 228962 76294 229018 76350
rect 228838 76170 228894 76226
rect 228962 76170 229018 76226
rect 228838 76046 228894 76102
rect 228962 76046 229018 76102
rect 228838 75922 228894 75978
rect 228962 75922 229018 75978
rect 259558 76294 259614 76350
rect 259682 76294 259738 76350
rect 259558 76170 259614 76226
rect 259682 76170 259738 76226
rect 259558 76046 259614 76102
rect 259682 76046 259738 76102
rect 259558 75922 259614 75978
rect 259682 75922 259738 75978
rect 59878 64294 59934 64350
rect 60002 64294 60058 64350
rect 59878 64170 59934 64226
rect 60002 64170 60058 64226
rect 59878 64046 59934 64102
rect 60002 64046 60058 64102
rect 59878 63922 59934 63978
rect 60002 63922 60058 63978
rect 90598 64294 90654 64350
rect 90722 64294 90778 64350
rect 90598 64170 90654 64226
rect 90722 64170 90778 64226
rect 90598 64046 90654 64102
rect 90722 64046 90778 64102
rect 90598 63922 90654 63978
rect 90722 63922 90778 63978
rect 121318 64294 121374 64350
rect 121442 64294 121498 64350
rect 121318 64170 121374 64226
rect 121442 64170 121498 64226
rect 121318 64046 121374 64102
rect 121442 64046 121498 64102
rect 121318 63922 121374 63978
rect 121442 63922 121498 63978
rect 152038 64294 152094 64350
rect 152162 64294 152218 64350
rect 152038 64170 152094 64226
rect 152162 64170 152218 64226
rect 152038 64046 152094 64102
rect 152162 64046 152218 64102
rect 152038 63922 152094 63978
rect 152162 63922 152218 63978
rect 182758 64294 182814 64350
rect 182882 64294 182938 64350
rect 182758 64170 182814 64226
rect 182882 64170 182938 64226
rect 182758 64046 182814 64102
rect 182882 64046 182938 64102
rect 182758 63922 182814 63978
rect 182882 63922 182938 63978
rect 213478 64294 213534 64350
rect 213602 64294 213658 64350
rect 213478 64170 213534 64226
rect 213602 64170 213658 64226
rect 213478 64046 213534 64102
rect 213602 64046 213658 64102
rect 213478 63922 213534 63978
rect 213602 63922 213658 63978
rect 244198 64294 244254 64350
rect 244322 64294 244378 64350
rect 244198 64170 244254 64226
rect 244322 64170 244378 64226
rect 244198 64046 244254 64102
rect 244322 64046 244378 64102
rect 244198 63922 244254 63978
rect 244322 63922 244378 63978
rect 44518 58294 44574 58350
rect 44642 58294 44698 58350
rect 44518 58170 44574 58226
rect 44642 58170 44698 58226
rect 44518 58046 44574 58102
rect 44642 58046 44698 58102
rect 44518 57922 44574 57978
rect 44642 57922 44698 57978
rect 75238 58294 75294 58350
rect 75362 58294 75418 58350
rect 75238 58170 75294 58226
rect 75362 58170 75418 58226
rect 75238 58046 75294 58102
rect 75362 58046 75418 58102
rect 75238 57922 75294 57978
rect 75362 57922 75418 57978
rect 105958 58294 106014 58350
rect 106082 58294 106138 58350
rect 105958 58170 106014 58226
rect 106082 58170 106138 58226
rect 105958 58046 106014 58102
rect 106082 58046 106138 58102
rect 105958 57922 106014 57978
rect 106082 57922 106138 57978
rect 136678 58294 136734 58350
rect 136802 58294 136858 58350
rect 136678 58170 136734 58226
rect 136802 58170 136858 58226
rect 136678 58046 136734 58102
rect 136802 58046 136858 58102
rect 136678 57922 136734 57978
rect 136802 57922 136858 57978
rect 167398 58294 167454 58350
rect 167522 58294 167578 58350
rect 167398 58170 167454 58226
rect 167522 58170 167578 58226
rect 167398 58046 167454 58102
rect 167522 58046 167578 58102
rect 167398 57922 167454 57978
rect 167522 57922 167578 57978
rect 198118 58294 198174 58350
rect 198242 58294 198298 58350
rect 198118 58170 198174 58226
rect 198242 58170 198298 58226
rect 198118 58046 198174 58102
rect 198242 58046 198298 58102
rect 198118 57922 198174 57978
rect 198242 57922 198298 57978
rect 228838 58294 228894 58350
rect 228962 58294 229018 58350
rect 228838 58170 228894 58226
rect 228962 58170 229018 58226
rect 228838 58046 228894 58102
rect 228962 58046 229018 58102
rect 228838 57922 228894 57978
rect 228962 57922 229018 57978
rect 259558 58294 259614 58350
rect 259682 58294 259738 58350
rect 259558 58170 259614 58226
rect 259682 58170 259738 58226
rect 259558 58046 259614 58102
rect 259682 58046 259738 58102
rect 259558 57922 259614 57978
rect 259682 57922 259738 57978
rect 66954 40294 67010 40350
rect 67078 40294 67134 40350
rect 67202 40294 67258 40350
rect 67326 40294 67382 40350
rect 66954 40170 67010 40226
rect 67078 40170 67134 40226
rect 67202 40170 67258 40226
rect 67326 40170 67382 40226
rect 66954 40046 67010 40102
rect 67078 40046 67134 40102
rect 67202 40046 67258 40102
rect 67326 40046 67382 40102
rect 66954 39922 67010 39978
rect 67078 39922 67134 39978
rect 67202 39922 67258 39978
rect 67326 39922 67382 39978
rect 66954 22294 67010 22350
rect 67078 22294 67134 22350
rect 67202 22294 67258 22350
rect 67326 22294 67382 22350
rect 66954 22170 67010 22226
rect 67078 22170 67134 22226
rect 67202 22170 67258 22226
rect 67326 22170 67382 22226
rect 66954 22046 67010 22102
rect 67078 22046 67134 22102
rect 67202 22046 67258 22102
rect 67326 22046 67382 22102
rect 66954 21922 67010 21978
rect 67078 21922 67134 21978
rect 67202 21922 67258 21978
rect 67326 21922 67382 21978
rect 57148 4922 57204 4978
rect 55132 4742 55188 4798
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 70674 46294 70730 46350
rect 70798 46294 70854 46350
rect 70922 46294 70978 46350
rect 71046 46294 71102 46350
rect 70674 46170 70730 46226
rect 70798 46170 70854 46226
rect 70922 46170 70978 46226
rect 71046 46170 71102 46226
rect 70674 46046 70730 46102
rect 70798 46046 70854 46102
rect 70922 46046 70978 46102
rect 71046 46046 71102 46102
rect 70674 45922 70730 45978
rect 70798 45922 70854 45978
rect 70922 45922 70978 45978
rect 71046 45922 71102 45978
rect 90636 47762 90692 47818
rect 70674 28294 70730 28350
rect 70798 28294 70854 28350
rect 70922 28294 70978 28350
rect 71046 28294 71102 28350
rect 70674 28170 70730 28226
rect 70798 28170 70854 28226
rect 70922 28170 70978 28226
rect 71046 28170 71102 28226
rect 70674 28046 70730 28102
rect 70798 28046 70854 28102
rect 70922 28046 70978 28102
rect 71046 28046 71102 28102
rect 70674 27922 70730 27978
rect 70798 27922 70854 27978
rect 70922 27922 70978 27978
rect 71046 27922 71102 27978
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 75516 41102 75572 41158
rect 97674 40294 97730 40350
rect 97798 40294 97854 40350
rect 97922 40294 97978 40350
rect 98046 40294 98102 40350
rect 97674 40170 97730 40226
rect 97798 40170 97854 40226
rect 97922 40170 97978 40226
rect 98046 40170 98102 40226
rect 97674 40046 97730 40102
rect 97798 40046 97854 40102
rect 97922 40046 97978 40102
rect 98046 40046 98102 40102
rect 97674 39922 97730 39978
rect 97798 39922 97854 39978
rect 97922 39922 97978 39978
rect 98046 39922 98102 39978
rect 97674 22294 97730 22350
rect 97798 22294 97854 22350
rect 97922 22294 97978 22350
rect 98046 22294 98102 22350
rect 97674 22170 97730 22226
rect 97798 22170 97854 22226
rect 97922 22170 97978 22226
rect 98046 22170 98102 22226
rect 97674 22046 97730 22102
rect 97798 22046 97854 22102
rect 97922 22046 97978 22102
rect 98046 22046 98102 22102
rect 97674 21922 97730 21978
rect 97798 21922 97854 21978
rect 97922 21922 97978 21978
rect 98046 21922 98102 21978
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 101394 46294 101450 46350
rect 101518 46294 101574 46350
rect 101642 46294 101698 46350
rect 101766 46294 101822 46350
rect 101394 46170 101450 46226
rect 101518 46170 101574 46226
rect 101642 46170 101698 46226
rect 101766 46170 101822 46226
rect 101394 46046 101450 46102
rect 101518 46046 101574 46102
rect 101642 46046 101698 46102
rect 101766 46046 101822 46102
rect 101394 45922 101450 45978
rect 101518 45922 101574 45978
rect 101642 45922 101698 45978
rect 101766 45922 101822 45978
rect 110796 47942 110852 47998
rect 101394 28294 101450 28350
rect 101518 28294 101574 28350
rect 101642 28294 101698 28350
rect 101766 28294 101822 28350
rect 101394 28170 101450 28226
rect 101518 28170 101574 28226
rect 101642 28170 101698 28226
rect 101766 28170 101822 28226
rect 101394 28046 101450 28102
rect 101518 28046 101574 28102
rect 101642 28046 101698 28102
rect 101766 28046 101822 28102
rect 101394 27922 101450 27978
rect 101518 27922 101574 27978
rect 101642 27922 101698 27978
rect 101766 27922 101822 27978
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 104076 44522 104132 44578
rect 128394 40294 128450 40350
rect 128518 40294 128574 40350
rect 128642 40294 128698 40350
rect 128766 40294 128822 40350
rect 128394 40170 128450 40226
rect 128518 40170 128574 40226
rect 128642 40170 128698 40226
rect 128766 40170 128822 40226
rect 128394 40046 128450 40102
rect 128518 40046 128574 40102
rect 128642 40046 128698 40102
rect 128766 40046 128822 40102
rect 128394 39922 128450 39978
rect 128518 39922 128574 39978
rect 128642 39922 128698 39978
rect 128766 39922 128822 39978
rect 128394 22294 128450 22350
rect 128518 22294 128574 22350
rect 128642 22294 128698 22350
rect 128766 22294 128822 22350
rect 128394 22170 128450 22226
rect 128518 22170 128574 22226
rect 128642 22170 128698 22226
rect 128766 22170 128822 22226
rect 128394 22046 128450 22102
rect 128518 22046 128574 22102
rect 128642 22046 128698 22102
rect 128766 22046 128822 22102
rect 128394 21922 128450 21978
rect 128518 21922 128574 21978
rect 128642 21922 128698 21978
rect 128766 21922 128822 21978
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 132114 46294 132170 46350
rect 132238 46294 132294 46350
rect 132362 46294 132418 46350
rect 132486 46294 132542 46350
rect 132114 46170 132170 46226
rect 132238 46170 132294 46226
rect 132362 46170 132418 46226
rect 132486 46170 132542 46226
rect 132114 46046 132170 46102
rect 132238 46046 132294 46102
rect 132362 46046 132418 46102
rect 132486 46046 132542 46102
rect 132114 45922 132170 45978
rect 132238 45922 132294 45978
rect 132362 45922 132418 45978
rect 132486 45922 132542 45978
rect 132114 28294 132170 28350
rect 132238 28294 132294 28350
rect 132362 28294 132418 28350
rect 132486 28294 132542 28350
rect 132114 28170 132170 28226
rect 132238 28170 132294 28226
rect 132362 28170 132418 28226
rect 132486 28170 132542 28226
rect 132114 28046 132170 28102
rect 132238 28046 132294 28102
rect 132362 28046 132418 28102
rect 132486 28046 132542 28102
rect 132114 27922 132170 27978
rect 132238 27922 132294 27978
rect 132362 27922 132418 27978
rect 132486 27922 132542 27978
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 154476 44702 154532 44758
rect 137228 4922 137284 4978
rect 148652 4742 148708 4798
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 189834 40294 189890 40350
rect 189958 40294 190014 40350
rect 190082 40294 190138 40350
rect 190206 40294 190262 40350
rect 189834 40170 189890 40226
rect 189958 40170 190014 40226
rect 190082 40170 190138 40226
rect 190206 40170 190262 40226
rect 189834 40046 189890 40102
rect 189958 40046 190014 40102
rect 190082 40046 190138 40102
rect 190206 40046 190262 40102
rect 189834 39922 189890 39978
rect 189958 39922 190014 39978
rect 190082 39922 190138 39978
rect 190206 39922 190262 39978
rect 189834 22294 189890 22350
rect 189958 22294 190014 22350
rect 190082 22294 190138 22350
rect 190206 22294 190262 22350
rect 189834 22170 189890 22226
rect 189958 22170 190014 22226
rect 190082 22170 190138 22226
rect 190206 22170 190262 22226
rect 189834 22046 189890 22102
rect 189958 22046 190014 22102
rect 190082 22046 190138 22102
rect 190206 22046 190262 22102
rect 189834 21922 189890 21978
rect 189958 21922 190014 21978
rect 190082 21922 190138 21978
rect 190206 21922 190262 21978
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 193554 46294 193610 46350
rect 193678 46294 193734 46350
rect 193802 46294 193858 46350
rect 193926 46294 193982 46350
rect 193554 46170 193610 46226
rect 193678 46170 193734 46226
rect 193802 46170 193858 46226
rect 193926 46170 193982 46226
rect 193554 46046 193610 46102
rect 193678 46046 193734 46102
rect 193802 46046 193858 46102
rect 193926 46046 193982 46102
rect 193554 45922 193610 45978
rect 193678 45922 193734 45978
rect 193802 45922 193858 45978
rect 193926 45922 193982 45978
rect 193554 28294 193610 28350
rect 193678 28294 193734 28350
rect 193802 28294 193858 28350
rect 193926 28294 193982 28350
rect 193554 28170 193610 28226
rect 193678 28170 193734 28226
rect 193802 28170 193858 28226
rect 193926 28170 193982 28226
rect 193554 28046 193610 28102
rect 193678 28046 193734 28102
rect 193802 28046 193858 28102
rect 193926 28046 193982 28102
rect 193554 27922 193610 27978
rect 193678 27922 193734 27978
rect 193802 27922 193858 27978
rect 193926 27922 193982 27978
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 220554 40294 220610 40350
rect 220678 40294 220734 40350
rect 220802 40294 220858 40350
rect 220926 40294 220982 40350
rect 220554 40170 220610 40226
rect 220678 40170 220734 40226
rect 220802 40170 220858 40226
rect 220926 40170 220982 40226
rect 220554 40046 220610 40102
rect 220678 40046 220734 40102
rect 220802 40046 220858 40102
rect 220926 40046 220982 40102
rect 220554 39922 220610 39978
rect 220678 39922 220734 39978
rect 220802 39922 220858 39978
rect 220926 39922 220982 39978
rect 220554 22294 220610 22350
rect 220678 22294 220734 22350
rect 220802 22294 220858 22350
rect 220926 22294 220982 22350
rect 220554 22170 220610 22226
rect 220678 22170 220734 22226
rect 220802 22170 220858 22226
rect 220926 22170 220982 22226
rect 220554 22046 220610 22102
rect 220678 22046 220734 22102
rect 220802 22046 220858 22102
rect 220926 22046 220982 22102
rect 220554 21922 220610 21978
rect 220678 21922 220734 21978
rect 220802 21922 220858 21978
rect 220926 21922 220982 21978
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 224274 46294 224330 46350
rect 224398 46294 224454 46350
rect 224522 46294 224578 46350
rect 224646 46294 224702 46350
rect 224274 46170 224330 46226
rect 224398 46170 224454 46226
rect 224522 46170 224578 46226
rect 224646 46170 224702 46226
rect 224274 46046 224330 46102
rect 224398 46046 224454 46102
rect 224522 46046 224578 46102
rect 224646 46046 224702 46102
rect 224274 45922 224330 45978
rect 224398 45922 224454 45978
rect 224522 45922 224578 45978
rect 224646 45922 224702 45978
rect 224274 28294 224330 28350
rect 224398 28294 224454 28350
rect 224522 28294 224578 28350
rect 224646 28294 224702 28350
rect 224274 28170 224330 28226
rect 224398 28170 224454 28226
rect 224522 28170 224578 28226
rect 224646 28170 224702 28226
rect 224274 28046 224330 28102
rect 224398 28046 224454 28102
rect 224522 28046 224578 28102
rect 224646 28046 224702 28102
rect 224274 27922 224330 27978
rect 224398 27922 224454 27978
rect 224522 27922 224578 27978
rect 224646 27922 224702 27978
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 251274 40294 251330 40350
rect 251398 40294 251454 40350
rect 251522 40294 251578 40350
rect 251646 40294 251702 40350
rect 251274 40170 251330 40226
rect 251398 40170 251454 40226
rect 251522 40170 251578 40226
rect 251646 40170 251702 40226
rect 251274 40046 251330 40102
rect 251398 40046 251454 40102
rect 251522 40046 251578 40102
rect 251646 40046 251702 40102
rect 251274 39922 251330 39978
rect 251398 39922 251454 39978
rect 251522 39922 251578 39978
rect 251646 39922 251702 39978
rect 251274 22294 251330 22350
rect 251398 22294 251454 22350
rect 251522 22294 251578 22350
rect 251646 22294 251702 22350
rect 251274 22170 251330 22226
rect 251398 22170 251454 22226
rect 251522 22170 251578 22226
rect 251646 22170 251702 22226
rect 251274 22046 251330 22102
rect 251398 22046 251454 22102
rect 251522 22046 251578 22102
rect 251646 22046 251702 22102
rect 251274 21922 251330 21978
rect 251398 21922 251454 21978
rect 251522 21922 251578 21978
rect 251646 21922 251702 21978
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 267036 209042 267092 209098
rect 267148 231002 267204 231058
rect 254994 46294 255050 46350
rect 255118 46294 255174 46350
rect 255242 46294 255298 46350
rect 255366 46294 255422 46350
rect 254994 46170 255050 46226
rect 255118 46170 255174 46226
rect 255242 46170 255298 46226
rect 255366 46170 255422 46226
rect 254994 46046 255050 46102
rect 255118 46046 255174 46102
rect 255242 46046 255298 46102
rect 255366 46046 255422 46102
rect 254994 45922 255050 45978
rect 255118 45922 255174 45978
rect 255242 45922 255298 45978
rect 255366 45922 255422 45978
rect 254994 28294 255050 28350
rect 255118 28294 255174 28350
rect 255242 28294 255298 28350
rect 255366 28294 255422 28350
rect 254994 28170 255050 28226
rect 255118 28170 255174 28226
rect 255242 28170 255298 28226
rect 255366 28170 255422 28226
rect 254994 28046 255050 28102
rect 255118 28046 255174 28102
rect 255242 28046 255298 28102
rect 255366 28046 255422 28102
rect 254994 27922 255050 27978
rect 255118 27922 255174 27978
rect 255242 27922 255298 27978
rect 255366 27922 255422 27978
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 267372 224522 267428 224578
rect 267484 47942 267540 47998
rect 267596 211382 267652 211438
rect 268604 110042 268660 110098
rect 269164 211202 269220 211258
rect 268716 106622 268772 106678
rect 269724 231182 269780 231238
rect 269948 231362 270004 231418
rect 270060 47762 270116 47818
rect 270732 227942 270788 227998
rect 270844 227762 270900 227818
rect 270956 227582 271012 227638
rect 273868 224162 273924 224218
rect 272300 153636 272356 153658
rect 272300 153602 272356 153636
rect 277228 236942 277284 236998
rect 275548 224342 275604 224398
rect 274092 210122 274148 210178
rect 274204 208682 274260 208738
rect 274652 153422 274708 153478
rect 281372 4742 281428 4798
rect 281994 238294 282050 238350
rect 282118 238294 282174 238350
rect 282242 238294 282298 238350
rect 282366 238294 282422 238350
rect 281994 238170 282050 238226
rect 282118 238170 282174 238226
rect 282242 238170 282298 238226
rect 282366 238170 282422 238226
rect 281994 238046 282050 238102
rect 282118 238046 282174 238102
rect 282242 238046 282298 238102
rect 282366 238046 282422 238102
rect 281994 237922 282050 237978
rect 282118 237922 282174 237978
rect 282242 237922 282298 237978
rect 282366 237922 282422 237978
rect 281994 220294 282050 220350
rect 282118 220294 282174 220350
rect 282242 220294 282298 220350
rect 282366 220294 282422 220350
rect 281994 220170 282050 220226
rect 282118 220170 282174 220226
rect 282242 220170 282298 220226
rect 282366 220170 282422 220226
rect 281994 220046 282050 220102
rect 282118 220046 282174 220102
rect 282242 220046 282298 220102
rect 282366 220046 282422 220102
rect 281994 219922 282050 219978
rect 282118 219922 282174 219978
rect 282242 219922 282298 219978
rect 282366 219922 282422 219978
rect 281994 202294 282050 202350
rect 282118 202294 282174 202350
rect 282242 202294 282298 202350
rect 282366 202294 282422 202350
rect 281994 202170 282050 202226
rect 282118 202170 282174 202226
rect 282242 202170 282298 202226
rect 282366 202170 282422 202226
rect 281994 202046 282050 202102
rect 282118 202046 282174 202102
rect 282242 202046 282298 202102
rect 282366 202046 282422 202102
rect 281994 201922 282050 201978
rect 282118 201922 282174 201978
rect 282242 201922 282298 201978
rect 282366 201922 282422 201978
rect 281994 184294 282050 184350
rect 282118 184294 282174 184350
rect 282242 184294 282298 184350
rect 282366 184294 282422 184350
rect 281994 184170 282050 184226
rect 282118 184170 282174 184226
rect 282242 184170 282298 184226
rect 282366 184170 282422 184226
rect 281994 184046 282050 184102
rect 282118 184046 282174 184102
rect 282242 184046 282298 184102
rect 282366 184046 282422 184102
rect 281994 183922 282050 183978
rect 282118 183922 282174 183978
rect 282242 183922 282298 183978
rect 282366 183922 282422 183978
rect 281994 166294 282050 166350
rect 282118 166294 282174 166350
rect 282242 166294 282298 166350
rect 282366 166294 282422 166350
rect 281994 166170 282050 166226
rect 282118 166170 282174 166226
rect 282242 166170 282298 166226
rect 282366 166170 282422 166226
rect 281994 166046 282050 166102
rect 282118 166046 282174 166102
rect 282242 166046 282298 166102
rect 282366 166046 282422 166102
rect 281994 165922 282050 165978
rect 282118 165922 282174 165978
rect 282242 165922 282298 165978
rect 282366 165922 282422 165978
rect 281994 148294 282050 148350
rect 282118 148294 282174 148350
rect 282242 148294 282298 148350
rect 282366 148294 282422 148350
rect 281994 148170 282050 148226
rect 282118 148170 282174 148226
rect 282242 148170 282298 148226
rect 282366 148170 282422 148226
rect 281994 148046 282050 148102
rect 282118 148046 282174 148102
rect 282242 148046 282298 148102
rect 282366 148046 282422 148102
rect 281994 147922 282050 147978
rect 282118 147922 282174 147978
rect 282242 147922 282298 147978
rect 282366 147922 282422 147978
rect 281994 130294 282050 130350
rect 282118 130294 282174 130350
rect 282242 130294 282298 130350
rect 282366 130294 282422 130350
rect 281994 130170 282050 130226
rect 282118 130170 282174 130226
rect 282242 130170 282298 130226
rect 282366 130170 282422 130226
rect 281994 130046 282050 130102
rect 282118 130046 282174 130102
rect 282242 130046 282298 130102
rect 282366 130046 282422 130102
rect 281994 129922 282050 129978
rect 282118 129922 282174 129978
rect 282242 129922 282298 129978
rect 282366 129922 282422 129978
rect 281994 112294 282050 112350
rect 282118 112294 282174 112350
rect 282242 112294 282298 112350
rect 282366 112294 282422 112350
rect 281994 112170 282050 112226
rect 282118 112170 282174 112226
rect 282242 112170 282298 112226
rect 282366 112170 282422 112226
rect 281994 112046 282050 112102
rect 282118 112046 282174 112102
rect 282242 112046 282298 112102
rect 282366 112046 282422 112102
rect 281994 111922 282050 111978
rect 282118 111922 282174 111978
rect 282242 111922 282298 111978
rect 282366 111922 282422 111978
rect 281994 94294 282050 94350
rect 282118 94294 282174 94350
rect 282242 94294 282298 94350
rect 282366 94294 282422 94350
rect 281994 94170 282050 94226
rect 282118 94170 282174 94226
rect 282242 94170 282298 94226
rect 282366 94170 282422 94226
rect 281994 94046 282050 94102
rect 282118 94046 282174 94102
rect 282242 94046 282298 94102
rect 282366 94046 282422 94102
rect 281994 93922 282050 93978
rect 282118 93922 282174 93978
rect 282242 93922 282298 93978
rect 282366 93922 282422 93978
rect 281994 76294 282050 76350
rect 282118 76294 282174 76350
rect 282242 76294 282298 76350
rect 282366 76294 282422 76350
rect 281994 76170 282050 76226
rect 282118 76170 282174 76226
rect 282242 76170 282298 76226
rect 282366 76170 282422 76226
rect 281994 76046 282050 76102
rect 282118 76046 282174 76102
rect 282242 76046 282298 76102
rect 282366 76046 282422 76102
rect 281994 75922 282050 75978
rect 282118 75922 282174 75978
rect 282242 75922 282298 75978
rect 282366 75922 282422 75978
rect 281994 58294 282050 58350
rect 282118 58294 282174 58350
rect 282242 58294 282298 58350
rect 282366 58294 282422 58350
rect 281994 58170 282050 58226
rect 282118 58170 282174 58226
rect 282242 58170 282298 58226
rect 282366 58170 282422 58226
rect 281994 58046 282050 58102
rect 282118 58046 282174 58102
rect 282242 58046 282298 58102
rect 282366 58046 282422 58102
rect 281994 57922 282050 57978
rect 282118 57922 282174 57978
rect 282242 57922 282298 57978
rect 282366 57922 282422 57978
rect 283052 44702 283108 44758
rect 285714 226294 285770 226350
rect 285838 226294 285894 226350
rect 285962 226294 286018 226350
rect 286086 226294 286142 226350
rect 285714 226170 285770 226226
rect 285838 226170 285894 226226
rect 285962 226170 286018 226226
rect 286086 226170 286142 226226
rect 285714 226046 285770 226102
rect 285838 226046 285894 226102
rect 285962 226046 286018 226102
rect 286086 226046 286142 226102
rect 285714 225922 285770 225978
rect 285838 225922 285894 225978
rect 285962 225922 286018 225978
rect 286086 225922 286142 225978
rect 285714 208294 285770 208350
rect 285838 208294 285894 208350
rect 285962 208294 286018 208350
rect 286086 208294 286142 208350
rect 285714 208170 285770 208226
rect 285838 208170 285894 208226
rect 285962 208170 286018 208226
rect 286086 208170 286142 208226
rect 285714 208046 285770 208102
rect 285838 208046 285894 208102
rect 285962 208046 286018 208102
rect 286086 208046 286142 208102
rect 285714 207922 285770 207978
rect 285838 207922 285894 207978
rect 285962 207922 286018 207978
rect 286086 207922 286142 207978
rect 285714 190294 285770 190350
rect 285838 190294 285894 190350
rect 285962 190294 286018 190350
rect 286086 190294 286142 190350
rect 285714 190170 285770 190226
rect 285838 190170 285894 190226
rect 285962 190170 286018 190226
rect 286086 190170 286142 190226
rect 285714 190046 285770 190102
rect 285838 190046 285894 190102
rect 285962 190046 286018 190102
rect 286086 190046 286142 190102
rect 285714 189922 285770 189978
rect 285838 189922 285894 189978
rect 285962 189922 286018 189978
rect 286086 189922 286142 189978
rect 285714 172294 285770 172350
rect 285838 172294 285894 172350
rect 285962 172294 286018 172350
rect 286086 172294 286142 172350
rect 285714 172170 285770 172226
rect 285838 172170 285894 172226
rect 285962 172170 286018 172226
rect 286086 172170 286142 172226
rect 285714 172046 285770 172102
rect 285838 172046 285894 172102
rect 285962 172046 286018 172102
rect 286086 172046 286142 172102
rect 285714 171922 285770 171978
rect 285838 171922 285894 171978
rect 285962 171922 286018 171978
rect 286086 171922 286142 171978
rect 285714 154294 285770 154350
rect 285838 154294 285894 154350
rect 285962 154294 286018 154350
rect 286086 154294 286142 154350
rect 285714 154170 285770 154226
rect 285838 154170 285894 154226
rect 285962 154170 286018 154226
rect 286086 154170 286142 154226
rect 285714 154046 285770 154102
rect 285838 154046 285894 154102
rect 285962 154046 286018 154102
rect 286086 154046 286142 154102
rect 285714 153922 285770 153978
rect 285838 153922 285894 153978
rect 285962 153922 286018 153978
rect 286086 153922 286142 153978
rect 285714 136294 285770 136350
rect 285838 136294 285894 136350
rect 285962 136294 286018 136350
rect 286086 136294 286142 136350
rect 285714 136170 285770 136226
rect 285838 136170 285894 136226
rect 285962 136170 286018 136226
rect 286086 136170 286142 136226
rect 285714 136046 285770 136102
rect 285838 136046 285894 136102
rect 285962 136046 286018 136102
rect 286086 136046 286142 136102
rect 285714 135922 285770 135978
rect 285838 135922 285894 135978
rect 285962 135922 286018 135978
rect 286086 135922 286142 135978
rect 285714 118294 285770 118350
rect 285838 118294 285894 118350
rect 285962 118294 286018 118350
rect 286086 118294 286142 118350
rect 285714 118170 285770 118226
rect 285838 118170 285894 118226
rect 285962 118170 286018 118226
rect 286086 118170 286142 118226
rect 285714 118046 285770 118102
rect 285838 118046 285894 118102
rect 285962 118046 286018 118102
rect 286086 118046 286142 118102
rect 285714 117922 285770 117978
rect 285838 117922 285894 117978
rect 285962 117922 286018 117978
rect 286086 117922 286142 117978
rect 285714 100294 285770 100350
rect 285838 100294 285894 100350
rect 285962 100294 286018 100350
rect 286086 100294 286142 100350
rect 285714 100170 285770 100226
rect 285838 100170 285894 100226
rect 285962 100170 286018 100226
rect 286086 100170 286142 100226
rect 285714 100046 285770 100102
rect 285838 100046 285894 100102
rect 285962 100046 286018 100102
rect 286086 100046 286142 100102
rect 285714 99922 285770 99978
rect 285838 99922 285894 99978
rect 285962 99922 286018 99978
rect 286086 99922 286142 99978
rect 285714 82294 285770 82350
rect 285838 82294 285894 82350
rect 285962 82294 286018 82350
rect 286086 82294 286142 82350
rect 285714 82170 285770 82226
rect 285838 82170 285894 82226
rect 285962 82170 286018 82226
rect 286086 82170 286142 82226
rect 285714 82046 285770 82102
rect 285838 82046 285894 82102
rect 285962 82046 286018 82102
rect 286086 82046 286142 82102
rect 285714 81922 285770 81978
rect 285838 81922 285894 81978
rect 285962 81922 286018 81978
rect 286086 81922 286142 81978
rect 285714 64294 285770 64350
rect 285838 64294 285894 64350
rect 285962 64294 286018 64350
rect 286086 64294 286142 64350
rect 285714 64170 285770 64226
rect 285838 64170 285894 64226
rect 285962 64170 286018 64226
rect 286086 64170 286142 64226
rect 285714 64046 285770 64102
rect 285838 64046 285894 64102
rect 285962 64046 286018 64102
rect 286086 64046 286142 64102
rect 285714 63922 285770 63978
rect 285838 63922 285894 63978
rect 285962 63922 286018 63978
rect 286086 63922 286142 63978
rect 285714 46294 285770 46350
rect 285838 46294 285894 46350
rect 285962 46294 286018 46350
rect 286086 46294 286142 46350
rect 285714 46170 285770 46226
rect 285838 46170 285894 46226
rect 285962 46170 286018 46226
rect 286086 46170 286142 46226
rect 285714 46046 285770 46102
rect 285838 46046 285894 46102
rect 285962 46046 286018 46102
rect 286086 46046 286142 46102
rect 285714 45922 285770 45978
rect 285838 45922 285894 45978
rect 285962 45922 286018 45978
rect 286086 45922 286142 45978
rect 281994 40294 282050 40350
rect 282118 40294 282174 40350
rect 282242 40294 282298 40350
rect 282366 40294 282422 40350
rect 281994 40170 282050 40226
rect 282118 40170 282174 40226
rect 282242 40170 282298 40226
rect 282366 40170 282422 40226
rect 281994 40046 282050 40102
rect 282118 40046 282174 40102
rect 282242 40046 282298 40102
rect 282366 40046 282422 40102
rect 281994 39922 282050 39978
rect 282118 39922 282174 39978
rect 282242 39922 282298 39978
rect 282366 39922 282422 39978
rect 281994 22294 282050 22350
rect 282118 22294 282174 22350
rect 282242 22294 282298 22350
rect 282366 22294 282422 22350
rect 281994 22170 282050 22226
rect 282118 22170 282174 22226
rect 282242 22170 282298 22226
rect 282366 22170 282422 22226
rect 281994 22046 282050 22102
rect 282118 22046 282174 22102
rect 282242 22046 282298 22102
rect 282366 22046 282422 22102
rect 281994 21922 282050 21978
rect 282118 21922 282174 21978
rect 282242 21922 282298 21978
rect 282366 21922 282422 21978
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 285714 28294 285770 28350
rect 285838 28294 285894 28350
rect 285962 28294 286018 28350
rect 286086 28294 286142 28350
rect 285714 28170 285770 28226
rect 285838 28170 285894 28226
rect 285962 28170 286018 28226
rect 286086 28170 286142 28226
rect 285714 28046 285770 28102
rect 285838 28046 285894 28102
rect 285962 28046 286018 28102
rect 286086 28046 286142 28102
rect 285714 27922 285770 27978
rect 285838 27922 285894 27978
rect 285962 27922 286018 27978
rect 286086 27922 286142 27978
rect 285714 10294 285770 10350
rect 285838 10294 285894 10350
rect 285962 10294 286018 10350
rect 286086 10294 286142 10350
rect 285714 10170 285770 10226
rect 285838 10170 285894 10226
rect 285962 10170 286018 10226
rect 286086 10170 286142 10226
rect 285714 10046 285770 10102
rect 285838 10046 285894 10102
rect 285962 10046 286018 10102
rect 286086 10046 286142 10102
rect 285714 9922 285770 9978
rect 285838 9922 285894 9978
rect 285962 9922 286018 9978
rect 286086 9922 286142 9978
rect 288316 4922 288372 4978
rect 312714 238294 312770 238350
rect 312838 238294 312894 238350
rect 312962 238294 313018 238350
rect 313086 238294 313142 238350
rect 312714 238170 312770 238226
rect 312838 238170 312894 238226
rect 312962 238170 313018 238226
rect 313086 238170 313142 238226
rect 312714 238046 312770 238102
rect 312838 238046 312894 238102
rect 312962 238046 313018 238102
rect 313086 238046 313142 238102
rect 312714 237922 312770 237978
rect 312838 237922 312894 237978
rect 312962 237922 313018 237978
rect 313086 237922 313142 237978
rect 293244 141902 293300 141958
rect 293132 104102 293188 104158
rect 296604 152702 296660 152758
rect 298172 209042 298228 209098
rect 298956 157382 299012 157438
rect 296492 103922 296548 103978
rect 305538 184294 305594 184350
rect 305662 184294 305718 184350
rect 305538 184170 305594 184226
rect 305662 184170 305718 184226
rect 305538 184046 305594 184102
rect 305662 184046 305718 184102
rect 305538 183922 305594 183978
rect 305662 183922 305718 183978
rect 305538 166294 305594 166350
rect 305662 166294 305718 166350
rect 305538 166170 305594 166226
rect 305662 166170 305718 166226
rect 305538 166046 305594 166102
rect 305662 166046 305718 166102
rect 305538 165922 305594 165978
rect 305662 165922 305718 165978
rect 309036 197522 309092 197578
rect 310716 197342 310772 197398
rect 312714 220294 312770 220350
rect 312838 220294 312894 220350
rect 312962 220294 313018 220350
rect 313086 220294 313142 220350
rect 312714 220170 312770 220226
rect 312838 220170 312894 220226
rect 312962 220170 313018 220226
rect 313086 220170 313142 220226
rect 312714 220046 312770 220102
rect 312838 220046 312894 220102
rect 312962 220046 313018 220102
rect 313086 220046 313142 220102
rect 312714 219922 312770 219978
rect 312838 219922 312894 219978
rect 312962 219922 313018 219978
rect 313086 219922 313142 219978
rect 312714 202294 312770 202350
rect 312838 202294 312894 202350
rect 312962 202294 313018 202350
rect 313086 202294 313142 202350
rect 312714 202170 312770 202226
rect 312838 202170 312894 202226
rect 312962 202170 313018 202226
rect 313086 202170 313142 202226
rect 312714 202046 312770 202102
rect 312838 202046 312894 202102
rect 312962 202046 313018 202102
rect 313086 202046 313142 202102
rect 312714 201922 312770 201978
rect 312838 201922 312894 201978
rect 312962 201922 313018 201978
rect 313086 201922 313142 201978
rect 336812 238562 336868 238618
rect 316434 226294 316490 226350
rect 316558 226294 316614 226350
rect 316682 226294 316738 226350
rect 316806 226294 316862 226350
rect 316434 226170 316490 226226
rect 316558 226170 316614 226226
rect 316682 226170 316738 226226
rect 316806 226170 316862 226226
rect 316434 226046 316490 226102
rect 316558 226046 316614 226102
rect 316682 226046 316738 226102
rect 316806 226046 316862 226102
rect 316434 225922 316490 225978
rect 316558 225922 316614 225978
rect 316682 225922 316738 225978
rect 316806 225922 316862 225978
rect 316434 208294 316490 208350
rect 316558 208294 316614 208350
rect 316682 208294 316738 208350
rect 316806 208294 316862 208350
rect 316434 208170 316490 208226
rect 316558 208170 316614 208226
rect 316682 208170 316738 208226
rect 316806 208170 316862 208226
rect 316434 208046 316490 208102
rect 316558 208046 316614 208102
rect 316682 208046 316738 208102
rect 316806 208046 316862 208102
rect 316434 207922 316490 207978
rect 316558 207922 316614 207978
rect 316682 207922 316738 207978
rect 316806 207922 316862 207978
rect 319116 193922 319172 193978
rect 334236 192302 334292 192358
rect 309822 190294 309878 190350
rect 309946 190294 310002 190350
rect 309822 190170 309878 190226
rect 309946 190170 310002 190226
rect 309822 190046 309878 190102
rect 309946 190046 310002 190102
rect 309822 189922 309878 189978
rect 309946 189922 310002 189978
rect 318390 190294 318446 190350
rect 318514 190294 318570 190350
rect 318390 190170 318446 190226
rect 318514 190170 318570 190226
rect 318390 190046 318446 190102
rect 318514 190046 318570 190102
rect 318390 189922 318446 189978
rect 318514 189922 318570 189978
rect 326958 190294 327014 190350
rect 327082 190294 327138 190350
rect 326958 190170 327014 190226
rect 327082 190170 327138 190226
rect 326958 190046 327014 190102
rect 327082 190046 327138 190102
rect 326958 189922 327014 189978
rect 327082 189922 327138 189978
rect 335526 190294 335582 190350
rect 335650 190294 335706 190350
rect 335526 190170 335582 190226
rect 335650 190170 335706 190226
rect 335526 190046 335582 190102
rect 335650 190046 335706 190102
rect 335526 189922 335582 189978
rect 335650 189922 335706 189978
rect 314106 184294 314162 184350
rect 314230 184294 314286 184350
rect 314106 184170 314162 184226
rect 314230 184170 314286 184226
rect 314106 184046 314162 184102
rect 314230 184046 314286 184102
rect 314106 183922 314162 183978
rect 314230 183922 314286 183978
rect 322674 184294 322730 184350
rect 322798 184294 322854 184350
rect 322674 184170 322730 184226
rect 322798 184170 322854 184226
rect 322674 184046 322730 184102
rect 322798 184046 322854 184102
rect 322674 183922 322730 183978
rect 322798 183922 322854 183978
rect 331242 184294 331298 184350
rect 331366 184294 331422 184350
rect 331242 184170 331298 184226
rect 331366 184170 331422 184226
rect 331242 184046 331298 184102
rect 331366 184046 331422 184102
rect 331242 183922 331298 183978
rect 331366 183922 331422 183978
rect 309822 172294 309878 172350
rect 309946 172294 310002 172350
rect 309822 172170 309878 172226
rect 309946 172170 310002 172226
rect 309822 172046 309878 172102
rect 309946 172046 310002 172102
rect 309822 171922 309878 171978
rect 309946 171922 310002 171978
rect 318390 172294 318446 172350
rect 318514 172294 318570 172350
rect 318390 172170 318446 172226
rect 318514 172170 318570 172226
rect 318390 172046 318446 172102
rect 318514 172046 318570 172102
rect 318390 171922 318446 171978
rect 318514 171922 318570 171978
rect 326958 172294 327014 172350
rect 327082 172294 327138 172350
rect 326958 172170 327014 172226
rect 327082 172170 327138 172226
rect 326958 172046 327014 172102
rect 327082 172046 327138 172102
rect 326958 171922 327014 171978
rect 327082 171922 327138 171978
rect 335526 172294 335582 172350
rect 335650 172294 335706 172350
rect 335526 172170 335582 172226
rect 335650 172170 335706 172226
rect 335526 172046 335582 172102
rect 335650 172046 335706 172102
rect 335526 171922 335582 171978
rect 335650 171922 335706 171978
rect 314106 166294 314162 166350
rect 314230 166294 314286 166350
rect 314106 166170 314162 166226
rect 314230 166170 314286 166226
rect 314106 166046 314162 166102
rect 314230 166046 314286 166102
rect 314106 165922 314162 165978
rect 314230 165922 314286 165978
rect 322674 166294 322730 166350
rect 322798 166294 322854 166350
rect 322674 166170 322730 166226
rect 322798 166170 322854 166226
rect 322674 166046 322730 166102
rect 322798 166046 322854 166102
rect 322674 165922 322730 165978
rect 322798 165922 322854 165978
rect 331242 166294 331298 166350
rect 331366 166294 331422 166350
rect 331242 166170 331298 166226
rect 331366 166170 331422 166226
rect 331242 166046 331298 166102
rect 331366 166046 331422 166102
rect 331242 165922 331298 165978
rect 331366 165922 331422 165978
rect 306572 157382 306628 157438
rect 312714 148294 312770 148350
rect 312838 148294 312894 148350
rect 312962 148294 313018 148350
rect 313086 148294 313142 148350
rect 312714 148170 312770 148226
rect 312838 148170 312894 148226
rect 312962 148170 313018 148226
rect 313086 148170 313142 148226
rect 312714 148046 312770 148102
rect 312838 148046 312894 148102
rect 312962 148046 313018 148102
rect 313086 148046 313142 148102
rect 312714 147922 312770 147978
rect 312838 147922 312894 147978
rect 312962 147922 313018 147978
rect 313086 147922 313142 147978
rect 311612 146942 311668 146998
rect 312714 130294 312770 130350
rect 312838 130294 312894 130350
rect 312962 130294 313018 130350
rect 313086 130294 313142 130350
rect 312714 130170 312770 130226
rect 312838 130170 312894 130226
rect 312962 130170 313018 130226
rect 313086 130170 313142 130226
rect 312714 130046 312770 130102
rect 312838 130046 312894 130102
rect 312962 130046 313018 130102
rect 313086 130046 313142 130102
rect 312714 129922 312770 129978
rect 312838 129922 312894 129978
rect 312962 129922 313018 129978
rect 313086 129922 313142 129978
rect 312714 112294 312770 112350
rect 312838 112294 312894 112350
rect 312962 112294 313018 112350
rect 313086 112294 313142 112350
rect 312714 112170 312770 112226
rect 312838 112170 312894 112226
rect 312962 112170 313018 112226
rect 313086 112170 313142 112226
rect 312714 112046 312770 112102
rect 312838 112046 312894 112102
rect 312962 112046 313018 112102
rect 313086 112046 313142 112102
rect 312714 111922 312770 111978
rect 312838 111922 312894 111978
rect 312962 111922 313018 111978
rect 313086 111922 313142 111978
rect 312714 94294 312770 94350
rect 312838 94294 312894 94350
rect 312962 94294 313018 94350
rect 313086 94294 313142 94350
rect 312714 94170 312770 94226
rect 312838 94170 312894 94226
rect 312962 94170 313018 94226
rect 313086 94170 313142 94226
rect 312714 94046 312770 94102
rect 312838 94046 312894 94102
rect 312962 94046 313018 94102
rect 313086 94046 313142 94102
rect 312714 93922 312770 93978
rect 312838 93922 312894 93978
rect 312962 93922 313018 93978
rect 313086 93922 313142 93978
rect 299528 82091 299584 82147
rect 299632 82091 299688 82147
rect 299736 82091 299792 82147
rect 299528 81987 299584 82043
rect 299632 81987 299688 82043
rect 299736 81987 299792 82043
rect 299528 81883 299584 81939
rect 299632 81883 299688 81939
rect 299736 81883 299792 81939
rect 307844 82091 307900 82147
rect 307948 82091 308004 82147
rect 308052 82091 308108 82147
rect 307844 81987 307900 82043
rect 307948 81987 308004 82043
rect 308052 81987 308108 82043
rect 307844 81883 307900 81939
rect 307948 81883 308004 81939
rect 308052 81883 308108 81939
rect 295412 76294 295468 76350
rect 295536 76294 295592 76350
rect 295412 76170 295468 76226
rect 295536 76170 295592 76226
rect 295412 76046 295468 76102
rect 295536 76046 295592 76102
rect 295412 75922 295468 75978
rect 295536 75922 295592 75978
rect 303728 76294 303784 76350
rect 303852 76294 303908 76350
rect 303728 76170 303784 76226
rect 303852 76170 303908 76226
rect 303728 76046 303784 76102
rect 303852 76046 303908 76102
rect 303728 75922 303784 75978
rect 303852 75922 303908 75978
rect 312044 76294 312100 76350
rect 312168 76294 312224 76350
rect 312044 76170 312100 76226
rect 312168 76170 312224 76226
rect 312044 76046 312100 76102
rect 312168 76046 312224 76102
rect 312044 75922 312100 75978
rect 312168 75922 312224 75978
rect 316434 154294 316490 154350
rect 316558 154294 316614 154350
rect 316682 154294 316738 154350
rect 316806 154294 316862 154350
rect 316434 154170 316490 154226
rect 316558 154170 316614 154226
rect 316682 154170 316738 154226
rect 316806 154170 316862 154226
rect 316434 154046 316490 154102
rect 316558 154046 316614 154102
rect 316682 154046 316738 154102
rect 316806 154046 316862 154102
rect 316434 153922 316490 153978
rect 316558 153922 316614 153978
rect 316682 153922 316738 153978
rect 316806 153922 316862 153978
rect 316434 136294 316490 136350
rect 316558 136294 316614 136350
rect 316682 136294 316738 136350
rect 316806 136294 316862 136350
rect 316434 136170 316490 136226
rect 316558 136170 316614 136226
rect 316682 136170 316738 136226
rect 316806 136170 316862 136226
rect 316434 136046 316490 136102
rect 316558 136046 316614 136102
rect 316682 136046 316738 136102
rect 316806 136046 316862 136102
rect 316434 135922 316490 135978
rect 316558 135922 316614 135978
rect 316682 135922 316738 135978
rect 316806 135922 316862 135978
rect 316434 118294 316490 118350
rect 316558 118294 316614 118350
rect 316682 118294 316738 118350
rect 316806 118294 316862 118350
rect 316434 118170 316490 118226
rect 316558 118170 316614 118226
rect 316682 118170 316738 118226
rect 316806 118170 316862 118226
rect 316434 118046 316490 118102
rect 316558 118046 316614 118102
rect 316682 118046 316738 118102
rect 316806 118046 316862 118102
rect 316434 117922 316490 117978
rect 316558 117922 316614 117978
rect 316682 117922 316738 117978
rect 316806 117922 316862 117978
rect 316434 100294 316490 100350
rect 316558 100294 316614 100350
rect 316682 100294 316738 100350
rect 316806 100294 316862 100350
rect 316434 100170 316490 100226
rect 316558 100170 316614 100226
rect 316682 100170 316738 100226
rect 316806 100170 316862 100226
rect 316434 100046 316490 100102
rect 316558 100046 316614 100102
rect 316682 100046 316738 100102
rect 316806 100046 316862 100102
rect 316434 99922 316490 99978
rect 316558 99922 316614 99978
rect 316682 99922 316738 99978
rect 316806 99922 316862 99978
rect 316160 82091 316216 82147
rect 316264 82091 316320 82147
rect 316368 82091 316424 82147
rect 316160 81987 316216 82043
rect 316264 81987 316320 82043
rect 316368 81987 316424 82043
rect 316160 81883 316216 81939
rect 316264 81883 316320 81939
rect 316368 81883 316424 81939
rect 324476 82091 324532 82147
rect 324580 82091 324636 82147
rect 324684 82091 324740 82147
rect 324476 81987 324532 82043
rect 324580 81987 324636 82043
rect 324684 81987 324740 82043
rect 324476 81883 324532 81939
rect 324580 81883 324636 81939
rect 324684 81883 324740 81939
rect 312714 76294 312770 76350
rect 312838 76294 312894 76350
rect 312962 76294 313018 76350
rect 313086 76294 313142 76350
rect 312714 76170 312770 76226
rect 312838 76170 312894 76226
rect 312962 76170 313018 76226
rect 313086 76170 313142 76226
rect 312714 76046 312770 76102
rect 312838 76046 312894 76102
rect 312962 76046 313018 76102
rect 313086 76046 313142 76102
rect 312714 75922 312770 75978
rect 312838 75922 312894 75978
rect 312962 75922 313018 75978
rect 313086 75922 313142 75978
rect 299570 64294 299626 64350
rect 299694 64294 299750 64350
rect 299570 64170 299626 64226
rect 299694 64170 299750 64226
rect 299570 64046 299626 64102
rect 299694 64046 299750 64102
rect 299570 63922 299626 63978
rect 299694 63922 299750 63978
rect 307886 64294 307942 64350
rect 308010 64294 308066 64350
rect 307886 64170 307942 64226
rect 308010 64170 308066 64226
rect 307886 64046 307942 64102
rect 308010 64046 308066 64102
rect 307886 63922 307942 63978
rect 308010 63922 308066 63978
rect 295412 58294 295468 58350
rect 295536 58294 295592 58350
rect 295412 58170 295468 58226
rect 295536 58170 295592 58226
rect 295412 58046 295468 58102
rect 295536 58046 295592 58102
rect 295412 57922 295468 57978
rect 295536 57922 295592 57978
rect 303728 58294 303784 58350
rect 303852 58294 303908 58350
rect 303728 58170 303784 58226
rect 303852 58170 303908 58226
rect 303728 58046 303784 58102
rect 303852 58046 303908 58102
rect 303728 57922 303784 57978
rect 303852 57922 303908 57978
rect 312044 58294 312100 58350
rect 312168 58294 312224 58350
rect 312044 58170 312100 58226
rect 312168 58170 312224 58226
rect 312044 58046 312100 58102
rect 312168 58046 312224 58102
rect 312044 57922 312100 57978
rect 312168 57922 312224 57978
rect 320360 76294 320416 76350
rect 320484 76294 320540 76350
rect 320360 76170 320416 76226
rect 320484 76170 320540 76226
rect 320360 76046 320416 76102
rect 320484 76046 320540 76102
rect 320360 75922 320416 75978
rect 320484 75922 320540 75978
rect 316202 64294 316258 64350
rect 316326 64294 316382 64350
rect 316202 64170 316258 64226
rect 316326 64170 316382 64226
rect 316202 64046 316258 64102
rect 316326 64046 316382 64102
rect 316202 63922 316258 63978
rect 316326 63922 316382 63978
rect 324518 64294 324574 64350
rect 324642 64294 324698 64350
rect 324518 64170 324574 64226
rect 324642 64170 324698 64226
rect 324518 64046 324574 64102
rect 324642 64046 324698 64102
rect 324518 63922 324574 63978
rect 324642 63922 324698 63978
rect 312714 58294 312770 58350
rect 312838 58294 312894 58350
rect 312962 58294 313018 58350
rect 313086 58294 313142 58350
rect 312714 58170 312770 58226
rect 312838 58170 312894 58226
rect 312962 58170 313018 58226
rect 313086 58170 313142 58226
rect 312714 58046 312770 58102
rect 312838 58046 312894 58102
rect 312962 58046 313018 58102
rect 313086 58046 313142 58102
rect 312714 57922 312770 57978
rect 312838 57922 312894 57978
rect 312962 57922 313018 57978
rect 313086 57922 313142 57978
rect 320360 58294 320416 58350
rect 320484 58294 320540 58350
rect 320360 58170 320416 58226
rect 320484 58170 320540 58226
rect 320360 58046 320416 58102
rect 320484 58046 320540 58102
rect 320360 57922 320416 57978
rect 320484 57922 320540 57978
rect 312714 40294 312770 40350
rect 312838 40294 312894 40350
rect 312962 40294 313018 40350
rect 313086 40294 313142 40350
rect 312714 40170 312770 40226
rect 312838 40170 312894 40226
rect 312962 40170 313018 40226
rect 313086 40170 313142 40226
rect 312714 40046 312770 40102
rect 312838 40046 312894 40102
rect 312962 40046 313018 40102
rect 313086 40046 313142 40102
rect 312714 39922 312770 39978
rect 312838 39922 312894 39978
rect 312962 39922 313018 39978
rect 313086 39922 313142 39978
rect 312714 22294 312770 22350
rect 312838 22294 312894 22350
rect 312962 22294 313018 22350
rect 313086 22294 313142 22350
rect 312714 22170 312770 22226
rect 312838 22170 312894 22226
rect 312962 22170 313018 22226
rect 313086 22170 313142 22226
rect 312714 22046 312770 22102
rect 312838 22046 312894 22102
rect 312962 22046 313018 22102
rect 313086 22046 313142 22102
rect 312714 21922 312770 21978
rect 312838 21922 312894 21978
rect 312962 21922 313018 21978
rect 313086 21922 313142 21978
rect 285714 -1176 285770 -1120
rect 285838 -1176 285894 -1120
rect 285962 -1176 286018 -1120
rect 286086 -1176 286142 -1120
rect 285714 -1300 285770 -1244
rect 285838 -1300 285894 -1244
rect 285962 -1300 286018 -1244
rect 286086 -1300 286142 -1244
rect 285714 -1424 285770 -1368
rect 285838 -1424 285894 -1368
rect 285962 -1424 286018 -1368
rect 286086 -1424 286142 -1368
rect 285714 -1548 285770 -1492
rect 285838 -1548 285894 -1492
rect 285962 -1548 286018 -1492
rect 286086 -1548 286142 -1492
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 316434 46294 316490 46350
rect 316558 46294 316614 46350
rect 316682 46294 316738 46350
rect 316806 46294 316862 46350
rect 316434 46170 316490 46226
rect 316558 46170 316614 46226
rect 316682 46170 316738 46226
rect 316806 46170 316862 46226
rect 316434 46046 316490 46102
rect 316558 46046 316614 46102
rect 316682 46046 316738 46102
rect 316806 46046 316862 46102
rect 316434 45922 316490 45978
rect 316558 45922 316614 45978
rect 316682 45922 316738 45978
rect 316806 45922 316862 45978
rect 337260 241262 337316 241318
rect 337148 240182 337204 240238
rect 337036 164582 337092 164638
rect 338604 258362 338660 258418
rect 338268 245402 338324 245458
rect 338492 247022 338548 247078
rect 338492 245042 338548 245098
rect 338380 197522 338436 197578
rect 339276 258412 339332 258418
rect 339276 258362 339332 258412
rect 338716 256562 338772 256618
rect 339388 256562 339444 256618
rect 338716 44522 338772 44578
rect 339276 253682 339332 253738
rect 339276 247022 339332 247078
rect 339388 245402 339444 245458
rect 339388 245084 339444 245098
rect 339388 245042 339444 245084
rect 339388 244916 339444 244918
rect 339388 244862 339444 244916
rect 339724 407582 339780 407638
rect 343434 400294 343490 400350
rect 343558 400294 343614 400350
rect 343682 400294 343738 400350
rect 343806 400294 343862 400350
rect 343434 400170 343490 400226
rect 343558 400170 343614 400226
rect 343682 400170 343738 400226
rect 343806 400170 343862 400226
rect 343434 400046 343490 400102
rect 343558 400046 343614 400102
rect 343682 400046 343738 400102
rect 343806 400046 343862 400102
rect 343434 399922 343490 399978
rect 343558 399922 343614 399978
rect 343682 399922 343738 399978
rect 343806 399922 343862 399978
rect 339948 397322 340004 397378
rect 339724 241622 339780 241678
rect 339612 240182 339668 240238
rect 339724 210842 339780 210898
rect 339500 157742 339556 157798
rect 339164 139382 339220 139438
rect 343196 395162 343252 395218
rect 342748 390662 342804 390718
rect 341852 380762 341908 380818
rect 340060 249902 340116 249958
rect 339948 238742 340004 238798
rect 340060 234422 340116 234478
rect 340284 193922 340340 193978
rect 340620 161162 340676 161218
rect 340284 160442 340340 160498
rect 340844 238562 340900 238618
rect 341292 241442 341348 241498
rect 341068 192302 341124 192358
rect 342076 160622 342132 160678
rect 341964 156122 342020 156178
rect 342076 149642 342132 149698
rect 347154 406294 347210 406350
rect 347278 406294 347334 406350
rect 347402 406294 347458 406350
rect 347526 406294 347582 406350
rect 347154 406170 347210 406226
rect 347278 406170 347334 406226
rect 347402 406170 347458 406226
rect 347526 406170 347582 406226
rect 347154 406046 347210 406102
rect 347278 406046 347334 406102
rect 347402 406046 347458 406102
rect 347526 406046 347582 406102
rect 347154 405922 347210 405978
rect 347278 405922 347334 405978
rect 347402 405922 347458 405978
rect 347526 405922 347582 405978
rect 343434 382294 343490 382350
rect 343558 382294 343614 382350
rect 343682 382294 343738 382350
rect 343806 382294 343862 382350
rect 343434 382170 343490 382226
rect 343558 382170 343614 382226
rect 343682 382170 343738 382226
rect 343806 382170 343862 382226
rect 343434 382046 343490 382102
rect 343558 382046 343614 382102
rect 343682 382046 343738 382102
rect 343806 382046 343862 382102
rect 343434 381922 343490 381978
rect 343558 381922 343614 381978
rect 343682 381922 343738 381978
rect 343806 381922 343862 381978
rect 344092 398582 344148 398638
rect 344204 395342 344260 395398
rect 347154 388294 347210 388350
rect 347278 388294 347334 388350
rect 347402 388294 347458 388350
rect 347526 388294 347582 388350
rect 347154 388170 347210 388226
rect 347278 388170 347334 388226
rect 347402 388170 347458 388226
rect 347526 388170 347582 388226
rect 347154 388046 347210 388102
rect 347278 388046 347334 388102
rect 347402 388046 347458 388102
rect 347526 388046 347582 388102
rect 347154 387922 347210 387978
rect 347278 387922 347334 387978
rect 347402 387922 347458 387978
rect 347526 387922 347582 387978
rect 348572 407222 348628 407278
rect 347154 370294 347210 370350
rect 347278 370294 347334 370350
rect 347402 370294 347458 370350
rect 347526 370294 347582 370350
rect 347154 370170 347210 370226
rect 347278 370170 347334 370226
rect 347402 370170 347458 370226
rect 347526 370170 347582 370226
rect 347154 370046 347210 370102
rect 347278 370046 347334 370102
rect 347402 370046 347458 370102
rect 347526 370046 347582 370102
rect 347154 369922 347210 369978
rect 347278 369922 347334 369978
rect 347402 369922 347458 369978
rect 347526 369922 347582 369978
rect 343434 364294 343490 364350
rect 343558 364294 343614 364350
rect 343682 364294 343738 364350
rect 343806 364294 343862 364350
rect 343434 364170 343490 364226
rect 343558 364170 343614 364226
rect 343682 364170 343738 364226
rect 343806 364170 343862 364226
rect 343434 364046 343490 364102
rect 343558 364046 343614 364102
rect 343682 364046 343738 364102
rect 343806 364046 343862 364102
rect 343434 363922 343490 363978
rect 343558 363922 343614 363978
rect 343682 363922 343738 363978
rect 343806 363922 343862 363978
rect 343434 346294 343490 346350
rect 343558 346294 343614 346350
rect 343682 346294 343738 346350
rect 343806 346294 343862 346350
rect 343434 346170 343490 346226
rect 343558 346170 343614 346226
rect 343682 346170 343738 346226
rect 343806 346170 343862 346226
rect 343434 346046 343490 346102
rect 343558 346046 343614 346102
rect 343682 346046 343738 346102
rect 343806 346046 343862 346102
rect 343434 345922 343490 345978
rect 343558 345922 343614 345978
rect 343682 345922 343738 345978
rect 343806 345922 343862 345978
rect 343434 328294 343490 328350
rect 343558 328294 343614 328350
rect 343682 328294 343738 328350
rect 343806 328294 343862 328350
rect 343434 328170 343490 328226
rect 343558 328170 343614 328226
rect 343682 328170 343738 328226
rect 343806 328170 343862 328226
rect 343434 328046 343490 328102
rect 343558 328046 343614 328102
rect 343682 328046 343738 328102
rect 343806 328046 343862 328102
rect 343434 327922 343490 327978
rect 343558 327922 343614 327978
rect 343682 327922 343738 327978
rect 343806 327922 343862 327978
rect 343434 310294 343490 310350
rect 343558 310294 343614 310350
rect 343682 310294 343738 310350
rect 343806 310294 343862 310350
rect 343434 310170 343490 310226
rect 343558 310170 343614 310226
rect 343682 310170 343738 310226
rect 343806 310170 343862 310226
rect 343434 310046 343490 310102
rect 343558 310046 343614 310102
rect 343682 310046 343738 310102
rect 343806 310046 343862 310102
rect 343434 309922 343490 309978
rect 343558 309922 343614 309978
rect 343682 309922 343738 309978
rect 343806 309922 343862 309978
rect 343434 292294 343490 292350
rect 343558 292294 343614 292350
rect 343682 292294 343738 292350
rect 343806 292294 343862 292350
rect 343434 292170 343490 292226
rect 343558 292170 343614 292226
rect 343682 292170 343738 292226
rect 343806 292170 343862 292226
rect 343434 292046 343490 292102
rect 343558 292046 343614 292102
rect 343682 292046 343738 292102
rect 343806 292046 343862 292102
rect 343434 291922 343490 291978
rect 343558 291922 343614 291978
rect 343682 291922 343738 291978
rect 343806 291922 343862 291978
rect 343434 274294 343490 274350
rect 343558 274294 343614 274350
rect 343682 274294 343738 274350
rect 343806 274294 343862 274350
rect 343434 274170 343490 274226
rect 343558 274170 343614 274226
rect 343682 274170 343738 274226
rect 343806 274170 343862 274226
rect 343434 274046 343490 274102
rect 343558 274046 343614 274102
rect 343682 274046 343738 274102
rect 343806 274046 343862 274102
rect 343434 273922 343490 273978
rect 343558 273922 343614 273978
rect 343682 273922 343738 273978
rect 343806 273922 343862 273978
rect 342412 241262 342468 241318
rect 342860 241082 342916 241138
rect 343434 256294 343490 256350
rect 343558 256294 343614 256350
rect 343682 256294 343738 256350
rect 343806 256294 343862 256350
rect 343434 256170 343490 256226
rect 343558 256170 343614 256226
rect 343682 256170 343738 256226
rect 343806 256170 343862 256226
rect 343434 256046 343490 256102
rect 343558 256046 343614 256102
rect 343682 256046 343738 256102
rect 343806 256046 343862 256102
rect 343434 255922 343490 255978
rect 343558 255922 343614 255978
rect 343682 255922 343738 255978
rect 343806 255922 343862 255978
rect 342636 238922 342692 238978
rect 344316 262862 344372 262918
rect 344764 241802 344820 241858
rect 344764 240362 344820 240418
rect 343434 238294 343490 238350
rect 343558 238294 343614 238350
rect 343682 238294 343738 238350
rect 343806 238294 343862 238350
rect 343434 238170 343490 238226
rect 343558 238170 343614 238226
rect 343682 238170 343738 238226
rect 343806 238170 343862 238226
rect 343434 238046 343490 238102
rect 343558 238046 343614 238102
rect 343682 238046 343738 238102
rect 343806 238046 343862 238102
rect 343434 237922 343490 237978
rect 343558 237922 343614 237978
rect 343682 237922 343738 237978
rect 343806 237922 343862 237978
rect 343434 220294 343490 220350
rect 343558 220294 343614 220350
rect 343682 220294 343738 220350
rect 343806 220294 343862 220350
rect 343434 220170 343490 220226
rect 343558 220170 343614 220226
rect 343682 220170 343738 220226
rect 343806 220170 343862 220226
rect 343434 220046 343490 220102
rect 343558 220046 343614 220102
rect 343682 220046 343738 220102
rect 343806 220046 343862 220102
rect 343434 219922 343490 219978
rect 343558 219922 343614 219978
rect 343682 219922 343738 219978
rect 343806 219922 343862 219978
rect 343434 202294 343490 202350
rect 343558 202294 343614 202350
rect 343682 202294 343738 202350
rect 343806 202294 343862 202350
rect 343434 202170 343490 202226
rect 343558 202170 343614 202226
rect 343682 202170 343738 202226
rect 343806 202170 343862 202226
rect 343434 202046 343490 202102
rect 343558 202046 343614 202102
rect 343682 202046 343738 202102
rect 343806 202046 343862 202102
rect 343434 201922 343490 201978
rect 343558 201922 343614 201978
rect 343682 201922 343738 201978
rect 343806 201922 343862 201978
rect 343434 184294 343490 184350
rect 343558 184294 343614 184350
rect 343682 184294 343738 184350
rect 343806 184294 343862 184350
rect 343434 184170 343490 184226
rect 343558 184170 343614 184226
rect 343682 184170 343738 184226
rect 343806 184170 343862 184226
rect 343434 184046 343490 184102
rect 343558 184046 343614 184102
rect 343682 184046 343738 184102
rect 343806 184046 343862 184102
rect 343434 183922 343490 183978
rect 343558 183922 343614 183978
rect 343682 183922 343738 183978
rect 343806 183922 343862 183978
rect 343434 166294 343490 166350
rect 343558 166294 343614 166350
rect 343682 166294 343738 166350
rect 343806 166294 343862 166350
rect 343434 166170 343490 166226
rect 343558 166170 343614 166226
rect 343682 166170 343738 166226
rect 343806 166170 343862 166226
rect 343434 166046 343490 166102
rect 343558 166046 343614 166102
rect 343682 166046 343738 166102
rect 343806 166046 343862 166102
rect 343434 165922 343490 165978
rect 343558 165922 343614 165978
rect 343682 165922 343738 165978
rect 343806 165922 343862 165978
rect 343434 148294 343490 148350
rect 343558 148294 343614 148350
rect 343682 148294 343738 148350
rect 343806 148294 343862 148350
rect 343434 148170 343490 148226
rect 343558 148170 343614 148226
rect 343682 148170 343738 148226
rect 343806 148170 343862 148226
rect 343434 148046 343490 148102
rect 343558 148046 343614 148102
rect 343682 148046 343738 148102
rect 343806 148046 343862 148102
rect 343434 147922 343490 147978
rect 343558 147922 343614 147978
rect 343682 147922 343738 147978
rect 343806 147922 343862 147978
rect 344092 197342 344148 197398
rect 344204 158642 344260 158698
rect 343434 130294 343490 130350
rect 343558 130294 343614 130350
rect 343682 130294 343738 130350
rect 343806 130294 343862 130350
rect 343434 130170 343490 130226
rect 343558 130170 343614 130226
rect 343682 130170 343738 130226
rect 343806 130170 343862 130226
rect 343434 130046 343490 130102
rect 343558 130046 343614 130102
rect 343682 130046 343738 130102
rect 343806 130046 343862 130102
rect 343434 129922 343490 129978
rect 343558 129922 343614 129978
rect 343682 129922 343738 129978
rect 343806 129922 343862 129978
rect 343434 112294 343490 112350
rect 343558 112294 343614 112350
rect 343682 112294 343738 112350
rect 343806 112294 343862 112350
rect 343434 112170 343490 112226
rect 343558 112170 343614 112226
rect 343682 112170 343738 112226
rect 343806 112170 343862 112226
rect 343434 112046 343490 112102
rect 343558 112046 343614 112102
rect 343682 112046 343738 112102
rect 343806 112046 343862 112102
rect 343434 111922 343490 111978
rect 343558 111922 343614 111978
rect 343682 111922 343738 111978
rect 343806 111922 343862 111978
rect 342524 94922 342580 94978
rect 345324 155402 345380 155458
rect 345548 240362 345604 240418
rect 345772 211022 345828 211078
rect 343434 94294 343490 94350
rect 343558 94294 343614 94350
rect 343682 94294 343738 94350
rect 343806 94294 343862 94350
rect 343434 94170 343490 94226
rect 343558 94170 343614 94226
rect 343682 94170 343738 94226
rect 343806 94170 343862 94226
rect 343434 94046 343490 94102
rect 343558 94046 343614 94102
rect 343682 94046 343738 94102
rect 343806 94046 343862 94102
rect 343434 93922 343490 93978
rect 343558 93922 343614 93978
rect 343682 93922 343738 93978
rect 343806 93922 343862 93978
rect 343434 76294 343490 76350
rect 343558 76294 343614 76350
rect 343682 76294 343738 76350
rect 343806 76294 343862 76350
rect 343434 76170 343490 76226
rect 343558 76170 343614 76226
rect 343682 76170 343738 76226
rect 343806 76170 343862 76226
rect 343434 76046 343490 76102
rect 343558 76046 343614 76102
rect 343682 76046 343738 76102
rect 343806 76046 343862 76102
rect 343434 75922 343490 75978
rect 343558 75922 343614 75978
rect 343682 75922 343738 75978
rect 343806 75922 343862 75978
rect 343434 58294 343490 58350
rect 343558 58294 343614 58350
rect 343682 58294 343738 58350
rect 343806 58294 343862 58350
rect 343434 58170 343490 58226
rect 343558 58170 343614 58226
rect 343682 58170 343738 58226
rect 343806 58170 343862 58226
rect 343434 58046 343490 58102
rect 343558 58046 343614 58102
rect 343682 58046 343738 58102
rect 343806 58046 343862 58102
rect 343434 57922 343490 57978
rect 343558 57922 343614 57978
rect 343682 57922 343738 57978
rect 343806 57922 343862 57978
rect 340172 41102 340228 41158
rect 346108 234242 346164 234298
rect 346332 160802 346388 160858
rect 346108 157382 346164 157438
rect 346556 150362 346612 150418
rect 346892 162782 346948 162838
rect 347154 352294 347210 352350
rect 347278 352294 347334 352350
rect 347402 352294 347458 352350
rect 347526 352294 347582 352350
rect 347154 352170 347210 352226
rect 347278 352170 347334 352226
rect 347402 352170 347458 352226
rect 347526 352170 347582 352226
rect 347154 352046 347210 352102
rect 347278 352046 347334 352102
rect 347402 352046 347458 352102
rect 347526 352046 347582 352102
rect 347154 351922 347210 351978
rect 347278 351922 347334 351978
rect 347402 351922 347458 351978
rect 347526 351922 347582 351978
rect 347154 334294 347210 334350
rect 347278 334294 347334 334350
rect 347402 334294 347458 334350
rect 347526 334294 347582 334350
rect 347154 334170 347210 334226
rect 347278 334170 347334 334226
rect 347402 334170 347458 334226
rect 347526 334170 347582 334226
rect 347154 334046 347210 334102
rect 347278 334046 347334 334102
rect 347402 334046 347458 334102
rect 347526 334046 347582 334102
rect 347154 333922 347210 333978
rect 347278 333922 347334 333978
rect 347402 333922 347458 333978
rect 347526 333922 347582 333978
rect 347154 316294 347210 316350
rect 347278 316294 347334 316350
rect 347402 316294 347458 316350
rect 347526 316294 347582 316350
rect 347154 316170 347210 316226
rect 347278 316170 347334 316226
rect 347402 316170 347458 316226
rect 347526 316170 347582 316226
rect 347154 316046 347210 316102
rect 347278 316046 347334 316102
rect 347402 316046 347458 316102
rect 347526 316046 347582 316102
rect 347154 315922 347210 315978
rect 347278 315922 347334 315978
rect 347402 315922 347458 315978
rect 347526 315922 347582 315978
rect 347154 298294 347210 298350
rect 347278 298294 347334 298350
rect 347402 298294 347458 298350
rect 347526 298294 347582 298350
rect 347154 298170 347210 298226
rect 347278 298170 347334 298226
rect 347402 298170 347458 298226
rect 347526 298170 347582 298226
rect 347154 298046 347210 298102
rect 347278 298046 347334 298102
rect 347402 298046 347458 298102
rect 347526 298046 347582 298102
rect 347154 297922 347210 297978
rect 347278 297922 347334 297978
rect 347402 297922 347458 297978
rect 347526 297922 347582 297978
rect 347154 280294 347210 280350
rect 347278 280294 347334 280350
rect 347402 280294 347458 280350
rect 347526 280294 347582 280350
rect 347154 280170 347210 280226
rect 347278 280170 347334 280226
rect 347402 280170 347458 280226
rect 347526 280170 347582 280226
rect 347154 280046 347210 280102
rect 347278 280046 347334 280102
rect 347402 280046 347458 280102
rect 347526 280046 347582 280102
rect 347154 279922 347210 279978
rect 347278 279922 347334 279978
rect 347402 279922 347458 279978
rect 347526 279922 347582 279978
rect 347154 262294 347210 262350
rect 347278 262294 347334 262350
rect 347402 262294 347458 262350
rect 347526 262294 347582 262350
rect 347154 262170 347210 262226
rect 347278 262170 347334 262226
rect 347402 262170 347458 262226
rect 347526 262170 347582 262226
rect 347154 262046 347210 262102
rect 347278 262046 347334 262102
rect 347402 262046 347458 262102
rect 347526 262046 347582 262102
rect 347154 261922 347210 261978
rect 347278 261922 347334 261978
rect 347402 261922 347458 261978
rect 347526 261922 347582 261978
rect 347154 244294 347210 244350
rect 347278 244294 347334 244350
rect 347402 244294 347458 244350
rect 347526 244294 347582 244350
rect 347154 244170 347210 244226
rect 347278 244170 347334 244226
rect 347402 244170 347458 244226
rect 347526 244170 347582 244226
rect 347154 244046 347210 244102
rect 347278 244046 347334 244102
rect 347402 244046 347458 244102
rect 347526 244046 347582 244102
rect 347154 243922 347210 243978
rect 347278 243922 347334 243978
rect 347402 243922 347458 243978
rect 347526 243922 347582 243978
rect 347154 226294 347210 226350
rect 347278 226294 347334 226350
rect 347402 226294 347458 226350
rect 347526 226294 347582 226350
rect 347154 226170 347210 226226
rect 347278 226170 347334 226226
rect 347402 226170 347458 226226
rect 347526 226170 347582 226226
rect 347154 226046 347210 226102
rect 347278 226046 347334 226102
rect 347402 226046 347458 226102
rect 347526 226046 347582 226102
rect 347154 225922 347210 225978
rect 347278 225922 347334 225978
rect 347402 225922 347458 225978
rect 347526 225922 347582 225978
rect 347154 208294 347210 208350
rect 347278 208294 347334 208350
rect 347402 208294 347458 208350
rect 347526 208294 347582 208350
rect 347154 208170 347210 208226
rect 347278 208170 347334 208226
rect 347402 208170 347458 208226
rect 347526 208170 347582 208226
rect 347154 208046 347210 208102
rect 347278 208046 347334 208102
rect 347402 208046 347458 208102
rect 347526 208046 347582 208102
rect 347154 207922 347210 207978
rect 347278 207922 347334 207978
rect 347402 207922 347458 207978
rect 347526 207922 347582 207978
rect 347154 190294 347210 190350
rect 347278 190294 347334 190350
rect 347402 190294 347458 190350
rect 347526 190294 347582 190350
rect 347154 190170 347210 190226
rect 347278 190170 347334 190226
rect 347402 190170 347458 190226
rect 347526 190170 347582 190226
rect 347154 190046 347210 190102
rect 347278 190046 347334 190102
rect 347402 190046 347458 190102
rect 347526 190046 347582 190102
rect 347154 189922 347210 189978
rect 347278 189922 347334 189978
rect 347402 189922 347458 189978
rect 347526 189922 347582 189978
rect 347154 172294 347210 172350
rect 347278 172294 347334 172350
rect 347402 172294 347458 172350
rect 347526 172294 347582 172350
rect 347154 172170 347210 172226
rect 347278 172170 347334 172226
rect 347402 172170 347458 172226
rect 347526 172170 347582 172226
rect 347154 172046 347210 172102
rect 347278 172046 347334 172102
rect 347402 172046 347458 172102
rect 347526 172046 347582 172102
rect 347154 171922 347210 171978
rect 347278 171922 347334 171978
rect 347402 171922 347458 171978
rect 347526 171922 347582 171978
rect 346892 157922 346948 157978
rect 346780 148562 346836 148618
rect 348460 162062 348516 162118
rect 347154 154294 347210 154350
rect 347278 154294 347334 154350
rect 347402 154294 347458 154350
rect 347526 154294 347582 154350
rect 347154 154170 347210 154226
rect 347278 154170 347334 154226
rect 347402 154170 347458 154226
rect 347526 154170 347582 154226
rect 347154 154046 347210 154102
rect 347278 154046 347334 154102
rect 347402 154046 347458 154102
rect 347526 154046 347582 154102
rect 347154 153922 347210 153978
rect 347278 153922 347334 153978
rect 347402 153922 347458 153978
rect 347526 153922 347582 153978
rect 347154 136294 347210 136350
rect 347278 136294 347334 136350
rect 347402 136294 347458 136350
rect 347526 136294 347582 136350
rect 347154 136170 347210 136226
rect 347278 136170 347334 136226
rect 347402 136170 347458 136226
rect 347526 136170 347582 136226
rect 347154 136046 347210 136102
rect 347278 136046 347334 136102
rect 347402 136046 347458 136102
rect 347526 136046 347582 136102
rect 347154 135922 347210 135978
rect 347278 135922 347334 135978
rect 347402 135922 347458 135978
rect 347526 135922 347582 135978
rect 347154 118294 347210 118350
rect 347278 118294 347334 118350
rect 347402 118294 347458 118350
rect 347526 118294 347582 118350
rect 347154 118170 347210 118226
rect 347278 118170 347334 118226
rect 347402 118170 347458 118226
rect 347526 118170 347582 118226
rect 347154 118046 347210 118102
rect 347278 118046 347334 118102
rect 347402 118046 347458 118102
rect 347526 118046 347582 118102
rect 347154 117922 347210 117978
rect 347278 117922 347334 117978
rect 347402 117922 347458 117978
rect 347526 117922 347582 117978
rect 347154 100294 347210 100350
rect 347278 100294 347334 100350
rect 347402 100294 347458 100350
rect 347526 100294 347582 100350
rect 347154 100170 347210 100226
rect 347278 100170 347334 100226
rect 347402 100170 347458 100226
rect 347526 100170 347582 100226
rect 347154 100046 347210 100102
rect 347278 100046 347334 100102
rect 347402 100046 347458 100102
rect 347526 100046 347582 100102
rect 347154 99922 347210 99978
rect 347278 99922 347334 99978
rect 347402 99922 347458 99978
rect 347526 99922 347582 99978
rect 348684 152522 348740 152578
rect 350140 151982 350196 152038
rect 350028 147662 350084 147718
rect 349356 145682 349412 145738
rect 350364 150542 350420 150598
rect 350588 152162 350644 152218
rect 350812 163682 350868 163738
rect 350812 146042 350868 146098
rect 351820 167282 351876 167338
rect 353836 406862 353892 406918
rect 353612 406682 353668 406738
rect 355292 407042 355348 407098
rect 355180 397322 355236 397378
rect 355068 397142 355124 397198
rect 355292 394982 355348 395038
rect 357756 409562 357812 409618
rect 356076 409022 356132 409078
rect 355740 400562 355796 400618
rect 356076 396962 356132 397018
rect 356412 392462 356468 392518
rect 356524 392282 356580 392338
rect 356076 391022 356132 391078
rect 356636 390842 356692 390898
rect 351036 141002 351092 141058
rect 351932 143882 351988 143938
rect 352044 140822 352100 140878
rect 352492 144242 352548 144298
rect 352604 144422 352660 144478
rect 352604 143882 352660 143938
rect 352940 262862 352996 262918
rect 353500 234602 353556 234658
rect 353500 162422 353556 162478
rect 353612 157562 353668 157618
rect 352716 142622 352772 142678
rect 354284 165482 354340 165538
rect 354396 162242 354452 162298
rect 354172 158822 354228 158878
rect 354956 164042 355012 164098
rect 355068 163862 355124 163918
rect 355404 236628 355460 236638
rect 355404 236582 355460 236628
rect 355404 213542 355460 213598
rect 355292 159542 355348 159598
rect 355180 155582 355236 155638
rect 353948 98162 354004 98218
rect 356636 236582 356692 236638
rect 356524 167282 356580 167338
rect 356076 164762 356132 164818
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 466314 562294 466370 562350
rect 466438 562294 466494 562350
rect 466562 562294 466618 562350
rect 466686 562294 466742 562350
rect 466314 562170 466370 562226
rect 466438 562170 466494 562226
rect 466562 562170 466618 562226
rect 466686 562170 466742 562226
rect 466314 562046 466370 562102
rect 466438 562046 466494 562102
rect 466562 562046 466618 562102
rect 466686 562046 466742 562102
rect 466314 561922 466370 561978
rect 466438 561922 466494 561978
rect 466562 561922 466618 561978
rect 466686 561922 466742 561978
rect 455638 550294 455694 550350
rect 455762 550294 455818 550350
rect 455638 550170 455694 550226
rect 455762 550170 455818 550226
rect 455638 550046 455694 550102
rect 455762 550046 455818 550102
rect 455638 549922 455694 549978
rect 455762 549922 455818 549978
rect 466314 544294 466370 544350
rect 466438 544294 466494 544350
rect 466562 544294 466618 544350
rect 466686 544294 466742 544350
rect 466314 544170 466370 544226
rect 466438 544170 466494 544226
rect 466562 544170 466618 544226
rect 466686 544170 466742 544226
rect 466314 544046 466370 544102
rect 466438 544046 466494 544102
rect 466562 544046 466618 544102
rect 466686 544046 466742 544102
rect 466314 543922 466370 543978
rect 466438 543922 466494 543978
rect 466562 543922 466618 543978
rect 466686 543922 466742 543978
rect 455638 532294 455694 532350
rect 455762 532294 455818 532350
rect 455638 532170 455694 532226
rect 455762 532170 455818 532226
rect 455638 532046 455694 532102
rect 455762 532046 455818 532102
rect 455638 531922 455694 531978
rect 455762 531922 455818 531978
rect 466314 526294 466370 526350
rect 466438 526294 466494 526350
rect 466562 526294 466618 526350
rect 466686 526294 466742 526350
rect 466314 526170 466370 526226
rect 466438 526170 466494 526226
rect 466562 526170 466618 526226
rect 466686 526170 466742 526226
rect 466314 526046 466370 526102
rect 466438 526046 466494 526102
rect 466562 526046 466618 526102
rect 466686 526046 466742 526102
rect 466314 525922 466370 525978
rect 466438 525922 466494 525978
rect 466562 525922 466618 525978
rect 466686 525922 466742 525978
rect 455638 514294 455694 514350
rect 455762 514294 455818 514350
rect 455638 514170 455694 514226
rect 455762 514170 455818 514226
rect 455638 514046 455694 514102
rect 455762 514046 455818 514102
rect 455638 513922 455694 513978
rect 455762 513922 455818 513978
rect 466314 508294 466370 508350
rect 466438 508294 466494 508350
rect 466562 508294 466618 508350
rect 466686 508294 466742 508350
rect 466314 508170 466370 508226
rect 466438 508170 466494 508226
rect 466562 508170 466618 508226
rect 466686 508170 466742 508226
rect 466314 508046 466370 508102
rect 466438 508046 466494 508102
rect 466562 508046 466618 508102
rect 466686 508046 466742 508102
rect 466314 507922 466370 507978
rect 466438 507922 466494 507978
rect 466562 507922 466618 507978
rect 466686 507922 466742 507978
rect 455638 496294 455694 496350
rect 455762 496294 455818 496350
rect 455638 496170 455694 496226
rect 455762 496170 455818 496226
rect 455638 496046 455694 496102
rect 455762 496046 455818 496102
rect 455638 495922 455694 495978
rect 455762 495922 455818 495978
rect 466314 490294 466370 490350
rect 466438 490294 466494 490350
rect 466562 490294 466618 490350
rect 466686 490294 466742 490350
rect 466314 490170 466370 490226
rect 466438 490170 466494 490226
rect 466562 490170 466618 490226
rect 466686 490170 466742 490226
rect 466314 490046 466370 490102
rect 466438 490046 466494 490102
rect 466562 490046 466618 490102
rect 466686 490046 466742 490102
rect 466314 489922 466370 489978
rect 466438 489922 466494 489978
rect 466562 489922 466618 489978
rect 466686 489922 466742 489978
rect 455638 478294 455694 478350
rect 455762 478294 455818 478350
rect 455638 478170 455694 478226
rect 455762 478170 455818 478226
rect 455638 478046 455694 478102
rect 455762 478046 455818 478102
rect 455638 477922 455694 477978
rect 455762 477922 455818 477978
rect 466314 472294 466370 472350
rect 466438 472294 466494 472350
rect 466562 472294 466618 472350
rect 466686 472294 466742 472350
rect 466314 472170 466370 472226
rect 466438 472170 466494 472226
rect 466562 472170 466618 472226
rect 466686 472170 466742 472226
rect 466314 472046 466370 472102
rect 466438 472046 466494 472102
rect 466562 472046 466618 472102
rect 466686 472046 466742 472102
rect 466314 471922 466370 471978
rect 466438 471922 466494 471978
rect 466562 471922 466618 471978
rect 466686 471922 466742 471978
rect 455638 460294 455694 460350
rect 455762 460294 455818 460350
rect 455638 460170 455694 460226
rect 455762 460170 455818 460226
rect 455638 460046 455694 460102
rect 455762 460046 455818 460102
rect 455638 459922 455694 459978
rect 455762 459922 455818 459978
rect 466314 454294 466370 454350
rect 466438 454294 466494 454350
rect 466562 454294 466618 454350
rect 466686 454294 466742 454350
rect 466314 454170 466370 454226
rect 466438 454170 466494 454226
rect 466562 454170 466618 454226
rect 466686 454170 466742 454226
rect 466314 454046 466370 454102
rect 466438 454046 466494 454102
rect 466562 454046 466618 454102
rect 466686 454046 466742 454102
rect 466314 453922 466370 453978
rect 466438 453922 466494 453978
rect 466562 453922 466618 453978
rect 466686 453922 466742 453978
rect 455638 442294 455694 442350
rect 455762 442294 455818 442350
rect 455638 442170 455694 442226
rect 455762 442170 455818 442226
rect 455638 442046 455694 442102
rect 455762 442046 455818 442102
rect 455638 441922 455694 441978
rect 455762 441922 455818 441978
rect 466314 436294 466370 436350
rect 466438 436294 466494 436350
rect 466562 436294 466618 436350
rect 466686 436294 466742 436350
rect 466314 436170 466370 436226
rect 466438 436170 466494 436226
rect 466562 436170 466618 436226
rect 466686 436170 466742 436226
rect 466314 436046 466370 436102
rect 466438 436046 466494 436102
rect 466562 436046 466618 436102
rect 466686 436046 466742 436102
rect 466314 435922 466370 435978
rect 466438 435922 466494 435978
rect 466562 435922 466618 435978
rect 466686 435922 466742 435978
rect 446012 428462 446068 428518
rect 444892 407222 444948 407278
rect 455638 424294 455694 424350
rect 455762 424294 455818 424350
rect 455638 424170 455694 424226
rect 455762 424170 455818 424226
rect 455638 424046 455694 424102
rect 455762 424046 455818 424102
rect 455638 423922 455694 423978
rect 455762 423922 455818 423978
rect 466314 418294 466370 418350
rect 466438 418294 466494 418350
rect 466562 418294 466618 418350
rect 466686 418294 466742 418350
rect 466314 418170 466370 418226
rect 466438 418170 466494 418226
rect 466562 418170 466618 418226
rect 466686 418170 466742 418226
rect 466314 418046 466370 418102
rect 466438 418046 466494 418102
rect 466562 418046 466618 418102
rect 466686 418046 466742 418102
rect 466314 417922 466370 417978
rect 466438 417922 466494 417978
rect 466562 417922 466618 417978
rect 466686 417922 466742 417978
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 470034 568294 470090 568350
rect 470158 568294 470214 568350
rect 470282 568294 470338 568350
rect 470406 568294 470462 568350
rect 470034 568170 470090 568226
rect 470158 568170 470214 568226
rect 470282 568170 470338 568226
rect 470406 568170 470462 568226
rect 470034 568046 470090 568102
rect 470158 568046 470214 568102
rect 470282 568046 470338 568102
rect 470406 568046 470462 568102
rect 470034 567922 470090 567978
rect 470158 567922 470214 567978
rect 470282 567922 470338 567978
rect 470406 567922 470462 567978
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 470998 562294 471054 562350
rect 471122 562294 471178 562350
rect 470998 562170 471054 562226
rect 471122 562170 471178 562226
rect 470998 562046 471054 562102
rect 471122 562046 471178 562102
rect 470998 561922 471054 561978
rect 471122 561922 471178 561978
rect 497034 562294 497090 562350
rect 497158 562294 497214 562350
rect 497282 562294 497338 562350
rect 497406 562294 497462 562350
rect 497034 562170 497090 562226
rect 497158 562170 497214 562226
rect 497282 562170 497338 562226
rect 497406 562170 497462 562226
rect 497034 562046 497090 562102
rect 497158 562046 497214 562102
rect 497282 562046 497338 562102
rect 497406 562046 497462 562102
rect 497034 561922 497090 561978
rect 497158 561922 497214 561978
rect 497282 561922 497338 561978
rect 497406 561922 497462 561978
rect 470034 550294 470090 550350
rect 470158 550294 470214 550350
rect 470282 550294 470338 550350
rect 470406 550294 470462 550350
rect 470034 550170 470090 550226
rect 470158 550170 470214 550226
rect 470282 550170 470338 550226
rect 470406 550170 470462 550226
rect 470034 550046 470090 550102
rect 470158 550046 470214 550102
rect 470282 550046 470338 550102
rect 470406 550046 470462 550102
rect 470034 549922 470090 549978
rect 470158 549922 470214 549978
rect 470282 549922 470338 549978
rect 470406 549922 470462 549978
rect 486358 550294 486414 550350
rect 486482 550294 486538 550350
rect 486358 550170 486414 550226
rect 486482 550170 486538 550226
rect 486358 550046 486414 550102
rect 486482 550046 486538 550102
rect 486358 549922 486414 549978
rect 486482 549922 486538 549978
rect 470998 544294 471054 544350
rect 471122 544294 471178 544350
rect 470998 544170 471054 544226
rect 471122 544170 471178 544226
rect 470998 544046 471054 544102
rect 471122 544046 471178 544102
rect 470998 543922 471054 543978
rect 471122 543922 471178 543978
rect 497034 544294 497090 544350
rect 497158 544294 497214 544350
rect 497282 544294 497338 544350
rect 497406 544294 497462 544350
rect 497034 544170 497090 544226
rect 497158 544170 497214 544226
rect 497282 544170 497338 544226
rect 497406 544170 497462 544226
rect 497034 544046 497090 544102
rect 497158 544046 497214 544102
rect 497282 544046 497338 544102
rect 497406 544046 497462 544102
rect 497034 543922 497090 543978
rect 497158 543922 497214 543978
rect 497282 543922 497338 543978
rect 497406 543922 497462 543978
rect 470034 532294 470090 532350
rect 470158 532294 470214 532350
rect 470282 532294 470338 532350
rect 470406 532294 470462 532350
rect 470034 532170 470090 532226
rect 470158 532170 470214 532226
rect 470282 532170 470338 532226
rect 470406 532170 470462 532226
rect 470034 532046 470090 532102
rect 470158 532046 470214 532102
rect 470282 532046 470338 532102
rect 470406 532046 470462 532102
rect 470034 531922 470090 531978
rect 470158 531922 470214 531978
rect 470282 531922 470338 531978
rect 470406 531922 470462 531978
rect 486358 532294 486414 532350
rect 486482 532294 486538 532350
rect 486358 532170 486414 532226
rect 486482 532170 486538 532226
rect 486358 532046 486414 532102
rect 486482 532046 486538 532102
rect 486358 531922 486414 531978
rect 486482 531922 486538 531978
rect 470998 526294 471054 526350
rect 471122 526294 471178 526350
rect 470998 526170 471054 526226
rect 471122 526170 471178 526226
rect 470998 526046 471054 526102
rect 471122 526046 471178 526102
rect 470998 525922 471054 525978
rect 471122 525922 471178 525978
rect 497034 526294 497090 526350
rect 497158 526294 497214 526350
rect 497282 526294 497338 526350
rect 497406 526294 497462 526350
rect 497034 526170 497090 526226
rect 497158 526170 497214 526226
rect 497282 526170 497338 526226
rect 497406 526170 497462 526226
rect 497034 526046 497090 526102
rect 497158 526046 497214 526102
rect 497282 526046 497338 526102
rect 497406 526046 497462 526102
rect 497034 525922 497090 525978
rect 497158 525922 497214 525978
rect 497282 525922 497338 525978
rect 497406 525922 497462 525978
rect 470034 514294 470090 514350
rect 470158 514294 470214 514350
rect 470282 514294 470338 514350
rect 470406 514294 470462 514350
rect 470034 514170 470090 514226
rect 470158 514170 470214 514226
rect 470282 514170 470338 514226
rect 470406 514170 470462 514226
rect 470034 514046 470090 514102
rect 470158 514046 470214 514102
rect 470282 514046 470338 514102
rect 470406 514046 470462 514102
rect 470034 513922 470090 513978
rect 470158 513922 470214 513978
rect 470282 513922 470338 513978
rect 470406 513922 470462 513978
rect 486358 514294 486414 514350
rect 486482 514294 486538 514350
rect 486358 514170 486414 514226
rect 486482 514170 486538 514226
rect 486358 514046 486414 514102
rect 486482 514046 486538 514102
rect 486358 513922 486414 513978
rect 486482 513922 486538 513978
rect 470998 508294 471054 508350
rect 471122 508294 471178 508350
rect 470998 508170 471054 508226
rect 471122 508170 471178 508226
rect 470998 508046 471054 508102
rect 471122 508046 471178 508102
rect 470998 507922 471054 507978
rect 471122 507922 471178 507978
rect 497034 508294 497090 508350
rect 497158 508294 497214 508350
rect 497282 508294 497338 508350
rect 497406 508294 497462 508350
rect 497034 508170 497090 508226
rect 497158 508170 497214 508226
rect 497282 508170 497338 508226
rect 497406 508170 497462 508226
rect 497034 508046 497090 508102
rect 497158 508046 497214 508102
rect 497282 508046 497338 508102
rect 497406 508046 497462 508102
rect 497034 507922 497090 507978
rect 497158 507922 497214 507978
rect 497282 507922 497338 507978
rect 497406 507922 497462 507978
rect 470034 496294 470090 496350
rect 470158 496294 470214 496350
rect 470282 496294 470338 496350
rect 470406 496294 470462 496350
rect 470034 496170 470090 496226
rect 470158 496170 470214 496226
rect 470282 496170 470338 496226
rect 470406 496170 470462 496226
rect 470034 496046 470090 496102
rect 470158 496046 470214 496102
rect 470282 496046 470338 496102
rect 470406 496046 470462 496102
rect 470034 495922 470090 495978
rect 470158 495922 470214 495978
rect 470282 495922 470338 495978
rect 470406 495922 470462 495978
rect 486358 496294 486414 496350
rect 486482 496294 486538 496350
rect 486358 496170 486414 496226
rect 486482 496170 486538 496226
rect 486358 496046 486414 496102
rect 486482 496046 486538 496102
rect 486358 495922 486414 495978
rect 486482 495922 486538 495978
rect 470998 490294 471054 490350
rect 471122 490294 471178 490350
rect 470998 490170 471054 490226
rect 471122 490170 471178 490226
rect 470998 490046 471054 490102
rect 471122 490046 471178 490102
rect 470998 489922 471054 489978
rect 471122 489922 471178 489978
rect 497034 490294 497090 490350
rect 497158 490294 497214 490350
rect 497282 490294 497338 490350
rect 497406 490294 497462 490350
rect 497034 490170 497090 490226
rect 497158 490170 497214 490226
rect 497282 490170 497338 490226
rect 497406 490170 497462 490226
rect 497034 490046 497090 490102
rect 497158 490046 497214 490102
rect 497282 490046 497338 490102
rect 497406 490046 497462 490102
rect 497034 489922 497090 489978
rect 497158 489922 497214 489978
rect 497282 489922 497338 489978
rect 497406 489922 497462 489978
rect 470034 478294 470090 478350
rect 470158 478294 470214 478350
rect 470282 478294 470338 478350
rect 470406 478294 470462 478350
rect 470034 478170 470090 478226
rect 470158 478170 470214 478226
rect 470282 478170 470338 478226
rect 470406 478170 470462 478226
rect 470034 478046 470090 478102
rect 470158 478046 470214 478102
rect 470282 478046 470338 478102
rect 470406 478046 470462 478102
rect 470034 477922 470090 477978
rect 470158 477922 470214 477978
rect 470282 477922 470338 477978
rect 470406 477922 470462 477978
rect 486358 478294 486414 478350
rect 486482 478294 486538 478350
rect 486358 478170 486414 478226
rect 486482 478170 486538 478226
rect 486358 478046 486414 478102
rect 486482 478046 486538 478102
rect 486358 477922 486414 477978
rect 486482 477922 486538 477978
rect 470998 472294 471054 472350
rect 471122 472294 471178 472350
rect 470998 472170 471054 472226
rect 471122 472170 471178 472226
rect 470998 472046 471054 472102
rect 471122 472046 471178 472102
rect 470998 471922 471054 471978
rect 471122 471922 471178 471978
rect 497034 472294 497090 472350
rect 497158 472294 497214 472350
rect 497282 472294 497338 472350
rect 497406 472294 497462 472350
rect 497034 472170 497090 472226
rect 497158 472170 497214 472226
rect 497282 472170 497338 472226
rect 497406 472170 497462 472226
rect 497034 472046 497090 472102
rect 497158 472046 497214 472102
rect 497282 472046 497338 472102
rect 497406 472046 497462 472102
rect 497034 471922 497090 471978
rect 497158 471922 497214 471978
rect 497282 471922 497338 471978
rect 497406 471922 497462 471978
rect 470034 460294 470090 460350
rect 470158 460294 470214 460350
rect 470282 460294 470338 460350
rect 470406 460294 470462 460350
rect 470034 460170 470090 460226
rect 470158 460170 470214 460226
rect 470282 460170 470338 460226
rect 470406 460170 470462 460226
rect 470034 460046 470090 460102
rect 470158 460046 470214 460102
rect 470282 460046 470338 460102
rect 470406 460046 470462 460102
rect 470034 459922 470090 459978
rect 470158 459922 470214 459978
rect 470282 459922 470338 459978
rect 470406 459922 470462 459978
rect 486358 460294 486414 460350
rect 486482 460294 486538 460350
rect 486358 460170 486414 460226
rect 486482 460170 486538 460226
rect 486358 460046 486414 460102
rect 486482 460046 486538 460102
rect 486358 459922 486414 459978
rect 486482 459922 486538 459978
rect 470998 454294 471054 454350
rect 471122 454294 471178 454350
rect 470998 454170 471054 454226
rect 471122 454170 471178 454226
rect 470998 454046 471054 454102
rect 471122 454046 471178 454102
rect 470998 453922 471054 453978
rect 471122 453922 471178 453978
rect 497034 454294 497090 454350
rect 497158 454294 497214 454350
rect 497282 454294 497338 454350
rect 497406 454294 497462 454350
rect 497034 454170 497090 454226
rect 497158 454170 497214 454226
rect 497282 454170 497338 454226
rect 497406 454170 497462 454226
rect 497034 454046 497090 454102
rect 497158 454046 497214 454102
rect 497282 454046 497338 454102
rect 497406 454046 497462 454102
rect 497034 453922 497090 453978
rect 497158 453922 497214 453978
rect 497282 453922 497338 453978
rect 497406 453922 497462 453978
rect 470034 442294 470090 442350
rect 470158 442294 470214 442350
rect 470282 442294 470338 442350
rect 470406 442294 470462 442350
rect 470034 442170 470090 442226
rect 470158 442170 470214 442226
rect 470282 442170 470338 442226
rect 470406 442170 470462 442226
rect 470034 442046 470090 442102
rect 470158 442046 470214 442102
rect 470282 442046 470338 442102
rect 470406 442046 470462 442102
rect 470034 441922 470090 441978
rect 470158 441922 470214 441978
rect 470282 441922 470338 441978
rect 470406 441922 470462 441978
rect 486358 442294 486414 442350
rect 486482 442294 486538 442350
rect 486358 442170 486414 442226
rect 486482 442170 486538 442226
rect 486358 442046 486414 442102
rect 486482 442046 486538 442102
rect 486358 441922 486414 441978
rect 486482 441922 486538 441978
rect 470998 436294 471054 436350
rect 471122 436294 471178 436350
rect 470998 436170 471054 436226
rect 471122 436170 471178 436226
rect 470998 436046 471054 436102
rect 471122 436046 471178 436102
rect 470998 435922 471054 435978
rect 471122 435922 471178 435978
rect 497034 436294 497090 436350
rect 497158 436294 497214 436350
rect 497282 436294 497338 436350
rect 497406 436294 497462 436350
rect 497034 436170 497090 436226
rect 497158 436170 497214 436226
rect 497282 436170 497338 436226
rect 497406 436170 497462 436226
rect 497034 436046 497090 436102
rect 497158 436046 497214 436102
rect 497282 436046 497338 436102
rect 497406 436046 497462 436102
rect 497034 435922 497090 435978
rect 497158 435922 497214 435978
rect 497282 435922 497338 435978
rect 497406 435922 497462 435978
rect 470034 424294 470090 424350
rect 470158 424294 470214 424350
rect 470282 424294 470338 424350
rect 470406 424294 470462 424350
rect 470034 424170 470090 424226
rect 470158 424170 470214 424226
rect 470282 424170 470338 424226
rect 470406 424170 470462 424226
rect 470034 424046 470090 424102
rect 470158 424046 470214 424102
rect 470282 424046 470338 424102
rect 470406 424046 470462 424102
rect 470034 423922 470090 423978
rect 470158 423922 470214 423978
rect 470282 423922 470338 423978
rect 470406 423922 470462 423978
rect 466314 400294 466370 400350
rect 466438 400294 466494 400350
rect 466562 400294 466618 400350
rect 466686 400294 466742 400350
rect 466314 400170 466370 400226
rect 466438 400170 466494 400226
rect 466562 400170 466618 400226
rect 466686 400170 466742 400226
rect 466314 400046 466370 400102
rect 466438 400046 466494 400102
rect 466562 400046 466618 400102
rect 466686 400046 466742 400102
rect 466314 399922 466370 399978
rect 466438 399922 466494 399978
rect 466562 399922 466618 399978
rect 466686 399922 466742 399978
rect 486358 424294 486414 424350
rect 486482 424294 486538 424350
rect 486358 424170 486414 424226
rect 486482 424170 486538 424226
rect 486358 424046 486414 424102
rect 486482 424046 486538 424102
rect 486358 423922 486414 423978
rect 486482 423922 486538 423978
rect 470998 418294 471054 418350
rect 471122 418294 471178 418350
rect 470998 418170 471054 418226
rect 471122 418170 471178 418226
rect 470998 418046 471054 418102
rect 471122 418046 471178 418102
rect 470998 417922 471054 417978
rect 471122 417922 471178 417978
rect 497034 418294 497090 418350
rect 497158 418294 497214 418350
rect 497282 418294 497338 418350
rect 497406 418294 497462 418350
rect 497034 418170 497090 418226
rect 497158 418170 497214 418226
rect 497282 418170 497338 418226
rect 497406 418170 497462 418226
rect 497034 418046 497090 418102
rect 497158 418046 497214 418102
rect 497282 418046 497338 418102
rect 497406 418046 497462 418102
rect 497034 417922 497090 417978
rect 497158 417922 497214 417978
rect 497282 417922 497338 417978
rect 497406 417922 497462 417978
rect 496412 407042 496468 407098
rect 470034 406294 470090 406350
rect 470158 406294 470214 406350
rect 470282 406294 470338 406350
rect 470406 406294 470462 406350
rect 470034 406170 470090 406226
rect 470158 406170 470214 406226
rect 470282 406170 470338 406226
rect 470406 406170 470462 406226
rect 470034 406046 470090 406102
rect 470158 406046 470214 406102
rect 470282 406046 470338 406102
rect 470406 406046 470462 406102
rect 470034 405922 470090 405978
rect 470158 405922 470214 405978
rect 470282 405922 470338 405978
rect 470406 405922 470462 405978
rect 490588 395522 490644 395578
rect 497034 400294 497090 400350
rect 497158 400294 497214 400350
rect 497282 400294 497338 400350
rect 497406 400294 497462 400350
rect 497034 400170 497090 400226
rect 497158 400170 497214 400226
rect 497282 400170 497338 400226
rect 497406 400170 497462 400226
rect 497034 400046 497090 400102
rect 497158 400046 497214 400102
rect 497282 400046 497338 400102
rect 497406 400046 497462 400102
rect 497034 399922 497090 399978
rect 497158 399922 497214 399978
rect 497282 399922 497338 399978
rect 497406 399922 497462 399978
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 500754 568294 500810 568350
rect 500878 568294 500934 568350
rect 501002 568294 501058 568350
rect 501126 568294 501182 568350
rect 500754 568170 500810 568226
rect 500878 568170 500934 568226
rect 501002 568170 501058 568226
rect 501126 568170 501182 568226
rect 500754 568046 500810 568102
rect 500878 568046 500934 568102
rect 501002 568046 501058 568102
rect 501126 568046 501182 568102
rect 500754 567922 500810 567978
rect 500878 567922 500934 567978
rect 501002 567922 501058 567978
rect 501126 567922 501182 567978
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 501718 562294 501774 562350
rect 501842 562294 501898 562350
rect 501718 562170 501774 562226
rect 501842 562170 501898 562226
rect 501718 562046 501774 562102
rect 501842 562046 501898 562102
rect 501718 561922 501774 561978
rect 501842 561922 501898 561978
rect 527754 562294 527810 562350
rect 527878 562294 527934 562350
rect 528002 562294 528058 562350
rect 528126 562294 528182 562350
rect 527754 562170 527810 562226
rect 527878 562170 527934 562226
rect 528002 562170 528058 562226
rect 528126 562170 528182 562226
rect 527754 562046 527810 562102
rect 527878 562046 527934 562102
rect 528002 562046 528058 562102
rect 528126 562046 528182 562102
rect 527754 561922 527810 561978
rect 527878 561922 527934 561978
rect 528002 561922 528058 561978
rect 528126 561922 528182 561978
rect 500754 550294 500810 550350
rect 500878 550294 500934 550350
rect 501002 550294 501058 550350
rect 501126 550294 501182 550350
rect 500754 550170 500810 550226
rect 500878 550170 500934 550226
rect 501002 550170 501058 550226
rect 501126 550170 501182 550226
rect 500754 550046 500810 550102
rect 500878 550046 500934 550102
rect 501002 550046 501058 550102
rect 501126 550046 501182 550102
rect 500754 549922 500810 549978
rect 500878 549922 500934 549978
rect 501002 549922 501058 549978
rect 501126 549922 501182 549978
rect 517078 550294 517134 550350
rect 517202 550294 517258 550350
rect 517078 550170 517134 550226
rect 517202 550170 517258 550226
rect 517078 550046 517134 550102
rect 517202 550046 517258 550102
rect 517078 549922 517134 549978
rect 517202 549922 517258 549978
rect 501718 544294 501774 544350
rect 501842 544294 501898 544350
rect 501718 544170 501774 544226
rect 501842 544170 501898 544226
rect 501718 544046 501774 544102
rect 501842 544046 501898 544102
rect 501718 543922 501774 543978
rect 501842 543922 501898 543978
rect 527754 544294 527810 544350
rect 527878 544294 527934 544350
rect 528002 544294 528058 544350
rect 528126 544294 528182 544350
rect 527754 544170 527810 544226
rect 527878 544170 527934 544226
rect 528002 544170 528058 544226
rect 528126 544170 528182 544226
rect 527754 544046 527810 544102
rect 527878 544046 527934 544102
rect 528002 544046 528058 544102
rect 528126 544046 528182 544102
rect 527754 543922 527810 543978
rect 527878 543922 527934 543978
rect 528002 543922 528058 543978
rect 528126 543922 528182 543978
rect 500754 532294 500810 532350
rect 500878 532294 500934 532350
rect 501002 532294 501058 532350
rect 501126 532294 501182 532350
rect 500754 532170 500810 532226
rect 500878 532170 500934 532226
rect 501002 532170 501058 532226
rect 501126 532170 501182 532226
rect 500754 532046 500810 532102
rect 500878 532046 500934 532102
rect 501002 532046 501058 532102
rect 501126 532046 501182 532102
rect 500754 531922 500810 531978
rect 500878 531922 500934 531978
rect 501002 531922 501058 531978
rect 501126 531922 501182 531978
rect 517078 532294 517134 532350
rect 517202 532294 517258 532350
rect 517078 532170 517134 532226
rect 517202 532170 517258 532226
rect 517078 532046 517134 532102
rect 517202 532046 517258 532102
rect 517078 531922 517134 531978
rect 517202 531922 517258 531978
rect 501718 526294 501774 526350
rect 501842 526294 501898 526350
rect 501718 526170 501774 526226
rect 501842 526170 501898 526226
rect 501718 526046 501774 526102
rect 501842 526046 501898 526102
rect 501718 525922 501774 525978
rect 501842 525922 501898 525978
rect 527754 526294 527810 526350
rect 527878 526294 527934 526350
rect 528002 526294 528058 526350
rect 528126 526294 528182 526350
rect 527754 526170 527810 526226
rect 527878 526170 527934 526226
rect 528002 526170 528058 526226
rect 528126 526170 528182 526226
rect 527754 526046 527810 526102
rect 527878 526046 527934 526102
rect 528002 526046 528058 526102
rect 528126 526046 528182 526102
rect 527754 525922 527810 525978
rect 527878 525922 527934 525978
rect 528002 525922 528058 525978
rect 528126 525922 528182 525978
rect 500754 514294 500810 514350
rect 500878 514294 500934 514350
rect 501002 514294 501058 514350
rect 501126 514294 501182 514350
rect 500754 514170 500810 514226
rect 500878 514170 500934 514226
rect 501002 514170 501058 514226
rect 501126 514170 501182 514226
rect 500754 514046 500810 514102
rect 500878 514046 500934 514102
rect 501002 514046 501058 514102
rect 501126 514046 501182 514102
rect 500754 513922 500810 513978
rect 500878 513922 500934 513978
rect 501002 513922 501058 513978
rect 501126 513922 501182 513978
rect 517078 514294 517134 514350
rect 517202 514294 517258 514350
rect 517078 514170 517134 514226
rect 517202 514170 517258 514226
rect 517078 514046 517134 514102
rect 517202 514046 517258 514102
rect 517078 513922 517134 513978
rect 517202 513922 517258 513978
rect 501718 508294 501774 508350
rect 501842 508294 501898 508350
rect 501718 508170 501774 508226
rect 501842 508170 501898 508226
rect 501718 508046 501774 508102
rect 501842 508046 501898 508102
rect 501718 507922 501774 507978
rect 501842 507922 501898 507978
rect 527754 508294 527810 508350
rect 527878 508294 527934 508350
rect 528002 508294 528058 508350
rect 528126 508294 528182 508350
rect 527754 508170 527810 508226
rect 527878 508170 527934 508226
rect 528002 508170 528058 508226
rect 528126 508170 528182 508226
rect 527754 508046 527810 508102
rect 527878 508046 527934 508102
rect 528002 508046 528058 508102
rect 528126 508046 528182 508102
rect 527754 507922 527810 507978
rect 527878 507922 527934 507978
rect 528002 507922 528058 507978
rect 528126 507922 528182 507978
rect 500754 496294 500810 496350
rect 500878 496294 500934 496350
rect 501002 496294 501058 496350
rect 501126 496294 501182 496350
rect 500754 496170 500810 496226
rect 500878 496170 500934 496226
rect 501002 496170 501058 496226
rect 501126 496170 501182 496226
rect 500754 496046 500810 496102
rect 500878 496046 500934 496102
rect 501002 496046 501058 496102
rect 501126 496046 501182 496102
rect 500754 495922 500810 495978
rect 500878 495922 500934 495978
rect 501002 495922 501058 495978
rect 501126 495922 501182 495978
rect 517078 496294 517134 496350
rect 517202 496294 517258 496350
rect 517078 496170 517134 496226
rect 517202 496170 517258 496226
rect 517078 496046 517134 496102
rect 517202 496046 517258 496102
rect 517078 495922 517134 495978
rect 517202 495922 517258 495978
rect 501718 490294 501774 490350
rect 501842 490294 501898 490350
rect 501718 490170 501774 490226
rect 501842 490170 501898 490226
rect 501718 490046 501774 490102
rect 501842 490046 501898 490102
rect 501718 489922 501774 489978
rect 501842 489922 501898 489978
rect 527754 490294 527810 490350
rect 527878 490294 527934 490350
rect 528002 490294 528058 490350
rect 528126 490294 528182 490350
rect 527754 490170 527810 490226
rect 527878 490170 527934 490226
rect 528002 490170 528058 490226
rect 528126 490170 528182 490226
rect 527754 490046 527810 490102
rect 527878 490046 527934 490102
rect 528002 490046 528058 490102
rect 528126 490046 528182 490102
rect 527754 489922 527810 489978
rect 527878 489922 527934 489978
rect 528002 489922 528058 489978
rect 528126 489922 528182 489978
rect 500754 478294 500810 478350
rect 500878 478294 500934 478350
rect 501002 478294 501058 478350
rect 501126 478294 501182 478350
rect 500754 478170 500810 478226
rect 500878 478170 500934 478226
rect 501002 478170 501058 478226
rect 501126 478170 501182 478226
rect 500754 478046 500810 478102
rect 500878 478046 500934 478102
rect 501002 478046 501058 478102
rect 501126 478046 501182 478102
rect 500754 477922 500810 477978
rect 500878 477922 500934 477978
rect 501002 477922 501058 477978
rect 501126 477922 501182 477978
rect 517078 478294 517134 478350
rect 517202 478294 517258 478350
rect 517078 478170 517134 478226
rect 517202 478170 517258 478226
rect 517078 478046 517134 478102
rect 517202 478046 517258 478102
rect 517078 477922 517134 477978
rect 517202 477922 517258 477978
rect 501718 472294 501774 472350
rect 501842 472294 501898 472350
rect 501718 472170 501774 472226
rect 501842 472170 501898 472226
rect 501718 472046 501774 472102
rect 501842 472046 501898 472102
rect 501718 471922 501774 471978
rect 501842 471922 501898 471978
rect 527754 472294 527810 472350
rect 527878 472294 527934 472350
rect 528002 472294 528058 472350
rect 528126 472294 528182 472350
rect 527754 472170 527810 472226
rect 527878 472170 527934 472226
rect 528002 472170 528058 472226
rect 528126 472170 528182 472226
rect 527754 472046 527810 472102
rect 527878 472046 527934 472102
rect 528002 472046 528058 472102
rect 528126 472046 528182 472102
rect 527754 471922 527810 471978
rect 527878 471922 527934 471978
rect 528002 471922 528058 471978
rect 528126 471922 528182 471978
rect 500754 460294 500810 460350
rect 500878 460294 500934 460350
rect 501002 460294 501058 460350
rect 501126 460294 501182 460350
rect 500754 460170 500810 460226
rect 500878 460170 500934 460226
rect 501002 460170 501058 460226
rect 501126 460170 501182 460226
rect 500754 460046 500810 460102
rect 500878 460046 500934 460102
rect 501002 460046 501058 460102
rect 501126 460046 501182 460102
rect 500754 459922 500810 459978
rect 500878 459922 500934 459978
rect 501002 459922 501058 459978
rect 501126 459922 501182 459978
rect 517078 460294 517134 460350
rect 517202 460294 517258 460350
rect 517078 460170 517134 460226
rect 517202 460170 517258 460226
rect 517078 460046 517134 460102
rect 517202 460046 517258 460102
rect 517078 459922 517134 459978
rect 517202 459922 517258 459978
rect 501718 454294 501774 454350
rect 501842 454294 501898 454350
rect 501718 454170 501774 454226
rect 501842 454170 501898 454226
rect 501718 454046 501774 454102
rect 501842 454046 501898 454102
rect 501718 453922 501774 453978
rect 501842 453922 501898 453978
rect 527754 454294 527810 454350
rect 527878 454294 527934 454350
rect 528002 454294 528058 454350
rect 528126 454294 528182 454350
rect 527754 454170 527810 454226
rect 527878 454170 527934 454226
rect 528002 454170 528058 454226
rect 528126 454170 528182 454226
rect 527754 454046 527810 454102
rect 527878 454046 527934 454102
rect 528002 454046 528058 454102
rect 528126 454046 528182 454102
rect 527754 453922 527810 453978
rect 527878 453922 527934 453978
rect 528002 453922 528058 453978
rect 528126 453922 528182 453978
rect 500754 442294 500810 442350
rect 500878 442294 500934 442350
rect 501002 442294 501058 442350
rect 501126 442294 501182 442350
rect 500754 442170 500810 442226
rect 500878 442170 500934 442226
rect 501002 442170 501058 442226
rect 501126 442170 501182 442226
rect 500754 442046 500810 442102
rect 500878 442046 500934 442102
rect 501002 442046 501058 442102
rect 501126 442046 501182 442102
rect 500754 441922 500810 441978
rect 500878 441922 500934 441978
rect 501002 441922 501058 441978
rect 501126 441922 501182 441978
rect 517078 442294 517134 442350
rect 517202 442294 517258 442350
rect 517078 442170 517134 442226
rect 517202 442170 517258 442226
rect 517078 442046 517134 442102
rect 517202 442046 517258 442102
rect 517078 441922 517134 441978
rect 517202 441922 517258 441978
rect 501718 436294 501774 436350
rect 501842 436294 501898 436350
rect 501718 436170 501774 436226
rect 501842 436170 501898 436226
rect 501718 436046 501774 436102
rect 501842 436046 501898 436102
rect 501718 435922 501774 435978
rect 501842 435922 501898 435978
rect 527754 436294 527810 436350
rect 527878 436294 527934 436350
rect 528002 436294 528058 436350
rect 528126 436294 528182 436350
rect 527754 436170 527810 436226
rect 527878 436170 527934 436226
rect 528002 436170 528058 436226
rect 528126 436170 528182 436226
rect 527754 436046 527810 436102
rect 527878 436046 527934 436102
rect 528002 436046 528058 436102
rect 528126 436046 528182 436102
rect 527754 435922 527810 435978
rect 527878 435922 527934 435978
rect 528002 435922 528058 435978
rect 528126 435922 528182 435978
rect 500754 424294 500810 424350
rect 500878 424294 500934 424350
rect 501002 424294 501058 424350
rect 501126 424294 501182 424350
rect 500754 424170 500810 424226
rect 500878 424170 500934 424226
rect 501002 424170 501058 424226
rect 501126 424170 501182 424226
rect 500754 424046 500810 424102
rect 500878 424046 500934 424102
rect 501002 424046 501058 424102
rect 501126 424046 501182 424102
rect 500754 423922 500810 423978
rect 500878 423922 500934 423978
rect 501002 423922 501058 423978
rect 501126 423922 501182 423978
rect 517078 424294 517134 424350
rect 517202 424294 517258 424350
rect 517078 424170 517134 424226
rect 517202 424170 517258 424226
rect 517078 424046 517134 424102
rect 517202 424046 517258 424102
rect 517078 423922 517134 423978
rect 517202 423922 517258 423978
rect 501718 418294 501774 418350
rect 501842 418294 501898 418350
rect 501718 418170 501774 418226
rect 501842 418170 501898 418226
rect 501718 418046 501774 418102
rect 501842 418046 501898 418102
rect 501718 417922 501774 417978
rect 501842 417922 501898 417978
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 531474 568294 531530 568350
rect 531598 568294 531654 568350
rect 531722 568294 531778 568350
rect 531846 568294 531902 568350
rect 531474 568170 531530 568226
rect 531598 568170 531654 568226
rect 531722 568170 531778 568226
rect 531846 568170 531902 568226
rect 531474 568046 531530 568102
rect 531598 568046 531654 568102
rect 531722 568046 531778 568102
rect 531846 568046 531902 568102
rect 531474 567922 531530 567978
rect 531598 567922 531654 567978
rect 531722 567922 531778 567978
rect 531846 567922 531902 567978
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 531474 550294 531530 550350
rect 531598 550294 531654 550350
rect 531722 550294 531778 550350
rect 531846 550294 531902 550350
rect 531474 550170 531530 550226
rect 531598 550170 531654 550226
rect 531722 550170 531778 550226
rect 531846 550170 531902 550226
rect 531474 550046 531530 550102
rect 531598 550046 531654 550102
rect 531722 550046 531778 550102
rect 531846 550046 531902 550102
rect 531474 549922 531530 549978
rect 531598 549922 531654 549978
rect 531722 549922 531778 549978
rect 531846 549922 531902 549978
rect 531474 532294 531530 532350
rect 531598 532294 531654 532350
rect 531722 532294 531778 532350
rect 531846 532294 531902 532350
rect 531474 532170 531530 532226
rect 531598 532170 531654 532226
rect 531722 532170 531778 532226
rect 531846 532170 531902 532226
rect 531474 532046 531530 532102
rect 531598 532046 531654 532102
rect 531722 532046 531778 532102
rect 531846 532046 531902 532102
rect 531474 531922 531530 531978
rect 531598 531922 531654 531978
rect 531722 531922 531778 531978
rect 531846 531922 531902 531978
rect 531474 514294 531530 514350
rect 531598 514294 531654 514350
rect 531722 514294 531778 514350
rect 531846 514294 531902 514350
rect 531474 514170 531530 514226
rect 531598 514170 531654 514226
rect 531722 514170 531778 514226
rect 531846 514170 531902 514226
rect 531474 514046 531530 514102
rect 531598 514046 531654 514102
rect 531722 514046 531778 514102
rect 531846 514046 531902 514102
rect 531474 513922 531530 513978
rect 531598 513922 531654 513978
rect 531722 513922 531778 513978
rect 531846 513922 531902 513978
rect 531474 496294 531530 496350
rect 531598 496294 531654 496350
rect 531722 496294 531778 496350
rect 531846 496294 531902 496350
rect 531474 496170 531530 496226
rect 531598 496170 531654 496226
rect 531722 496170 531778 496226
rect 531846 496170 531902 496226
rect 531474 496046 531530 496102
rect 531598 496046 531654 496102
rect 531722 496046 531778 496102
rect 531846 496046 531902 496102
rect 531474 495922 531530 495978
rect 531598 495922 531654 495978
rect 531722 495922 531778 495978
rect 531846 495922 531902 495978
rect 531474 478294 531530 478350
rect 531598 478294 531654 478350
rect 531722 478294 531778 478350
rect 531846 478294 531902 478350
rect 531474 478170 531530 478226
rect 531598 478170 531654 478226
rect 531722 478170 531778 478226
rect 531846 478170 531902 478226
rect 531474 478046 531530 478102
rect 531598 478046 531654 478102
rect 531722 478046 531778 478102
rect 531846 478046 531902 478102
rect 531474 477922 531530 477978
rect 531598 477922 531654 477978
rect 531722 477922 531778 477978
rect 531846 477922 531902 477978
rect 531474 460294 531530 460350
rect 531598 460294 531654 460350
rect 531722 460294 531778 460350
rect 531846 460294 531902 460350
rect 531474 460170 531530 460226
rect 531598 460170 531654 460226
rect 531722 460170 531778 460226
rect 531846 460170 531902 460226
rect 531474 460046 531530 460102
rect 531598 460046 531654 460102
rect 531722 460046 531778 460102
rect 531846 460046 531902 460102
rect 531474 459922 531530 459978
rect 531598 459922 531654 459978
rect 531722 459922 531778 459978
rect 531846 459922 531902 459978
rect 531474 442294 531530 442350
rect 531598 442294 531654 442350
rect 531722 442294 531778 442350
rect 531846 442294 531902 442350
rect 531474 442170 531530 442226
rect 531598 442170 531654 442226
rect 531722 442170 531778 442226
rect 531846 442170 531902 442226
rect 531474 442046 531530 442102
rect 531598 442046 531654 442102
rect 531722 442046 531778 442102
rect 531846 442046 531902 442102
rect 531474 441922 531530 441978
rect 531598 441922 531654 441978
rect 531722 441922 531778 441978
rect 531846 441922 531902 441978
rect 529228 428652 529284 428698
rect 529228 428642 529284 428652
rect 527754 418294 527810 418350
rect 527878 418294 527934 418350
rect 528002 418294 528058 418350
rect 528126 418294 528182 418350
rect 527754 418170 527810 418226
rect 527878 418170 527934 418226
rect 528002 418170 528058 418226
rect 528126 418170 528182 418226
rect 527754 418046 527810 418102
rect 527878 418046 527934 418102
rect 528002 418046 528058 418102
rect 528126 418046 528182 418102
rect 527754 417922 527810 417978
rect 527878 417922 527934 417978
rect 528002 417922 528058 417978
rect 528126 417922 528182 417978
rect 522172 406862 522228 406918
rect 527324 406682 527380 406738
rect 500754 406294 500810 406350
rect 500878 406294 500934 406350
rect 501002 406294 501058 406350
rect 501126 406294 501182 406350
rect 500754 406170 500810 406226
rect 500878 406170 500934 406226
rect 501002 406170 501058 406226
rect 501126 406170 501182 406226
rect 500754 406046 500810 406102
rect 500878 406046 500934 406102
rect 501002 406046 501058 406102
rect 501126 406046 501182 406102
rect 500754 405922 500810 405978
rect 500878 405922 500934 405978
rect 501002 405922 501058 405978
rect 501126 405922 501182 405978
rect 527754 400294 527810 400350
rect 527878 400294 527934 400350
rect 528002 400294 528058 400350
rect 528126 400294 528182 400350
rect 527754 400170 527810 400226
rect 527878 400170 527934 400226
rect 528002 400170 528058 400226
rect 528126 400170 528182 400226
rect 527754 400046 527810 400102
rect 527878 400046 527934 400102
rect 528002 400046 528058 400102
rect 528126 400046 528182 400102
rect 527754 399922 527810 399978
rect 527878 399922 527934 399978
rect 528002 399922 528058 399978
rect 528126 399922 528182 399978
rect 525532 394996 525588 395038
rect 525532 394982 525588 394996
rect 531474 424294 531530 424350
rect 531598 424294 531654 424350
rect 531722 424294 531778 424350
rect 531846 424294 531902 424350
rect 531474 424170 531530 424226
rect 531598 424170 531654 424226
rect 531722 424170 531778 424226
rect 531846 424170 531902 424226
rect 531474 424046 531530 424102
rect 531598 424046 531654 424102
rect 531722 424046 531778 424102
rect 531846 424046 531902 424102
rect 531474 423922 531530 423978
rect 531598 423922 531654 423978
rect 531722 423922 531778 423978
rect 531846 423922 531902 423978
rect 532700 409382 532756 409438
rect 532812 407402 532868 407458
rect 531474 406294 531530 406350
rect 531598 406294 531654 406350
rect 531722 406294 531778 406350
rect 531846 406294 531902 406350
rect 531474 406170 531530 406226
rect 531598 406170 531654 406226
rect 531722 406170 531778 406226
rect 531846 406170 531902 406226
rect 531474 406046 531530 406102
rect 531598 406046 531654 406102
rect 531722 406046 531778 406102
rect 531846 406046 531902 406102
rect 531474 405922 531530 405978
rect 531598 405922 531654 405978
rect 531722 405922 531778 405978
rect 531846 405922 531902 405978
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 532924 405422 532980 405478
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 537628 409202 537684 409258
rect 535948 405602 536004 405658
rect 541772 404342 541828 404398
rect 540092 404162 540148 404218
rect 543452 402722 543508 402778
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 558474 472294 558530 472350
rect 558598 472294 558654 472350
rect 558722 472294 558778 472350
rect 558846 472294 558902 472350
rect 558474 472170 558530 472226
rect 558598 472170 558654 472226
rect 558722 472170 558778 472226
rect 558846 472170 558902 472226
rect 558474 472046 558530 472102
rect 558598 472046 558654 472102
rect 558722 472046 558778 472102
rect 558846 472046 558902 472102
rect 558474 471922 558530 471978
rect 558598 471922 558654 471978
rect 558722 471922 558778 471978
rect 558846 471922 558902 471978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 534268 398942 534324 398998
rect 558474 400294 558530 400350
rect 558598 400294 558654 400350
rect 558722 400294 558778 400350
rect 558846 400294 558902 400350
rect 558474 400170 558530 400226
rect 558598 400170 558654 400226
rect 558722 400170 558778 400226
rect 558846 400170 558902 400226
rect 558474 400046 558530 400102
rect 558598 400046 558654 400102
rect 558722 400046 558778 400102
rect 558846 400046 558902 400102
rect 558474 399922 558530 399978
rect 558598 399922 558654 399978
rect 558722 399922 558778 399978
rect 558846 399922 558902 399978
rect 546252 397322 546308 397378
rect 553196 396782 553252 396838
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 584668 409742 584724 409798
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 574028 397142 574084 397198
rect 580972 396962 581028 397018
rect 567084 396602 567140 396658
rect 364476 392642 364532 392698
rect 374878 388294 374934 388350
rect 375002 388294 375058 388350
rect 374878 388170 374934 388226
rect 375002 388170 375058 388226
rect 374878 388046 374934 388102
rect 375002 388046 375058 388102
rect 374878 387922 374934 387978
rect 375002 387922 375058 387978
rect 405598 388294 405654 388350
rect 405722 388294 405778 388350
rect 405598 388170 405654 388226
rect 405722 388170 405778 388226
rect 405598 388046 405654 388102
rect 405722 388046 405778 388102
rect 405598 387922 405654 387978
rect 405722 387922 405778 387978
rect 436318 388294 436374 388350
rect 436442 388294 436498 388350
rect 436318 388170 436374 388226
rect 436442 388170 436498 388226
rect 436318 388046 436374 388102
rect 436442 388046 436498 388102
rect 436318 387922 436374 387978
rect 436442 387922 436498 387978
rect 467038 388294 467094 388350
rect 467162 388294 467218 388350
rect 467038 388170 467094 388226
rect 467162 388170 467218 388226
rect 467038 388046 467094 388102
rect 467162 388046 467218 388102
rect 467038 387922 467094 387978
rect 467162 387922 467218 387978
rect 497758 388294 497814 388350
rect 497882 388294 497938 388350
rect 497758 388170 497814 388226
rect 497882 388170 497938 388226
rect 497758 388046 497814 388102
rect 497882 388046 497938 388102
rect 497758 387922 497814 387978
rect 497882 387922 497938 387978
rect 528478 388294 528534 388350
rect 528602 388294 528658 388350
rect 528478 388170 528534 388226
rect 528602 388170 528658 388226
rect 528478 388046 528534 388102
rect 528602 388046 528658 388102
rect 528478 387922 528534 387978
rect 528602 387922 528658 387978
rect 559198 388294 559254 388350
rect 559322 388294 559378 388350
rect 559198 388170 559254 388226
rect 559322 388170 559378 388226
rect 559198 388046 559254 388102
rect 559322 388046 559378 388102
rect 559198 387922 559254 387978
rect 559322 387922 559378 387978
rect 359518 382294 359574 382350
rect 359642 382294 359698 382350
rect 359518 382170 359574 382226
rect 359642 382170 359698 382226
rect 359518 382046 359574 382102
rect 359642 382046 359698 382102
rect 359518 381922 359574 381978
rect 359642 381922 359698 381978
rect 390238 382294 390294 382350
rect 390362 382294 390418 382350
rect 390238 382170 390294 382226
rect 390362 382170 390418 382226
rect 390238 382046 390294 382102
rect 390362 382046 390418 382102
rect 390238 381922 390294 381978
rect 390362 381922 390418 381978
rect 420958 382294 421014 382350
rect 421082 382294 421138 382350
rect 420958 382170 421014 382226
rect 421082 382170 421138 382226
rect 420958 382046 421014 382102
rect 421082 382046 421138 382102
rect 420958 381922 421014 381978
rect 421082 381922 421138 381978
rect 451678 382294 451734 382350
rect 451802 382294 451858 382350
rect 451678 382170 451734 382226
rect 451802 382170 451858 382226
rect 451678 382046 451734 382102
rect 451802 382046 451858 382102
rect 451678 381922 451734 381978
rect 451802 381922 451858 381978
rect 482398 382294 482454 382350
rect 482522 382294 482578 382350
rect 482398 382170 482454 382226
rect 482522 382170 482578 382226
rect 482398 382046 482454 382102
rect 482522 382046 482578 382102
rect 482398 381922 482454 381978
rect 482522 381922 482578 381978
rect 513118 382294 513174 382350
rect 513242 382294 513298 382350
rect 513118 382170 513174 382226
rect 513242 382170 513298 382226
rect 513118 382046 513174 382102
rect 513242 382046 513298 382102
rect 513118 381922 513174 381978
rect 513242 381922 513298 381978
rect 543838 382294 543894 382350
rect 543962 382294 544018 382350
rect 543838 382170 543894 382226
rect 543962 382170 544018 382226
rect 543838 382046 543894 382102
rect 543962 382046 544018 382102
rect 543838 381922 543894 381978
rect 543962 381922 544018 381978
rect 574558 382294 574614 382350
rect 574682 382294 574738 382350
rect 574558 382170 574614 382226
rect 574682 382170 574738 382226
rect 574558 382046 574614 382102
rect 574682 382046 574738 382102
rect 574558 381922 574614 381978
rect 574682 381922 574738 381978
rect 374878 370294 374934 370350
rect 375002 370294 375058 370350
rect 374878 370170 374934 370226
rect 375002 370170 375058 370226
rect 374878 370046 374934 370102
rect 375002 370046 375058 370102
rect 374878 369922 374934 369978
rect 375002 369922 375058 369978
rect 405598 370294 405654 370350
rect 405722 370294 405778 370350
rect 405598 370170 405654 370226
rect 405722 370170 405778 370226
rect 405598 370046 405654 370102
rect 405722 370046 405778 370102
rect 405598 369922 405654 369978
rect 405722 369922 405778 369978
rect 436318 370294 436374 370350
rect 436442 370294 436498 370350
rect 436318 370170 436374 370226
rect 436442 370170 436498 370226
rect 436318 370046 436374 370102
rect 436442 370046 436498 370102
rect 436318 369922 436374 369978
rect 436442 369922 436498 369978
rect 467038 370294 467094 370350
rect 467162 370294 467218 370350
rect 467038 370170 467094 370226
rect 467162 370170 467218 370226
rect 467038 370046 467094 370102
rect 467162 370046 467218 370102
rect 467038 369922 467094 369978
rect 467162 369922 467218 369978
rect 497758 370294 497814 370350
rect 497882 370294 497938 370350
rect 497758 370170 497814 370226
rect 497882 370170 497938 370226
rect 497758 370046 497814 370102
rect 497882 370046 497938 370102
rect 497758 369922 497814 369978
rect 497882 369922 497938 369978
rect 528478 370294 528534 370350
rect 528602 370294 528658 370350
rect 528478 370170 528534 370226
rect 528602 370170 528658 370226
rect 528478 370046 528534 370102
rect 528602 370046 528658 370102
rect 528478 369922 528534 369978
rect 528602 369922 528658 369978
rect 559198 370294 559254 370350
rect 559322 370294 559378 370350
rect 559198 370170 559254 370226
rect 559322 370170 559378 370226
rect 559198 370046 559254 370102
rect 559322 370046 559378 370102
rect 559198 369922 559254 369978
rect 559322 369922 559378 369978
rect 359518 364294 359574 364350
rect 359642 364294 359698 364350
rect 359518 364170 359574 364226
rect 359642 364170 359698 364226
rect 359518 364046 359574 364102
rect 359642 364046 359698 364102
rect 359518 363922 359574 363978
rect 359642 363922 359698 363978
rect 390238 364294 390294 364350
rect 390362 364294 390418 364350
rect 390238 364170 390294 364226
rect 390362 364170 390418 364226
rect 390238 364046 390294 364102
rect 390362 364046 390418 364102
rect 390238 363922 390294 363978
rect 390362 363922 390418 363978
rect 420958 364294 421014 364350
rect 421082 364294 421138 364350
rect 420958 364170 421014 364226
rect 421082 364170 421138 364226
rect 420958 364046 421014 364102
rect 421082 364046 421138 364102
rect 420958 363922 421014 363978
rect 421082 363922 421138 363978
rect 451678 364294 451734 364350
rect 451802 364294 451858 364350
rect 451678 364170 451734 364226
rect 451802 364170 451858 364226
rect 451678 364046 451734 364102
rect 451802 364046 451858 364102
rect 451678 363922 451734 363978
rect 451802 363922 451858 363978
rect 482398 364294 482454 364350
rect 482522 364294 482578 364350
rect 482398 364170 482454 364226
rect 482522 364170 482578 364226
rect 482398 364046 482454 364102
rect 482522 364046 482578 364102
rect 482398 363922 482454 363978
rect 482522 363922 482578 363978
rect 513118 364294 513174 364350
rect 513242 364294 513298 364350
rect 513118 364170 513174 364226
rect 513242 364170 513298 364226
rect 513118 364046 513174 364102
rect 513242 364046 513298 364102
rect 513118 363922 513174 363978
rect 513242 363922 513298 363978
rect 543838 364294 543894 364350
rect 543962 364294 544018 364350
rect 543838 364170 543894 364226
rect 543962 364170 544018 364226
rect 543838 364046 543894 364102
rect 543962 364046 544018 364102
rect 543838 363922 543894 363978
rect 543962 363922 544018 363978
rect 574558 364294 574614 364350
rect 574682 364294 574738 364350
rect 574558 364170 574614 364226
rect 574682 364170 574738 364226
rect 574558 364046 574614 364102
rect 574682 364046 574738 364102
rect 574558 363922 574614 363978
rect 574682 363922 574738 363978
rect 374878 352294 374934 352350
rect 375002 352294 375058 352350
rect 374878 352170 374934 352226
rect 375002 352170 375058 352226
rect 374878 352046 374934 352102
rect 375002 352046 375058 352102
rect 374878 351922 374934 351978
rect 375002 351922 375058 351978
rect 405598 352294 405654 352350
rect 405722 352294 405778 352350
rect 405598 352170 405654 352226
rect 405722 352170 405778 352226
rect 405598 352046 405654 352102
rect 405722 352046 405778 352102
rect 405598 351922 405654 351978
rect 405722 351922 405778 351978
rect 436318 352294 436374 352350
rect 436442 352294 436498 352350
rect 436318 352170 436374 352226
rect 436442 352170 436498 352226
rect 436318 352046 436374 352102
rect 436442 352046 436498 352102
rect 436318 351922 436374 351978
rect 436442 351922 436498 351978
rect 467038 352294 467094 352350
rect 467162 352294 467218 352350
rect 467038 352170 467094 352226
rect 467162 352170 467218 352226
rect 467038 352046 467094 352102
rect 467162 352046 467218 352102
rect 467038 351922 467094 351978
rect 467162 351922 467218 351978
rect 497758 352294 497814 352350
rect 497882 352294 497938 352350
rect 497758 352170 497814 352226
rect 497882 352170 497938 352226
rect 497758 352046 497814 352102
rect 497882 352046 497938 352102
rect 497758 351922 497814 351978
rect 497882 351922 497938 351978
rect 528478 352294 528534 352350
rect 528602 352294 528658 352350
rect 528478 352170 528534 352226
rect 528602 352170 528658 352226
rect 528478 352046 528534 352102
rect 528602 352046 528658 352102
rect 528478 351922 528534 351978
rect 528602 351922 528658 351978
rect 559198 352294 559254 352350
rect 559322 352294 559378 352350
rect 559198 352170 559254 352226
rect 559322 352170 559378 352226
rect 559198 352046 559254 352102
rect 559322 352046 559378 352102
rect 559198 351922 559254 351978
rect 559322 351922 559378 351978
rect 359518 346294 359574 346350
rect 359642 346294 359698 346350
rect 359518 346170 359574 346226
rect 359642 346170 359698 346226
rect 359518 346046 359574 346102
rect 359642 346046 359698 346102
rect 359518 345922 359574 345978
rect 359642 345922 359698 345978
rect 390238 346294 390294 346350
rect 390362 346294 390418 346350
rect 390238 346170 390294 346226
rect 390362 346170 390418 346226
rect 390238 346046 390294 346102
rect 390362 346046 390418 346102
rect 390238 345922 390294 345978
rect 390362 345922 390418 345978
rect 420958 346294 421014 346350
rect 421082 346294 421138 346350
rect 420958 346170 421014 346226
rect 421082 346170 421138 346226
rect 420958 346046 421014 346102
rect 421082 346046 421138 346102
rect 420958 345922 421014 345978
rect 421082 345922 421138 345978
rect 451678 346294 451734 346350
rect 451802 346294 451858 346350
rect 451678 346170 451734 346226
rect 451802 346170 451858 346226
rect 451678 346046 451734 346102
rect 451802 346046 451858 346102
rect 451678 345922 451734 345978
rect 451802 345922 451858 345978
rect 482398 346294 482454 346350
rect 482522 346294 482578 346350
rect 482398 346170 482454 346226
rect 482522 346170 482578 346226
rect 482398 346046 482454 346102
rect 482522 346046 482578 346102
rect 482398 345922 482454 345978
rect 482522 345922 482578 345978
rect 513118 346294 513174 346350
rect 513242 346294 513298 346350
rect 513118 346170 513174 346226
rect 513242 346170 513298 346226
rect 513118 346046 513174 346102
rect 513242 346046 513298 346102
rect 513118 345922 513174 345978
rect 513242 345922 513298 345978
rect 543838 346294 543894 346350
rect 543962 346294 544018 346350
rect 543838 346170 543894 346226
rect 543962 346170 544018 346226
rect 543838 346046 543894 346102
rect 543962 346046 544018 346102
rect 543838 345922 543894 345978
rect 543962 345922 544018 345978
rect 574558 346294 574614 346350
rect 574682 346294 574738 346350
rect 574558 346170 574614 346226
rect 574682 346170 574738 346226
rect 574558 346046 574614 346102
rect 574682 346046 574738 346102
rect 574558 345922 574614 345978
rect 574682 345922 574738 345978
rect 374878 334294 374934 334350
rect 375002 334294 375058 334350
rect 374878 334170 374934 334226
rect 375002 334170 375058 334226
rect 374878 334046 374934 334102
rect 375002 334046 375058 334102
rect 374878 333922 374934 333978
rect 375002 333922 375058 333978
rect 405598 334294 405654 334350
rect 405722 334294 405778 334350
rect 405598 334170 405654 334226
rect 405722 334170 405778 334226
rect 405598 334046 405654 334102
rect 405722 334046 405778 334102
rect 405598 333922 405654 333978
rect 405722 333922 405778 333978
rect 436318 334294 436374 334350
rect 436442 334294 436498 334350
rect 436318 334170 436374 334226
rect 436442 334170 436498 334226
rect 436318 334046 436374 334102
rect 436442 334046 436498 334102
rect 436318 333922 436374 333978
rect 436442 333922 436498 333978
rect 467038 334294 467094 334350
rect 467162 334294 467218 334350
rect 467038 334170 467094 334226
rect 467162 334170 467218 334226
rect 467038 334046 467094 334102
rect 467162 334046 467218 334102
rect 467038 333922 467094 333978
rect 467162 333922 467218 333978
rect 497758 334294 497814 334350
rect 497882 334294 497938 334350
rect 497758 334170 497814 334226
rect 497882 334170 497938 334226
rect 497758 334046 497814 334102
rect 497882 334046 497938 334102
rect 497758 333922 497814 333978
rect 497882 333922 497938 333978
rect 528478 334294 528534 334350
rect 528602 334294 528658 334350
rect 528478 334170 528534 334226
rect 528602 334170 528658 334226
rect 528478 334046 528534 334102
rect 528602 334046 528658 334102
rect 528478 333922 528534 333978
rect 528602 333922 528658 333978
rect 559198 334294 559254 334350
rect 559322 334294 559378 334350
rect 559198 334170 559254 334226
rect 559322 334170 559378 334226
rect 559198 334046 559254 334102
rect 559322 334046 559378 334102
rect 559198 333922 559254 333978
rect 559322 333922 559378 333978
rect 359518 328294 359574 328350
rect 359642 328294 359698 328350
rect 359518 328170 359574 328226
rect 359642 328170 359698 328226
rect 359518 328046 359574 328102
rect 359642 328046 359698 328102
rect 359518 327922 359574 327978
rect 359642 327922 359698 327978
rect 390238 328294 390294 328350
rect 390362 328294 390418 328350
rect 390238 328170 390294 328226
rect 390362 328170 390418 328226
rect 390238 328046 390294 328102
rect 390362 328046 390418 328102
rect 390238 327922 390294 327978
rect 390362 327922 390418 327978
rect 420958 328294 421014 328350
rect 421082 328294 421138 328350
rect 420958 328170 421014 328226
rect 421082 328170 421138 328226
rect 420958 328046 421014 328102
rect 421082 328046 421138 328102
rect 420958 327922 421014 327978
rect 421082 327922 421138 327978
rect 451678 328294 451734 328350
rect 451802 328294 451858 328350
rect 451678 328170 451734 328226
rect 451802 328170 451858 328226
rect 451678 328046 451734 328102
rect 451802 328046 451858 328102
rect 451678 327922 451734 327978
rect 451802 327922 451858 327978
rect 482398 328294 482454 328350
rect 482522 328294 482578 328350
rect 482398 328170 482454 328226
rect 482522 328170 482578 328226
rect 482398 328046 482454 328102
rect 482522 328046 482578 328102
rect 482398 327922 482454 327978
rect 482522 327922 482578 327978
rect 513118 328294 513174 328350
rect 513242 328294 513298 328350
rect 513118 328170 513174 328226
rect 513242 328170 513298 328226
rect 513118 328046 513174 328102
rect 513242 328046 513298 328102
rect 513118 327922 513174 327978
rect 513242 327922 513298 327978
rect 543838 328294 543894 328350
rect 543962 328294 544018 328350
rect 543838 328170 543894 328226
rect 543962 328170 544018 328226
rect 543838 328046 543894 328102
rect 543962 328046 544018 328102
rect 543838 327922 543894 327978
rect 543962 327922 544018 327978
rect 574558 328294 574614 328350
rect 574682 328294 574738 328350
rect 574558 328170 574614 328226
rect 574682 328170 574738 328226
rect 574558 328046 574614 328102
rect 574682 328046 574738 328102
rect 574558 327922 574614 327978
rect 574682 327922 574738 327978
rect 374878 316294 374934 316350
rect 375002 316294 375058 316350
rect 374878 316170 374934 316226
rect 375002 316170 375058 316226
rect 374878 316046 374934 316102
rect 375002 316046 375058 316102
rect 374878 315922 374934 315978
rect 375002 315922 375058 315978
rect 405598 316294 405654 316350
rect 405722 316294 405778 316350
rect 405598 316170 405654 316226
rect 405722 316170 405778 316226
rect 405598 316046 405654 316102
rect 405722 316046 405778 316102
rect 405598 315922 405654 315978
rect 405722 315922 405778 315978
rect 436318 316294 436374 316350
rect 436442 316294 436498 316350
rect 436318 316170 436374 316226
rect 436442 316170 436498 316226
rect 436318 316046 436374 316102
rect 436442 316046 436498 316102
rect 436318 315922 436374 315978
rect 436442 315922 436498 315978
rect 467038 316294 467094 316350
rect 467162 316294 467218 316350
rect 467038 316170 467094 316226
rect 467162 316170 467218 316226
rect 467038 316046 467094 316102
rect 467162 316046 467218 316102
rect 467038 315922 467094 315978
rect 467162 315922 467218 315978
rect 497758 316294 497814 316350
rect 497882 316294 497938 316350
rect 497758 316170 497814 316226
rect 497882 316170 497938 316226
rect 497758 316046 497814 316102
rect 497882 316046 497938 316102
rect 497758 315922 497814 315978
rect 497882 315922 497938 315978
rect 528478 316294 528534 316350
rect 528602 316294 528658 316350
rect 528478 316170 528534 316226
rect 528602 316170 528658 316226
rect 528478 316046 528534 316102
rect 528602 316046 528658 316102
rect 528478 315922 528534 315978
rect 528602 315922 528658 315978
rect 559198 316294 559254 316350
rect 559322 316294 559378 316350
rect 559198 316170 559254 316226
rect 559322 316170 559378 316226
rect 559198 316046 559254 316102
rect 559322 316046 559378 316102
rect 559198 315922 559254 315978
rect 559322 315922 559378 315978
rect 359518 310294 359574 310350
rect 359642 310294 359698 310350
rect 359518 310170 359574 310226
rect 359642 310170 359698 310226
rect 359518 310046 359574 310102
rect 359642 310046 359698 310102
rect 359518 309922 359574 309978
rect 359642 309922 359698 309978
rect 390238 310294 390294 310350
rect 390362 310294 390418 310350
rect 390238 310170 390294 310226
rect 390362 310170 390418 310226
rect 390238 310046 390294 310102
rect 390362 310046 390418 310102
rect 390238 309922 390294 309978
rect 390362 309922 390418 309978
rect 420958 310294 421014 310350
rect 421082 310294 421138 310350
rect 420958 310170 421014 310226
rect 421082 310170 421138 310226
rect 420958 310046 421014 310102
rect 421082 310046 421138 310102
rect 420958 309922 421014 309978
rect 421082 309922 421138 309978
rect 451678 310294 451734 310350
rect 451802 310294 451858 310350
rect 451678 310170 451734 310226
rect 451802 310170 451858 310226
rect 451678 310046 451734 310102
rect 451802 310046 451858 310102
rect 451678 309922 451734 309978
rect 451802 309922 451858 309978
rect 482398 310294 482454 310350
rect 482522 310294 482578 310350
rect 482398 310170 482454 310226
rect 482522 310170 482578 310226
rect 482398 310046 482454 310102
rect 482522 310046 482578 310102
rect 482398 309922 482454 309978
rect 482522 309922 482578 309978
rect 513118 310294 513174 310350
rect 513242 310294 513298 310350
rect 513118 310170 513174 310226
rect 513242 310170 513298 310226
rect 513118 310046 513174 310102
rect 513242 310046 513298 310102
rect 513118 309922 513174 309978
rect 513242 309922 513298 309978
rect 543838 310294 543894 310350
rect 543962 310294 544018 310350
rect 543838 310170 543894 310226
rect 543962 310170 544018 310226
rect 543838 310046 543894 310102
rect 543962 310046 544018 310102
rect 543838 309922 543894 309978
rect 543962 309922 544018 309978
rect 574558 310294 574614 310350
rect 574682 310294 574738 310350
rect 574558 310170 574614 310226
rect 574682 310170 574738 310226
rect 574558 310046 574614 310102
rect 574682 310046 574738 310102
rect 574558 309922 574614 309978
rect 574682 309922 574738 309978
rect 374878 298294 374934 298350
rect 375002 298294 375058 298350
rect 374878 298170 374934 298226
rect 375002 298170 375058 298226
rect 374878 298046 374934 298102
rect 375002 298046 375058 298102
rect 374878 297922 374934 297978
rect 375002 297922 375058 297978
rect 405598 298294 405654 298350
rect 405722 298294 405778 298350
rect 405598 298170 405654 298226
rect 405722 298170 405778 298226
rect 405598 298046 405654 298102
rect 405722 298046 405778 298102
rect 405598 297922 405654 297978
rect 405722 297922 405778 297978
rect 436318 298294 436374 298350
rect 436442 298294 436498 298350
rect 436318 298170 436374 298226
rect 436442 298170 436498 298226
rect 436318 298046 436374 298102
rect 436442 298046 436498 298102
rect 436318 297922 436374 297978
rect 436442 297922 436498 297978
rect 467038 298294 467094 298350
rect 467162 298294 467218 298350
rect 467038 298170 467094 298226
rect 467162 298170 467218 298226
rect 467038 298046 467094 298102
rect 467162 298046 467218 298102
rect 467038 297922 467094 297978
rect 467162 297922 467218 297978
rect 497758 298294 497814 298350
rect 497882 298294 497938 298350
rect 497758 298170 497814 298226
rect 497882 298170 497938 298226
rect 497758 298046 497814 298102
rect 497882 298046 497938 298102
rect 497758 297922 497814 297978
rect 497882 297922 497938 297978
rect 528478 298294 528534 298350
rect 528602 298294 528658 298350
rect 528478 298170 528534 298226
rect 528602 298170 528658 298226
rect 528478 298046 528534 298102
rect 528602 298046 528658 298102
rect 528478 297922 528534 297978
rect 528602 297922 528658 297978
rect 559198 298294 559254 298350
rect 559322 298294 559378 298350
rect 559198 298170 559254 298226
rect 559322 298170 559378 298226
rect 559198 298046 559254 298102
rect 559322 298046 559378 298102
rect 559198 297922 559254 297978
rect 559322 297922 559378 297978
rect 359518 292294 359574 292350
rect 359642 292294 359698 292350
rect 359518 292170 359574 292226
rect 359642 292170 359698 292226
rect 359518 292046 359574 292102
rect 359642 292046 359698 292102
rect 359518 291922 359574 291978
rect 359642 291922 359698 291978
rect 390238 292294 390294 292350
rect 390362 292294 390418 292350
rect 390238 292170 390294 292226
rect 390362 292170 390418 292226
rect 390238 292046 390294 292102
rect 390362 292046 390418 292102
rect 390238 291922 390294 291978
rect 390362 291922 390418 291978
rect 420958 292294 421014 292350
rect 421082 292294 421138 292350
rect 420958 292170 421014 292226
rect 421082 292170 421138 292226
rect 420958 292046 421014 292102
rect 421082 292046 421138 292102
rect 420958 291922 421014 291978
rect 421082 291922 421138 291978
rect 451678 292294 451734 292350
rect 451802 292294 451858 292350
rect 451678 292170 451734 292226
rect 451802 292170 451858 292226
rect 451678 292046 451734 292102
rect 451802 292046 451858 292102
rect 451678 291922 451734 291978
rect 451802 291922 451858 291978
rect 482398 292294 482454 292350
rect 482522 292294 482578 292350
rect 482398 292170 482454 292226
rect 482522 292170 482578 292226
rect 482398 292046 482454 292102
rect 482522 292046 482578 292102
rect 482398 291922 482454 291978
rect 482522 291922 482578 291978
rect 513118 292294 513174 292350
rect 513242 292294 513298 292350
rect 513118 292170 513174 292226
rect 513242 292170 513298 292226
rect 513118 292046 513174 292102
rect 513242 292046 513298 292102
rect 513118 291922 513174 291978
rect 513242 291922 513298 291978
rect 543838 292294 543894 292350
rect 543962 292294 544018 292350
rect 543838 292170 543894 292226
rect 543962 292170 544018 292226
rect 543838 292046 543894 292102
rect 543962 292046 544018 292102
rect 543838 291922 543894 291978
rect 543962 291922 544018 291978
rect 574558 292294 574614 292350
rect 574682 292294 574738 292350
rect 574558 292170 574614 292226
rect 574682 292170 574738 292226
rect 574558 292046 574614 292102
rect 574682 292046 574738 292102
rect 574558 291922 574614 291978
rect 574682 291922 574738 291978
rect 374878 280294 374934 280350
rect 375002 280294 375058 280350
rect 374878 280170 374934 280226
rect 375002 280170 375058 280226
rect 374878 280046 374934 280102
rect 375002 280046 375058 280102
rect 374878 279922 374934 279978
rect 375002 279922 375058 279978
rect 405598 280294 405654 280350
rect 405722 280294 405778 280350
rect 405598 280170 405654 280226
rect 405722 280170 405778 280226
rect 405598 280046 405654 280102
rect 405722 280046 405778 280102
rect 405598 279922 405654 279978
rect 405722 279922 405778 279978
rect 436318 280294 436374 280350
rect 436442 280294 436498 280350
rect 436318 280170 436374 280226
rect 436442 280170 436498 280226
rect 436318 280046 436374 280102
rect 436442 280046 436498 280102
rect 436318 279922 436374 279978
rect 436442 279922 436498 279978
rect 467038 280294 467094 280350
rect 467162 280294 467218 280350
rect 467038 280170 467094 280226
rect 467162 280170 467218 280226
rect 467038 280046 467094 280102
rect 467162 280046 467218 280102
rect 467038 279922 467094 279978
rect 467162 279922 467218 279978
rect 497758 280294 497814 280350
rect 497882 280294 497938 280350
rect 497758 280170 497814 280226
rect 497882 280170 497938 280226
rect 497758 280046 497814 280102
rect 497882 280046 497938 280102
rect 497758 279922 497814 279978
rect 497882 279922 497938 279978
rect 528478 280294 528534 280350
rect 528602 280294 528658 280350
rect 528478 280170 528534 280226
rect 528602 280170 528658 280226
rect 528478 280046 528534 280102
rect 528602 280046 528658 280102
rect 528478 279922 528534 279978
rect 528602 279922 528658 279978
rect 559198 280294 559254 280350
rect 559322 280294 559378 280350
rect 559198 280170 559254 280226
rect 559322 280170 559378 280226
rect 559198 280046 559254 280102
rect 559322 280046 559378 280102
rect 559198 279922 559254 279978
rect 559322 279922 559378 279978
rect 359518 274294 359574 274350
rect 359642 274294 359698 274350
rect 359518 274170 359574 274226
rect 359642 274170 359698 274226
rect 359518 274046 359574 274102
rect 359642 274046 359698 274102
rect 359518 273922 359574 273978
rect 359642 273922 359698 273978
rect 390238 274294 390294 274350
rect 390362 274294 390418 274350
rect 390238 274170 390294 274226
rect 390362 274170 390418 274226
rect 390238 274046 390294 274102
rect 390362 274046 390418 274102
rect 390238 273922 390294 273978
rect 390362 273922 390418 273978
rect 420958 274294 421014 274350
rect 421082 274294 421138 274350
rect 420958 274170 421014 274226
rect 421082 274170 421138 274226
rect 420958 274046 421014 274102
rect 421082 274046 421138 274102
rect 420958 273922 421014 273978
rect 421082 273922 421138 273978
rect 451678 274294 451734 274350
rect 451802 274294 451858 274350
rect 451678 274170 451734 274226
rect 451802 274170 451858 274226
rect 451678 274046 451734 274102
rect 451802 274046 451858 274102
rect 451678 273922 451734 273978
rect 451802 273922 451858 273978
rect 482398 274294 482454 274350
rect 482522 274294 482578 274350
rect 482398 274170 482454 274226
rect 482522 274170 482578 274226
rect 482398 274046 482454 274102
rect 482522 274046 482578 274102
rect 482398 273922 482454 273978
rect 482522 273922 482578 273978
rect 513118 274294 513174 274350
rect 513242 274294 513298 274350
rect 513118 274170 513174 274226
rect 513242 274170 513298 274226
rect 513118 274046 513174 274102
rect 513242 274046 513298 274102
rect 513118 273922 513174 273978
rect 513242 273922 513298 273978
rect 543838 274294 543894 274350
rect 543962 274294 544018 274350
rect 543838 274170 543894 274226
rect 543962 274170 544018 274226
rect 543838 274046 543894 274102
rect 543962 274046 544018 274102
rect 543838 273922 543894 273978
rect 543962 273922 544018 273978
rect 574558 274294 574614 274350
rect 574682 274294 574738 274350
rect 574558 274170 574614 274226
rect 574682 274170 574738 274226
rect 574558 274046 574614 274102
rect 574682 274046 574738 274102
rect 574558 273922 574614 273978
rect 574682 273922 574738 273978
rect 374878 262294 374934 262350
rect 375002 262294 375058 262350
rect 374878 262170 374934 262226
rect 375002 262170 375058 262226
rect 374878 262046 374934 262102
rect 375002 262046 375058 262102
rect 374878 261922 374934 261978
rect 375002 261922 375058 261978
rect 405598 262294 405654 262350
rect 405722 262294 405778 262350
rect 405598 262170 405654 262226
rect 405722 262170 405778 262226
rect 405598 262046 405654 262102
rect 405722 262046 405778 262102
rect 405598 261922 405654 261978
rect 405722 261922 405778 261978
rect 436318 262294 436374 262350
rect 436442 262294 436498 262350
rect 436318 262170 436374 262226
rect 436442 262170 436498 262226
rect 436318 262046 436374 262102
rect 436442 262046 436498 262102
rect 436318 261922 436374 261978
rect 436442 261922 436498 261978
rect 467038 262294 467094 262350
rect 467162 262294 467218 262350
rect 467038 262170 467094 262226
rect 467162 262170 467218 262226
rect 467038 262046 467094 262102
rect 467162 262046 467218 262102
rect 467038 261922 467094 261978
rect 467162 261922 467218 261978
rect 497758 262294 497814 262350
rect 497882 262294 497938 262350
rect 497758 262170 497814 262226
rect 497882 262170 497938 262226
rect 497758 262046 497814 262102
rect 497882 262046 497938 262102
rect 497758 261922 497814 261978
rect 497882 261922 497938 261978
rect 528478 262294 528534 262350
rect 528602 262294 528658 262350
rect 528478 262170 528534 262226
rect 528602 262170 528658 262226
rect 528478 262046 528534 262102
rect 528602 262046 528658 262102
rect 528478 261922 528534 261978
rect 528602 261922 528658 261978
rect 559198 262294 559254 262350
rect 559322 262294 559378 262350
rect 559198 262170 559254 262226
rect 559322 262170 559378 262226
rect 559198 262046 559254 262102
rect 559322 262046 559378 262102
rect 559198 261922 559254 261978
rect 559322 261922 559378 261978
rect 359518 256294 359574 256350
rect 359642 256294 359698 256350
rect 359518 256170 359574 256226
rect 359642 256170 359698 256226
rect 359518 256046 359574 256102
rect 359642 256046 359698 256102
rect 359518 255922 359574 255978
rect 359642 255922 359698 255978
rect 390238 256294 390294 256350
rect 390362 256294 390418 256350
rect 390238 256170 390294 256226
rect 390362 256170 390418 256226
rect 390238 256046 390294 256102
rect 390362 256046 390418 256102
rect 390238 255922 390294 255978
rect 390362 255922 390418 255978
rect 420958 256294 421014 256350
rect 421082 256294 421138 256350
rect 420958 256170 421014 256226
rect 421082 256170 421138 256226
rect 420958 256046 421014 256102
rect 421082 256046 421138 256102
rect 420958 255922 421014 255978
rect 421082 255922 421138 255978
rect 451678 256294 451734 256350
rect 451802 256294 451858 256350
rect 451678 256170 451734 256226
rect 451802 256170 451858 256226
rect 451678 256046 451734 256102
rect 451802 256046 451858 256102
rect 451678 255922 451734 255978
rect 451802 255922 451858 255978
rect 482398 256294 482454 256350
rect 482522 256294 482578 256350
rect 482398 256170 482454 256226
rect 482522 256170 482578 256226
rect 482398 256046 482454 256102
rect 482522 256046 482578 256102
rect 482398 255922 482454 255978
rect 482522 255922 482578 255978
rect 513118 256294 513174 256350
rect 513242 256294 513298 256350
rect 513118 256170 513174 256226
rect 513242 256170 513298 256226
rect 513118 256046 513174 256102
rect 513242 256046 513298 256102
rect 513118 255922 513174 255978
rect 513242 255922 513298 255978
rect 543838 256294 543894 256350
rect 543962 256294 544018 256350
rect 543838 256170 543894 256226
rect 543962 256170 544018 256226
rect 543838 256046 543894 256102
rect 543962 256046 544018 256102
rect 543838 255922 543894 255978
rect 543962 255922 544018 255978
rect 574558 256294 574614 256350
rect 574682 256294 574738 256350
rect 574558 256170 574614 256226
rect 574682 256170 574738 256226
rect 574558 256046 574614 256102
rect 574682 256046 574738 256102
rect 574558 255922 574614 255978
rect 574682 255922 574738 255978
rect 374878 244294 374934 244350
rect 375002 244294 375058 244350
rect 374878 244170 374934 244226
rect 375002 244170 375058 244226
rect 374878 244046 374934 244102
rect 375002 244046 375058 244102
rect 374878 243922 374934 243978
rect 375002 243922 375058 243978
rect 405598 244294 405654 244350
rect 405722 244294 405778 244350
rect 405598 244170 405654 244226
rect 405722 244170 405778 244226
rect 405598 244046 405654 244102
rect 405722 244046 405778 244102
rect 405598 243922 405654 243978
rect 405722 243922 405778 243978
rect 436318 244294 436374 244350
rect 436442 244294 436498 244350
rect 436318 244170 436374 244226
rect 436442 244170 436498 244226
rect 436318 244046 436374 244102
rect 436442 244046 436498 244102
rect 436318 243922 436374 243978
rect 436442 243922 436498 243978
rect 467038 244294 467094 244350
rect 467162 244294 467218 244350
rect 467038 244170 467094 244226
rect 467162 244170 467218 244226
rect 467038 244046 467094 244102
rect 467162 244046 467218 244102
rect 467038 243922 467094 243978
rect 467162 243922 467218 243978
rect 497758 244294 497814 244350
rect 497882 244294 497938 244350
rect 497758 244170 497814 244226
rect 497882 244170 497938 244226
rect 497758 244046 497814 244102
rect 497882 244046 497938 244102
rect 497758 243922 497814 243978
rect 497882 243922 497938 243978
rect 528478 244294 528534 244350
rect 528602 244294 528658 244350
rect 528478 244170 528534 244226
rect 528602 244170 528658 244226
rect 528478 244046 528534 244102
rect 528602 244046 528658 244102
rect 528478 243922 528534 243978
rect 528602 243922 528658 243978
rect 559198 244294 559254 244350
rect 559322 244294 559378 244350
rect 559198 244170 559254 244226
rect 559322 244170 559378 244226
rect 559198 244046 559254 244102
rect 559322 244046 559378 244102
rect 559198 243922 559254 243978
rect 559322 243922 559378 243978
rect 359518 238294 359574 238350
rect 359642 238294 359698 238350
rect 359518 238170 359574 238226
rect 359642 238170 359698 238226
rect 359518 238046 359574 238102
rect 359642 238046 359698 238102
rect 359518 237922 359574 237978
rect 359642 237922 359698 237978
rect 390238 238294 390294 238350
rect 390362 238294 390418 238350
rect 390238 238170 390294 238226
rect 390362 238170 390418 238226
rect 390238 238046 390294 238102
rect 390362 238046 390418 238102
rect 390238 237922 390294 237978
rect 390362 237922 390418 237978
rect 420958 238294 421014 238350
rect 421082 238294 421138 238350
rect 420958 238170 421014 238226
rect 421082 238170 421138 238226
rect 420958 238046 421014 238102
rect 421082 238046 421138 238102
rect 420958 237922 421014 237978
rect 421082 237922 421138 237978
rect 451678 238294 451734 238350
rect 451802 238294 451858 238350
rect 451678 238170 451734 238226
rect 451802 238170 451858 238226
rect 451678 238046 451734 238102
rect 451802 238046 451858 238102
rect 451678 237922 451734 237978
rect 451802 237922 451858 237978
rect 482398 238294 482454 238350
rect 482522 238294 482578 238350
rect 482398 238170 482454 238226
rect 482522 238170 482578 238226
rect 482398 238046 482454 238102
rect 482522 238046 482578 238102
rect 482398 237922 482454 237978
rect 482522 237922 482578 237978
rect 513118 238294 513174 238350
rect 513242 238294 513298 238350
rect 513118 238170 513174 238226
rect 513242 238170 513298 238226
rect 513118 238046 513174 238102
rect 513242 238046 513298 238102
rect 513118 237922 513174 237978
rect 513242 237922 513298 237978
rect 543838 238294 543894 238350
rect 543962 238294 544018 238350
rect 543838 238170 543894 238226
rect 543962 238170 544018 238226
rect 543838 238046 543894 238102
rect 543962 238046 544018 238102
rect 543838 237922 543894 237978
rect 543962 237922 544018 237978
rect 574558 238294 574614 238350
rect 574682 238294 574738 238350
rect 574558 238170 574614 238226
rect 574682 238170 574738 238226
rect 574558 238046 574614 238102
rect 574682 238046 574738 238102
rect 574558 237922 574614 237978
rect 574682 237922 574738 237978
rect 374878 226294 374934 226350
rect 375002 226294 375058 226350
rect 374878 226170 374934 226226
rect 375002 226170 375058 226226
rect 374878 226046 374934 226102
rect 375002 226046 375058 226102
rect 374878 225922 374934 225978
rect 375002 225922 375058 225978
rect 405598 226294 405654 226350
rect 405722 226294 405778 226350
rect 405598 226170 405654 226226
rect 405722 226170 405778 226226
rect 405598 226046 405654 226102
rect 405722 226046 405778 226102
rect 405598 225922 405654 225978
rect 405722 225922 405778 225978
rect 436318 226294 436374 226350
rect 436442 226294 436498 226350
rect 436318 226170 436374 226226
rect 436442 226170 436498 226226
rect 436318 226046 436374 226102
rect 436442 226046 436498 226102
rect 436318 225922 436374 225978
rect 436442 225922 436498 225978
rect 467038 226294 467094 226350
rect 467162 226294 467218 226350
rect 467038 226170 467094 226226
rect 467162 226170 467218 226226
rect 467038 226046 467094 226102
rect 467162 226046 467218 226102
rect 467038 225922 467094 225978
rect 467162 225922 467218 225978
rect 497758 226294 497814 226350
rect 497882 226294 497938 226350
rect 497758 226170 497814 226226
rect 497882 226170 497938 226226
rect 497758 226046 497814 226102
rect 497882 226046 497938 226102
rect 497758 225922 497814 225978
rect 497882 225922 497938 225978
rect 528478 226294 528534 226350
rect 528602 226294 528658 226350
rect 528478 226170 528534 226226
rect 528602 226170 528658 226226
rect 528478 226046 528534 226102
rect 528602 226046 528658 226102
rect 528478 225922 528534 225978
rect 528602 225922 528658 225978
rect 559198 226294 559254 226350
rect 559322 226294 559378 226350
rect 559198 226170 559254 226226
rect 559322 226170 559378 226226
rect 559198 226046 559254 226102
rect 559322 226046 559378 226102
rect 559198 225922 559254 225978
rect 559322 225922 559378 225978
rect 359518 220294 359574 220350
rect 359642 220294 359698 220350
rect 359518 220170 359574 220226
rect 359642 220170 359698 220226
rect 359518 220046 359574 220102
rect 359642 220046 359698 220102
rect 359518 219922 359574 219978
rect 359642 219922 359698 219978
rect 390238 220294 390294 220350
rect 390362 220294 390418 220350
rect 390238 220170 390294 220226
rect 390362 220170 390418 220226
rect 390238 220046 390294 220102
rect 390362 220046 390418 220102
rect 390238 219922 390294 219978
rect 390362 219922 390418 219978
rect 420958 220294 421014 220350
rect 421082 220294 421138 220350
rect 420958 220170 421014 220226
rect 421082 220170 421138 220226
rect 420958 220046 421014 220102
rect 421082 220046 421138 220102
rect 420958 219922 421014 219978
rect 421082 219922 421138 219978
rect 451678 220294 451734 220350
rect 451802 220294 451858 220350
rect 451678 220170 451734 220226
rect 451802 220170 451858 220226
rect 451678 220046 451734 220102
rect 451802 220046 451858 220102
rect 451678 219922 451734 219978
rect 451802 219922 451858 219978
rect 482398 220294 482454 220350
rect 482522 220294 482578 220350
rect 482398 220170 482454 220226
rect 482522 220170 482578 220226
rect 482398 220046 482454 220102
rect 482522 220046 482578 220102
rect 482398 219922 482454 219978
rect 482522 219922 482578 219978
rect 513118 220294 513174 220350
rect 513242 220294 513298 220350
rect 513118 220170 513174 220226
rect 513242 220170 513298 220226
rect 513118 220046 513174 220102
rect 513242 220046 513298 220102
rect 513118 219922 513174 219978
rect 513242 219922 513298 219978
rect 543838 220294 543894 220350
rect 543962 220294 544018 220350
rect 543838 220170 543894 220226
rect 543962 220170 544018 220226
rect 543838 220046 543894 220102
rect 543962 220046 544018 220102
rect 543838 219922 543894 219978
rect 543962 219922 544018 219978
rect 574558 220294 574614 220350
rect 574682 220294 574738 220350
rect 574558 220170 574614 220226
rect 574682 220170 574738 220226
rect 574558 220046 574614 220102
rect 574682 220046 574738 220102
rect 574558 219922 574614 219978
rect 574682 219922 574738 219978
rect 356748 213542 356804 213598
rect 374878 208294 374934 208350
rect 375002 208294 375058 208350
rect 374878 208170 374934 208226
rect 375002 208170 375058 208226
rect 374878 208046 374934 208102
rect 375002 208046 375058 208102
rect 374878 207922 374934 207978
rect 375002 207922 375058 207978
rect 405598 208294 405654 208350
rect 405722 208294 405778 208350
rect 405598 208170 405654 208226
rect 405722 208170 405778 208226
rect 405598 208046 405654 208102
rect 405722 208046 405778 208102
rect 405598 207922 405654 207978
rect 405722 207922 405778 207978
rect 436318 208294 436374 208350
rect 436442 208294 436498 208350
rect 436318 208170 436374 208226
rect 436442 208170 436498 208226
rect 436318 208046 436374 208102
rect 436442 208046 436498 208102
rect 436318 207922 436374 207978
rect 436442 207922 436498 207978
rect 467038 208294 467094 208350
rect 467162 208294 467218 208350
rect 467038 208170 467094 208226
rect 467162 208170 467218 208226
rect 467038 208046 467094 208102
rect 467162 208046 467218 208102
rect 467038 207922 467094 207978
rect 467162 207922 467218 207978
rect 497758 208294 497814 208350
rect 497882 208294 497938 208350
rect 497758 208170 497814 208226
rect 497882 208170 497938 208226
rect 497758 208046 497814 208102
rect 497882 208046 497938 208102
rect 497758 207922 497814 207978
rect 497882 207922 497938 207978
rect 528478 208294 528534 208350
rect 528602 208294 528658 208350
rect 528478 208170 528534 208226
rect 528602 208170 528658 208226
rect 528478 208046 528534 208102
rect 528602 208046 528658 208102
rect 528478 207922 528534 207978
rect 528602 207922 528658 207978
rect 559198 208294 559254 208350
rect 559322 208294 559378 208350
rect 559198 208170 559254 208226
rect 559322 208170 559378 208226
rect 559198 208046 559254 208102
rect 559322 208046 559378 208102
rect 559198 207922 559254 207978
rect 559322 207922 559378 207978
rect 359518 202294 359574 202350
rect 359642 202294 359698 202350
rect 359518 202170 359574 202226
rect 359642 202170 359698 202226
rect 359518 202046 359574 202102
rect 359642 202046 359698 202102
rect 359518 201922 359574 201978
rect 359642 201922 359698 201978
rect 390238 202294 390294 202350
rect 390362 202294 390418 202350
rect 390238 202170 390294 202226
rect 390362 202170 390418 202226
rect 390238 202046 390294 202102
rect 390362 202046 390418 202102
rect 390238 201922 390294 201978
rect 390362 201922 390418 201978
rect 420958 202294 421014 202350
rect 421082 202294 421138 202350
rect 420958 202170 421014 202226
rect 421082 202170 421138 202226
rect 420958 202046 421014 202102
rect 421082 202046 421138 202102
rect 420958 201922 421014 201978
rect 421082 201922 421138 201978
rect 451678 202294 451734 202350
rect 451802 202294 451858 202350
rect 451678 202170 451734 202226
rect 451802 202170 451858 202226
rect 451678 202046 451734 202102
rect 451802 202046 451858 202102
rect 451678 201922 451734 201978
rect 451802 201922 451858 201978
rect 482398 202294 482454 202350
rect 482522 202294 482578 202350
rect 482398 202170 482454 202226
rect 482522 202170 482578 202226
rect 482398 202046 482454 202102
rect 482522 202046 482578 202102
rect 482398 201922 482454 201978
rect 482522 201922 482578 201978
rect 513118 202294 513174 202350
rect 513242 202294 513298 202350
rect 513118 202170 513174 202226
rect 513242 202170 513298 202226
rect 513118 202046 513174 202102
rect 513242 202046 513298 202102
rect 513118 201922 513174 201978
rect 513242 201922 513298 201978
rect 543838 202294 543894 202350
rect 543962 202294 544018 202350
rect 543838 202170 543894 202226
rect 543962 202170 544018 202226
rect 543838 202046 543894 202102
rect 543962 202046 544018 202102
rect 543838 201922 543894 201978
rect 543962 201922 544018 201978
rect 574558 202294 574614 202350
rect 574682 202294 574738 202350
rect 574558 202170 574614 202226
rect 574682 202170 574738 202226
rect 574558 202046 574614 202102
rect 574682 202046 574738 202102
rect 574558 201922 574614 201978
rect 574682 201922 574738 201978
rect 374878 190294 374934 190350
rect 375002 190294 375058 190350
rect 374878 190170 374934 190226
rect 375002 190170 375058 190226
rect 374878 190046 374934 190102
rect 375002 190046 375058 190102
rect 374878 189922 374934 189978
rect 375002 189922 375058 189978
rect 405598 190294 405654 190350
rect 405722 190294 405778 190350
rect 405598 190170 405654 190226
rect 405722 190170 405778 190226
rect 405598 190046 405654 190102
rect 405722 190046 405778 190102
rect 405598 189922 405654 189978
rect 405722 189922 405778 189978
rect 436318 190294 436374 190350
rect 436442 190294 436498 190350
rect 436318 190170 436374 190226
rect 436442 190170 436498 190226
rect 436318 190046 436374 190102
rect 436442 190046 436498 190102
rect 436318 189922 436374 189978
rect 436442 189922 436498 189978
rect 467038 190294 467094 190350
rect 467162 190294 467218 190350
rect 467038 190170 467094 190226
rect 467162 190170 467218 190226
rect 467038 190046 467094 190102
rect 467162 190046 467218 190102
rect 467038 189922 467094 189978
rect 467162 189922 467218 189978
rect 497758 190294 497814 190350
rect 497882 190294 497938 190350
rect 497758 190170 497814 190226
rect 497882 190170 497938 190226
rect 497758 190046 497814 190102
rect 497882 190046 497938 190102
rect 497758 189922 497814 189978
rect 497882 189922 497938 189978
rect 528478 190294 528534 190350
rect 528602 190294 528658 190350
rect 528478 190170 528534 190226
rect 528602 190170 528658 190226
rect 528478 190046 528534 190102
rect 528602 190046 528658 190102
rect 528478 189922 528534 189978
rect 528602 189922 528658 189978
rect 559198 190294 559254 190350
rect 559322 190294 559378 190350
rect 559198 190170 559254 190226
rect 559322 190170 559378 190226
rect 559198 190046 559254 190102
rect 559322 190046 559378 190102
rect 559198 189922 559254 189978
rect 559322 189922 559378 189978
rect 359518 184294 359574 184350
rect 359642 184294 359698 184350
rect 359518 184170 359574 184226
rect 359642 184170 359698 184226
rect 359518 184046 359574 184102
rect 359642 184046 359698 184102
rect 359518 183922 359574 183978
rect 359642 183922 359698 183978
rect 390238 184294 390294 184350
rect 390362 184294 390418 184350
rect 390238 184170 390294 184226
rect 390362 184170 390418 184226
rect 390238 184046 390294 184102
rect 390362 184046 390418 184102
rect 390238 183922 390294 183978
rect 390362 183922 390418 183978
rect 420958 184294 421014 184350
rect 421082 184294 421138 184350
rect 420958 184170 421014 184226
rect 421082 184170 421138 184226
rect 420958 184046 421014 184102
rect 421082 184046 421138 184102
rect 420958 183922 421014 183978
rect 421082 183922 421138 183978
rect 451678 184294 451734 184350
rect 451802 184294 451858 184350
rect 451678 184170 451734 184226
rect 451802 184170 451858 184226
rect 451678 184046 451734 184102
rect 451802 184046 451858 184102
rect 451678 183922 451734 183978
rect 451802 183922 451858 183978
rect 482398 184294 482454 184350
rect 482522 184294 482578 184350
rect 482398 184170 482454 184226
rect 482522 184170 482578 184226
rect 482398 184046 482454 184102
rect 482522 184046 482578 184102
rect 482398 183922 482454 183978
rect 482522 183922 482578 183978
rect 513118 184294 513174 184350
rect 513242 184294 513298 184350
rect 513118 184170 513174 184226
rect 513242 184170 513298 184226
rect 513118 184046 513174 184102
rect 513242 184046 513298 184102
rect 513118 183922 513174 183978
rect 513242 183922 513298 183978
rect 543838 184294 543894 184350
rect 543962 184294 544018 184350
rect 543838 184170 543894 184226
rect 543962 184170 544018 184226
rect 543838 184046 543894 184102
rect 543962 184046 544018 184102
rect 543838 183922 543894 183978
rect 543962 183922 544018 183978
rect 574558 184294 574614 184350
rect 574682 184294 574738 184350
rect 574558 184170 574614 184226
rect 574682 184170 574738 184226
rect 574558 184046 574614 184102
rect 574682 184046 574738 184102
rect 574558 183922 574614 183978
rect 574682 183922 574738 183978
rect 374878 172294 374934 172350
rect 375002 172294 375058 172350
rect 374878 172170 374934 172226
rect 375002 172170 375058 172226
rect 374878 172046 374934 172102
rect 375002 172046 375058 172102
rect 374878 171922 374934 171978
rect 375002 171922 375058 171978
rect 405598 172294 405654 172350
rect 405722 172294 405778 172350
rect 405598 172170 405654 172226
rect 405722 172170 405778 172226
rect 405598 172046 405654 172102
rect 405722 172046 405778 172102
rect 405598 171922 405654 171978
rect 405722 171922 405778 171978
rect 436318 172294 436374 172350
rect 436442 172294 436498 172350
rect 436318 172170 436374 172226
rect 436442 172170 436498 172226
rect 436318 172046 436374 172102
rect 436442 172046 436498 172102
rect 436318 171922 436374 171978
rect 436442 171922 436498 171978
rect 467038 172294 467094 172350
rect 467162 172294 467218 172350
rect 467038 172170 467094 172226
rect 467162 172170 467218 172226
rect 467038 172046 467094 172102
rect 467162 172046 467218 172102
rect 467038 171922 467094 171978
rect 467162 171922 467218 171978
rect 497758 172294 497814 172350
rect 497882 172294 497938 172350
rect 497758 172170 497814 172226
rect 497882 172170 497938 172226
rect 497758 172046 497814 172102
rect 497882 172046 497938 172102
rect 497758 171922 497814 171978
rect 497882 171922 497938 171978
rect 528478 172294 528534 172350
rect 528602 172294 528658 172350
rect 528478 172170 528534 172226
rect 528602 172170 528658 172226
rect 528478 172046 528534 172102
rect 528602 172046 528658 172102
rect 528478 171922 528534 171978
rect 528602 171922 528658 171978
rect 559198 172294 559254 172350
rect 559322 172294 559378 172350
rect 559198 172170 559254 172226
rect 559322 172170 559378 172226
rect 559198 172046 559254 172102
rect 559322 172046 559378 172102
rect 559198 171922 559254 171978
rect 559322 171922 559378 171978
rect 488908 165482 488964 165538
rect 374154 148294 374210 148350
rect 374278 148294 374334 148350
rect 374402 148294 374458 148350
rect 374526 148294 374582 148350
rect 374154 148170 374210 148226
rect 374278 148170 374334 148226
rect 374402 148170 374458 148226
rect 374526 148170 374582 148226
rect 374154 148046 374210 148102
rect 374278 148046 374334 148102
rect 374402 148046 374458 148102
rect 374526 148046 374582 148102
rect 374154 147922 374210 147978
rect 374278 147922 374334 147978
rect 374402 147922 374458 147978
rect 374526 147922 374582 147978
rect 366268 145908 366324 145918
rect 366268 145862 366324 145908
rect 374154 130294 374210 130350
rect 374278 130294 374334 130350
rect 374402 130294 374458 130350
rect 374526 130294 374582 130350
rect 374154 130170 374210 130226
rect 374278 130170 374334 130226
rect 374402 130170 374458 130226
rect 374526 130170 374582 130226
rect 374154 130046 374210 130102
rect 374278 130046 374334 130102
rect 374402 130046 374458 130102
rect 374526 130046 374582 130102
rect 374154 129922 374210 129978
rect 374278 129922 374334 129978
rect 374402 129922 374458 129978
rect 374526 129922 374582 129978
rect 374154 112294 374210 112350
rect 374278 112294 374334 112350
rect 374402 112294 374458 112350
rect 374526 112294 374582 112350
rect 374154 112170 374210 112226
rect 374278 112170 374334 112226
rect 374402 112170 374458 112226
rect 374526 112170 374582 112226
rect 374154 112046 374210 112102
rect 374278 112046 374334 112102
rect 374402 112046 374458 112102
rect 374526 112046 374582 112102
rect 374154 111922 374210 111978
rect 374278 111922 374334 111978
rect 374402 111922 374458 111978
rect 374526 111922 374582 111978
rect 377874 154294 377930 154350
rect 377998 154294 378054 154350
rect 378122 154294 378178 154350
rect 378246 154294 378302 154350
rect 377874 154170 377930 154226
rect 377998 154170 378054 154226
rect 378122 154170 378178 154226
rect 378246 154170 378302 154226
rect 377874 154046 377930 154102
rect 377998 154046 378054 154102
rect 378122 154046 378178 154102
rect 378246 154046 378302 154102
rect 377874 153922 377930 153978
rect 377998 153922 378054 153978
rect 378122 153922 378178 153978
rect 378246 153922 378302 153978
rect 377874 136294 377930 136350
rect 377998 136294 378054 136350
rect 378122 136294 378178 136350
rect 378246 136294 378302 136350
rect 377874 136170 377930 136226
rect 377998 136170 378054 136226
rect 378122 136170 378178 136226
rect 378246 136170 378302 136226
rect 377874 136046 377930 136102
rect 377998 136046 378054 136102
rect 378122 136046 378178 136102
rect 378246 136046 378302 136102
rect 377874 135922 377930 135978
rect 377998 135922 378054 135978
rect 378122 135922 378178 135978
rect 378246 135922 378302 135978
rect 377874 118294 377930 118350
rect 377998 118294 378054 118350
rect 378122 118294 378178 118350
rect 378246 118294 378302 118350
rect 377874 118170 377930 118226
rect 377998 118170 378054 118226
rect 378122 118170 378178 118226
rect 378246 118170 378302 118226
rect 377874 118046 377930 118102
rect 377998 118046 378054 118102
rect 378122 118046 378178 118102
rect 378246 118046 378302 118102
rect 377874 117922 377930 117978
rect 377998 117922 378054 117978
rect 378122 117922 378178 117978
rect 378246 117922 378302 117978
rect 404874 148294 404930 148350
rect 404998 148294 405054 148350
rect 405122 148294 405178 148350
rect 405246 148294 405302 148350
rect 404874 148170 404930 148226
rect 404998 148170 405054 148226
rect 405122 148170 405178 148226
rect 405246 148170 405302 148226
rect 404874 148046 404930 148102
rect 404998 148046 405054 148102
rect 405122 148046 405178 148102
rect 405246 148046 405302 148102
rect 404874 147922 404930 147978
rect 404998 147922 405054 147978
rect 405122 147922 405178 147978
rect 405246 147922 405302 147978
rect 404874 130294 404930 130350
rect 404998 130294 405054 130350
rect 405122 130294 405178 130350
rect 405246 130294 405302 130350
rect 404874 130170 404930 130226
rect 404998 130170 405054 130226
rect 405122 130170 405178 130226
rect 405246 130170 405302 130226
rect 404874 130046 404930 130102
rect 404998 130046 405054 130102
rect 405122 130046 405178 130102
rect 405246 130046 405302 130102
rect 404874 129922 404930 129978
rect 404998 129922 405054 129978
rect 405122 129922 405178 129978
rect 405246 129922 405302 129978
rect 404874 112294 404930 112350
rect 404998 112294 405054 112350
rect 405122 112294 405178 112350
rect 405246 112294 405302 112350
rect 404874 112170 404930 112226
rect 404998 112170 405054 112226
rect 405122 112170 405178 112226
rect 405246 112170 405302 112226
rect 404874 112046 404930 112102
rect 404998 112046 405054 112102
rect 405122 112046 405178 112102
rect 405246 112046 405302 112102
rect 404874 111922 404930 111978
rect 404998 111922 405054 111978
rect 405122 111922 405178 111978
rect 405246 111922 405302 111978
rect 398188 110042 398244 110098
rect 396508 106622 396564 106678
rect 392364 104102 392420 104158
rect 389228 103922 389284 103978
rect 377874 100294 377930 100350
rect 377998 100294 378054 100350
rect 378122 100294 378178 100350
rect 378246 100294 378302 100350
rect 377874 100170 377930 100226
rect 377998 100170 378054 100226
rect 378122 100170 378178 100226
rect 378246 100170 378302 100226
rect 377874 100046 377930 100102
rect 377998 100046 378054 100102
rect 378122 100046 378178 100102
rect 378246 100046 378302 100102
rect 377874 99922 377930 99978
rect 377998 99922 378054 99978
rect 378122 99922 378178 99978
rect 378246 99922 378302 99978
rect 421596 156302 421652 156358
rect 408594 154294 408650 154350
rect 408718 154294 408774 154350
rect 408842 154294 408898 154350
rect 408966 154294 409022 154350
rect 408594 154170 408650 154226
rect 408718 154170 408774 154226
rect 408842 154170 408898 154226
rect 408966 154170 409022 154226
rect 408594 154046 408650 154102
rect 408718 154046 408774 154102
rect 408842 154046 408898 154102
rect 408966 154046 409022 154102
rect 408594 153922 408650 153978
rect 408718 153922 408774 153978
rect 408842 153922 408898 153978
rect 408966 153922 409022 153978
rect 421708 145682 421764 145738
rect 422492 145502 422548 145558
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 408594 136294 408650 136350
rect 408718 136294 408774 136350
rect 408842 136294 408898 136350
rect 408966 136294 409022 136350
rect 408594 136170 408650 136226
rect 408718 136170 408774 136226
rect 408842 136170 408898 136226
rect 408966 136170 409022 136226
rect 408594 136046 408650 136102
rect 408718 136046 408774 136102
rect 408842 136046 408898 136102
rect 408966 136046 409022 136102
rect 408594 135922 408650 135978
rect 408718 135922 408774 135978
rect 408842 135922 408898 135978
rect 408966 135922 409022 135978
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 423276 122462 423332 122518
rect 408594 118294 408650 118350
rect 408718 118294 408774 118350
rect 408842 118294 408898 118350
rect 408966 118294 409022 118350
rect 408594 118170 408650 118226
rect 408718 118170 408774 118226
rect 408842 118170 408898 118226
rect 408966 118170 409022 118226
rect 408594 118046 408650 118102
rect 408718 118046 408774 118102
rect 408842 118046 408898 118102
rect 408966 118046 409022 118102
rect 408594 117922 408650 117978
rect 408718 117922 408774 117978
rect 408842 117922 408898 117978
rect 408966 117922 409022 117978
rect 408594 100294 408650 100350
rect 408718 100294 408774 100350
rect 408842 100294 408898 100350
rect 408966 100294 409022 100350
rect 408594 100170 408650 100226
rect 408718 100170 408774 100226
rect 408842 100170 408898 100226
rect 408966 100170 409022 100226
rect 408594 100046 408650 100102
rect 408718 100046 408774 100102
rect 408842 100046 408898 100102
rect 408966 100046 409022 100102
rect 408594 99922 408650 99978
rect 408718 99922 408774 99978
rect 408842 99922 408898 99978
rect 408966 99922 409022 99978
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 374518 94294 374574 94350
rect 374642 94294 374698 94350
rect 374518 94170 374574 94226
rect 374642 94170 374698 94226
rect 374518 94046 374574 94102
rect 374642 94046 374698 94102
rect 374518 93922 374574 93978
rect 374642 93922 374698 93978
rect 405238 94294 405294 94350
rect 405362 94294 405418 94350
rect 405238 94170 405294 94226
rect 405362 94170 405418 94226
rect 405238 94046 405294 94102
rect 405362 94046 405418 94102
rect 405238 93922 405294 93978
rect 405362 93922 405418 93978
rect 347154 82294 347210 82350
rect 347278 82294 347334 82350
rect 347402 82294 347458 82350
rect 347526 82294 347582 82350
rect 347154 82170 347210 82226
rect 347278 82170 347334 82226
rect 347402 82170 347458 82226
rect 347526 82170 347582 82226
rect 347154 82046 347210 82102
rect 347278 82046 347334 82102
rect 347402 82046 347458 82102
rect 347526 82046 347582 82102
rect 347154 81922 347210 81978
rect 347278 81922 347334 81978
rect 347402 81922 347458 81978
rect 347526 81922 347582 81978
rect 389878 82294 389934 82350
rect 390002 82294 390058 82350
rect 389878 82170 389934 82226
rect 390002 82170 390058 82226
rect 389878 82046 389934 82102
rect 390002 82046 390058 82102
rect 389878 81922 389934 81978
rect 390002 81922 390058 81978
rect 374518 76294 374574 76350
rect 374642 76294 374698 76350
rect 374518 76170 374574 76226
rect 374642 76170 374698 76226
rect 374518 76046 374574 76102
rect 374642 76046 374698 76102
rect 374518 75922 374574 75978
rect 374642 75922 374698 75978
rect 405238 76294 405294 76350
rect 405362 76294 405418 76350
rect 405238 76170 405294 76226
rect 405362 76170 405418 76226
rect 405238 76046 405294 76102
rect 405362 76046 405418 76102
rect 405238 75922 405294 75978
rect 405362 75922 405418 75978
rect 347154 64294 347210 64350
rect 347278 64294 347334 64350
rect 347402 64294 347458 64350
rect 347526 64294 347582 64350
rect 347154 64170 347210 64226
rect 347278 64170 347334 64226
rect 347402 64170 347458 64226
rect 347526 64170 347582 64226
rect 347154 64046 347210 64102
rect 347278 64046 347334 64102
rect 347402 64046 347458 64102
rect 347526 64046 347582 64102
rect 347154 63922 347210 63978
rect 347278 63922 347334 63978
rect 347402 63922 347458 63978
rect 347526 63922 347582 63978
rect 343434 40294 343490 40350
rect 343558 40294 343614 40350
rect 343682 40294 343738 40350
rect 343806 40294 343862 40350
rect 343434 40170 343490 40226
rect 343558 40170 343614 40226
rect 343682 40170 343738 40226
rect 343806 40170 343862 40226
rect 343434 40046 343490 40102
rect 343558 40046 343614 40102
rect 343682 40046 343738 40102
rect 343806 40046 343862 40102
rect 343434 39922 343490 39978
rect 343558 39922 343614 39978
rect 343682 39922 343738 39978
rect 343806 39922 343862 39978
rect 316434 28294 316490 28350
rect 316558 28294 316614 28350
rect 316682 28294 316738 28350
rect 316806 28294 316862 28350
rect 316434 28170 316490 28226
rect 316558 28170 316614 28226
rect 316682 28170 316738 28226
rect 316806 28170 316862 28226
rect 316434 28046 316490 28102
rect 316558 28046 316614 28102
rect 316682 28046 316738 28102
rect 316806 28046 316862 28102
rect 316434 27922 316490 27978
rect 316558 27922 316614 27978
rect 316682 27922 316738 27978
rect 316806 27922 316862 27978
rect 316434 10294 316490 10350
rect 316558 10294 316614 10350
rect 316682 10294 316738 10350
rect 316806 10294 316862 10350
rect 316434 10170 316490 10226
rect 316558 10170 316614 10226
rect 316682 10170 316738 10226
rect 316806 10170 316862 10226
rect 316434 10046 316490 10102
rect 316558 10046 316614 10102
rect 316682 10046 316738 10102
rect 316806 10046 316862 10102
rect 316434 9922 316490 9978
rect 316558 9922 316614 9978
rect 316682 9922 316738 9978
rect 316806 9922 316862 9978
rect 316434 -1176 316490 -1120
rect 316558 -1176 316614 -1120
rect 316682 -1176 316738 -1120
rect 316806 -1176 316862 -1120
rect 316434 -1300 316490 -1244
rect 316558 -1300 316614 -1244
rect 316682 -1300 316738 -1244
rect 316806 -1300 316862 -1244
rect 316434 -1424 316490 -1368
rect 316558 -1424 316614 -1368
rect 316682 -1424 316738 -1368
rect 316806 -1424 316862 -1368
rect 316434 -1548 316490 -1492
rect 316558 -1548 316614 -1492
rect 316682 -1548 316738 -1492
rect 316806 -1548 316862 -1492
rect 343434 22294 343490 22350
rect 343558 22294 343614 22350
rect 343682 22294 343738 22350
rect 343806 22294 343862 22350
rect 343434 22170 343490 22226
rect 343558 22170 343614 22226
rect 343682 22170 343738 22226
rect 343806 22170 343862 22226
rect 343434 22046 343490 22102
rect 343558 22046 343614 22102
rect 343682 22046 343738 22102
rect 343806 22046 343862 22102
rect 343434 21922 343490 21978
rect 343558 21922 343614 21978
rect 343682 21922 343738 21978
rect 343806 21922 343862 21978
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 389878 64294 389934 64350
rect 390002 64294 390058 64350
rect 389878 64170 389934 64226
rect 390002 64170 390058 64226
rect 389878 64046 389934 64102
rect 390002 64046 390058 64102
rect 389878 63922 389934 63978
rect 390002 63922 390058 63978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 374518 58294 374574 58350
rect 374642 58294 374698 58350
rect 374518 58170 374574 58226
rect 374642 58170 374698 58226
rect 374518 58046 374574 58102
rect 374642 58046 374698 58102
rect 374518 57922 374574 57978
rect 374642 57922 374698 57978
rect 405238 58294 405294 58350
rect 405362 58294 405418 58350
rect 405238 58170 405294 58226
rect 405362 58170 405418 58226
rect 405238 58046 405294 58102
rect 405362 58046 405418 58102
rect 405238 57922 405294 57978
rect 405362 57922 405418 57978
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 347154 46294 347210 46350
rect 347278 46294 347334 46350
rect 347402 46294 347458 46350
rect 347526 46294 347582 46350
rect 347154 46170 347210 46226
rect 347278 46170 347334 46226
rect 347402 46170 347458 46226
rect 347526 46170 347582 46226
rect 347154 46046 347210 46102
rect 347278 46046 347334 46102
rect 347402 46046 347458 46102
rect 347526 46046 347582 46102
rect 347154 45922 347210 45978
rect 347278 45922 347334 45978
rect 347402 45922 347458 45978
rect 347526 45922 347582 45978
rect 347154 28294 347210 28350
rect 347278 28294 347334 28350
rect 347402 28294 347458 28350
rect 347526 28294 347582 28350
rect 347154 28170 347210 28226
rect 347278 28170 347334 28226
rect 347402 28170 347458 28226
rect 347526 28170 347582 28226
rect 347154 28046 347210 28102
rect 347278 28046 347334 28102
rect 347402 28046 347458 28102
rect 347526 28046 347582 28102
rect 347154 27922 347210 27978
rect 347278 27922 347334 27978
rect 347402 27922 347458 27978
rect 347526 27922 347582 27978
rect 347154 10294 347210 10350
rect 347278 10294 347334 10350
rect 347402 10294 347458 10350
rect 347526 10294 347582 10350
rect 347154 10170 347210 10226
rect 347278 10170 347334 10226
rect 347402 10170 347458 10226
rect 347526 10170 347582 10226
rect 347154 10046 347210 10102
rect 347278 10046 347334 10102
rect 347402 10046 347458 10102
rect 347526 10046 347582 10102
rect 347154 9922 347210 9978
rect 347278 9922 347334 9978
rect 347402 9922 347458 9978
rect 347526 9922 347582 9978
rect 347154 -1176 347210 -1120
rect 347278 -1176 347334 -1120
rect 347402 -1176 347458 -1120
rect 347526 -1176 347582 -1120
rect 347154 -1300 347210 -1244
rect 347278 -1300 347334 -1244
rect 347402 -1300 347458 -1244
rect 347526 -1300 347582 -1244
rect 347154 -1424 347210 -1368
rect 347278 -1424 347334 -1368
rect 347402 -1424 347458 -1368
rect 347526 -1424 347582 -1368
rect 347154 -1548 347210 -1492
rect 347278 -1548 347334 -1492
rect 347402 -1548 347458 -1492
rect 347526 -1548 347582 -1492
rect 374154 40294 374210 40350
rect 374278 40294 374334 40350
rect 374402 40294 374458 40350
rect 374526 40294 374582 40350
rect 374154 40170 374210 40226
rect 374278 40170 374334 40226
rect 374402 40170 374458 40226
rect 374526 40170 374582 40226
rect 374154 40046 374210 40102
rect 374278 40046 374334 40102
rect 374402 40046 374458 40102
rect 374526 40046 374582 40102
rect 374154 39922 374210 39978
rect 374278 39922 374334 39978
rect 374402 39922 374458 39978
rect 374526 39922 374582 39978
rect 374154 22294 374210 22350
rect 374278 22294 374334 22350
rect 374402 22294 374458 22350
rect 374526 22294 374582 22350
rect 374154 22170 374210 22226
rect 374278 22170 374334 22226
rect 374402 22170 374458 22226
rect 374526 22170 374582 22226
rect 374154 22046 374210 22102
rect 374278 22046 374334 22102
rect 374402 22046 374458 22102
rect 374526 22046 374582 22102
rect 374154 21922 374210 21978
rect 374278 21922 374334 21978
rect 374402 21922 374458 21978
rect 374526 21922 374582 21978
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 377874 46294 377930 46350
rect 377998 46294 378054 46350
rect 378122 46294 378178 46350
rect 378246 46294 378302 46350
rect 377874 46170 377930 46226
rect 377998 46170 378054 46226
rect 378122 46170 378178 46226
rect 378246 46170 378302 46226
rect 377874 46046 377930 46102
rect 377998 46046 378054 46102
rect 378122 46046 378178 46102
rect 378246 46046 378302 46102
rect 377874 45922 377930 45978
rect 377998 45922 378054 45978
rect 378122 45922 378178 45978
rect 378246 45922 378302 45978
rect 377874 28294 377930 28350
rect 377998 28294 378054 28350
rect 378122 28294 378178 28350
rect 378246 28294 378302 28350
rect 377874 28170 377930 28226
rect 377998 28170 378054 28226
rect 378122 28170 378178 28226
rect 378246 28170 378302 28226
rect 377874 28046 377930 28102
rect 377998 28046 378054 28102
rect 378122 28046 378178 28102
rect 378246 28046 378302 28102
rect 377874 27922 377930 27978
rect 377998 27922 378054 27978
rect 378122 27922 378178 27978
rect 378246 27922 378302 27978
rect 377874 10294 377930 10350
rect 377998 10294 378054 10350
rect 378122 10294 378178 10350
rect 378246 10294 378302 10350
rect 377874 10170 377930 10226
rect 377998 10170 378054 10226
rect 378122 10170 378178 10226
rect 378246 10170 378302 10226
rect 377874 10046 377930 10102
rect 377998 10046 378054 10102
rect 378122 10046 378178 10102
rect 378246 10046 378302 10102
rect 377874 9922 377930 9978
rect 377998 9922 378054 9978
rect 378122 9922 378178 9978
rect 378246 9922 378302 9978
rect 377874 -1176 377930 -1120
rect 377998 -1176 378054 -1120
rect 378122 -1176 378178 -1120
rect 378246 -1176 378302 -1120
rect 377874 -1300 377930 -1244
rect 377998 -1300 378054 -1244
rect 378122 -1300 378178 -1244
rect 378246 -1300 378302 -1244
rect 377874 -1424 377930 -1368
rect 377998 -1424 378054 -1368
rect 378122 -1424 378178 -1368
rect 378246 -1424 378302 -1368
rect 377874 -1548 377930 -1492
rect 377998 -1548 378054 -1492
rect 378122 -1548 378178 -1492
rect 378246 -1548 378302 -1492
rect 404874 40294 404930 40350
rect 404998 40294 405054 40350
rect 405122 40294 405178 40350
rect 405246 40294 405302 40350
rect 404874 40170 404930 40226
rect 404998 40170 405054 40226
rect 405122 40170 405178 40226
rect 405246 40170 405302 40226
rect 404874 40046 404930 40102
rect 404998 40046 405054 40102
rect 405122 40046 405178 40102
rect 405246 40046 405302 40102
rect 404874 39922 404930 39978
rect 404998 39922 405054 39978
rect 405122 39922 405178 39978
rect 405246 39922 405302 39978
rect 404874 22294 404930 22350
rect 404998 22294 405054 22350
rect 405122 22294 405178 22350
rect 405246 22294 405302 22350
rect 404874 22170 404930 22226
rect 404998 22170 405054 22226
rect 405122 22170 405178 22226
rect 405246 22170 405302 22226
rect 404874 22046 404930 22102
rect 404998 22046 405054 22102
rect 405122 22046 405178 22102
rect 405246 22046 405302 22102
rect 404874 21922 404930 21978
rect 404998 21922 405054 21978
rect 405122 21922 405178 21978
rect 405246 21922 405302 21978
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 408594 46294 408650 46350
rect 408718 46294 408774 46350
rect 408842 46294 408898 46350
rect 408966 46294 409022 46350
rect 408594 46170 408650 46226
rect 408718 46170 408774 46226
rect 408842 46170 408898 46226
rect 408966 46170 409022 46226
rect 408594 46046 408650 46102
rect 408718 46046 408774 46102
rect 408842 46046 408898 46102
rect 408966 46046 409022 46102
rect 408594 45922 408650 45978
rect 408718 45922 408774 45978
rect 408842 45922 408898 45978
rect 408966 45922 409022 45978
rect 408594 28294 408650 28350
rect 408718 28294 408774 28350
rect 408842 28294 408898 28350
rect 408966 28294 409022 28350
rect 408594 28170 408650 28226
rect 408718 28170 408774 28226
rect 408842 28170 408898 28226
rect 408966 28170 409022 28226
rect 408594 28046 408650 28102
rect 408718 28046 408774 28102
rect 408842 28046 408898 28102
rect 408966 28046 409022 28102
rect 408594 27922 408650 27978
rect 408718 27922 408774 27978
rect 408842 27922 408898 27978
rect 408966 27922 409022 27978
rect 408594 10294 408650 10350
rect 408718 10294 408774 10350
rect 408842 10294 408898 10350
rect 408966 10294 409022 10350
rect 408594 10170 408650 10226
rect 408718 10170 408774 10226
rect 408842 10170 408898 10226
rect 408966 10170 409022 10226
rect 408594 10046 408650 10102
rect 408718 10046 408774 10102
rect 408842 10046 408898 10102
rect 408966 10046 409022 10102
rect 408594 9922 408650 9978
rect 408718 9922 408774 9978
rect 408842 9922 408898 9978
rect 408966 9922 409022 9978
rect 408594 -1176 408650 -1120
rect 408718 -1176 408774 -1120
rect 408842 -1176 408898 -1120
rect 408966 -1176 409022 -1120
rect 408594 -1300 408650 -1244
rect 408718 -1300 408774 -1244
rect 408842 -1300 408898 -1244
rect 408966 -1300 409022 -1244
rect 408594 -1424 408650 -1368
rect 408718 -1424 408774 -1368
rect 408842 -1424 408898 -1368
rect 408966 -1424 409022 -1368
rect 408594 -1548 408650 -1492
rect 408718 -1548 408774 -1492
rect 408842 -1548 408898 -1492
rect 408966 -1548 409022 -1492
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 457212 151262 457268 151318
rect 456988 150002 457044 150058
rect 487788 164042 487844 164098
rect 460236 157382 460292 157438
rect 460124 156122 460180 156178
rect 460348 154862 460404 154918
rect 458444 154682 458500 154738
rect 461244 156482 461300 156538
rect 460460 145862 460516 145918
rect 460348 144422 460404 144478
rect 460572 144242 460628 144298
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 461132 149822 461188 149878
rect 461244 147662 461300 147718
rect 461692 145682 461748 145738
rect 461580 145502 461636 145558
rect 483756 162422 483812 162478
rect 480396 160802 480452 160858
rect 477036 157562 477092 157618
rect 475692 154862 475748 154918
rect 485100 155582 485156 155638
rect 489244 164762 489300 164818
rect 493164 163862 493220 163918
rect 491820 162242 491876 162298
rect 539308 162782 539364 162838
rect 546476 161162 546532 161218
rect 532364 159542 532420 159598
rect 497868 157742 497924 157798
rect 494508 156482 494564 156538
rect 499884 153602 499940 153658
rect 497308 152882 497364 152938
rect 498540 153422 498596 153478
rect 463708 152522 463764 152578
rect 462924 142622 462980 142678
rect 462812 141002 462868 141058
rect 461132 140822 461188 140878
rect 477036 149822 477092 149878
rect 463596 146042 463652 146098
rect 463036 139382 463092 139438
rect 479878 136294 479934 136350
rect 480002 136294 480058 136350
rect 479878 136170 479934 136226
rect 480002 136170 480058 136226
rect 479878 136046 479934 136102
rect 480002 136046 480058 136102
rect 479878 135922 479934 135978
rect 480002 135922 480058 135978
rect 510598 136294 510654 136350
rect 510722 136294 510778 136350
rect 510598 136170 510654 136226
rect 510722 136170 510778 136226
rect 510598 136046 510654 136102
rect 510722 136046 510778 136102
rect 510598 135922 510654 135978
rect 510722 135922 510778 135978
rect 541318 136294 541374 136350
rect 541442 136294 541498 136350
rect 541318 136170 541374 136226
rect 541442 136170 541498 136226
rect 541318 136046 541374 136102
rect 541442 136046 541498 136102
rect 541318 135922 541374 135978
rect 541442 135922 541498 135978
rect 464518 130294 464574 130350
rect 464642 130294 464698 130350
rect 464518 130170 464574 130226
rect 464642 130170 464698 130226
rect 464518 130046 464574 130102
rect 464642 130046 464698 130102
rect 464518 129922 464574 129978
rect 464642 129922 464698 129978
rect 495238 130294 495294 130350
rect 495362 130294 495418 130350
rect 495238 130170 495294 130226
rect 495362 130170 495418 130226
rect 495238 130046 495294 130102
rect 495362 130046 495418 130102
rect 495238 129922 495294 129978
rect 495362 129922 495418 129978
rect 525958 130294 526014 130350
rect 526082 130294 526138 130350
rect 525958 130170 526014 130226
rect 526082 130170 526138 130226
rect 525958 130046 526014 130102
rect 526082 130046 526138 130102
rect 525958 129922 526014 129978
rect 526082 129922 526138 129978
rect 460684 122462 460740 122518
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 479878 118294 479934 118350
rect 480002 118294 480058 118350
rect 479878 118170 479934 118226
rect 480002 118170 480058 118226
rect 479878 118046 479934 118102
rect 480002 118046 480058 118102
rect 479878 117922 479934 117978
rect 480002 117922 480058 117978
rect 510598 118294 510654 118350
rect 510722 118294 510778 118350
rect 510598 118170 510654 118226
rect 510722 118170 510778 118226
rect 510598 118046 510654 118102
rect 510722 118046 510778 118102
rect 510598 117922 510654 117978
rect 510722 117922 510778 117978
rect 541318 118294 541374 118350
rect 541442 118294 541498 118350
rect 541318 118170 541374 118226
rect 541442 118170 541498 118226
rect 541318 118046 541374 118102
rect 541442 118046 541498 118102
rect 541318 117922 541374 117978
rect 541442 117922 541498 117978
rect 554316 163682 554372 163738
rect 553868 157922 553924 157978
rect 553644 116882 553700 116938
rect 553756 150002 553812 150058
rect 464518 112294 464574 112350
rect 464642 112294 464698 112350
rect 464518 112170 464574 112226
rect 464642 112170 464698 112226
rect 464518 112046 464574 112102
rect 464642 112046 464698 112102
rect 464518 111922 464574 111978
rect 464642 111922 464698 111978
rect 495238 112294 495294 112350
rect 495362 112294 495418 112350
rect 495238 112170 495294 112226
rect 495362 112170 495418 112226
rect 495238 112046 495294 112102
rect 495362 112046 495418 112102
rect 495238 111922 495294 111978
rect 495362 111922 495418 111978
rect 525958 112294 526014 112350
rect 526082 112294 526138 112350
rect 525958 112170 526014 112226
rect 526082 112170 526138 112226
rect 525958 112046 526014 112102
rect 526082 112046 526138 112102
rect 525958 111922 526014 111978
rect 526082 111922 526138 111978
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 457660 98162 457716 98218
rect 457660 94922 457716 94978
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 479878 100294 479934 100350
rect 480002 100294 480058 100350
rect 479878 100170 479934 100226
rect 480002 100170 480058 100226
rect 479878 100046 479934 100102
rect 480002 100046 480058 100102
rect 479878 99922 479934 99978
rect 480002 99922 480058 99978
rect 510598 100294 510654 100350
rect 510722 100294 510778 100350
rect 510598 100170 510654 100226
rect 510722 100170 510778 100226
rect 510598 100046 510654 100102
rect 510722 100046 510778 100102
rect 510598 99922 510654 99978
rect 510722 99922 510778 99978
rect 541318 100294 541374 100350
rect 541442 100294 541498 100350
rect 541318 100170 541374 100226
rect 541442 100170 541498 100226
rect 541318 100046 541374 100102
rect 541442 100046 541498 100102
rect 541318 99922 541374 99978
rect 541442 99922 541498 99978
rect 553196 99602 553252 99658
rect 553308 105362 553364 105418
rect 464518 94294 464574 94350
rect 464642 94294 464698 94350
rect 464518 94170 464574 94226
rect 464642 94170 464698 94226
rect 464518 94046 464574 94102
rect 464642 94046 464698 94102
rect 464518 93922 464574 93978
rect 464642 93922 464698 93978
rect 495238 94294 495294 94350
rect 495362 94294 495418 94350
rect 495238 94170 495294 94226
rect 495362 94170 495418 94226
rect 495238 94046 495294 94102
rect 495362 94046 495418 94102
rect 495238 93922 495294 93978
rect 495362 93922 495418 93978
rect 525958 94294 526014 94350
rect 526082 94294 526138 94350
rect 525958 94170 526014 94226
rect 526082 94170 526138 94226
rect 525958 94046 526014 94102
rect 526082 94046 526138 94102
rect 553756 103922 553812 103978
rect 554540 158822 554596 158878
rect 554428 156302 554484 156358
rect 554092 105362 554148 105418
rect 554316 103922 554372 103978
rect 525958 93922 526014 93978
rect 526082 93922 526138 93978
rect 479878 82294 479934 82350
rect 480002 82294 480058 82350
rect 479878 82170 479934 82226
rect 480002 82170 480058 82226
rect 479878 82046 479934 82102
rect 480002 82046 480058 82102
rect 479878 81922 479934 81978
rect 480002 81922 480058 81978
rect 510598 82294 510654 82350
rect 510722 82294 510778 82350
rect 510598 82170 510654 82226
rect 510722 82170 510778 82226
rect 510598 82046 510654 82102
rect 510722 82046 510778 82102
rect 510598 81922 510654 81978
rect 510722 81922 510778 81978
rect 541318 82294 541374 82350
rect 541442 82294 541498 82350
rect 541318 82170 541374 82226
rect 541442 82170 541498 82226
rect 541318 82046 541374 82102
rect 541442 82046 541498 82102
rect 541318 81922 541374 81978
rect 541442 81922 541498 81978
rect 554316 99602 554372 99658
rect 464518 76294 464574 76350
rect 464642 76294 464698 76350
rect 464518 76170 464574 76226
rect 464642 76170 464698 76226
rect 464518 76046 464574 76102
rect 464642 76046 464698 76102
rect 464518 75922 464574 75978
rect 464642 75922 464698 75978
rect 495238 76294 495294 76350
rect 495362 76294 495418 76350
rect 495238 76170 495294 76226
rect 495362 76170 495418 76226
rect 495238 76046 495294 76102
rect 495362 76046 495418 76102
rect 495238 75922 495294 75978
rect 495362 75922 495418 75978
rect 525958 76294 526014 76350
rect 526082 76294 526138 76350
rect 525958 76170 526014 76226
rect 526082 76170 526138 76226
rect 525958 76046 526014 76102
rect 526082 76046 526138 76102
rect 525958 75922 526014 75978
rect 526082 75922 526138 75978
rect 554764 160622 554820 160678
rect 555212 160442 555268 160498
rect 555100 154682 555156 154738
rect 554988 150542 555044 150598
rect 554876 149642 554932 149698
rect 556108 152882 556164 152938
rect 555212 116900 555268 116938
rect 555212 116882 555268 116900
rect 556332 158642 556388 158698
rect 557788 155402 557844 155458
rect 557900 150362 557956 150418
rect 557788 148562 557844 148618
rect 558236 152162 558292 152218
rect 558124 151982 558180 152038
rect 558474 148294 558530 148350
rect 558598 148294 558654 148350
rect 558722 148294 558778 148350
rect 558846 148294 558902 148350
rect 558474 148170 558530 148226
rect 558598 148170 558654 148226
rect 558722 148170 558778 148226
rect 558846 148170 558902 148226
rect 558474 148046 558530 148102
rect 558598 148046 558654 148102
rect 558722 148046 558778 148102
rect 558846 148046 558902 148102
rect 558474 147922 558530 147978
rect 558598 147922 558654 147978
rect 558722 147922 558778 147978
rect 558846 147922 558902 147978
rect 558474 130294 558530 130350
rect 558598 130294 558654 130350
rect 558722 130294 558778 130350
rect 558846 130294 558902 130350
rect 558474 130170 558530 130226
rect 558598 130170 558654 130226
rect 558722 130170 558778 130226
rect 558846 130170 558902 130226
rect 558474 130046 558530 130102
rect 558598 130046 558654 130102
rect 558722 130046 558778 130102
rect 558846 130046 558902 130102
rect 558474 129922 558530 129978
rect 558598 129922 558654 129978
rect 558722 129922 558778 129978
rect 558846 129922 558902 129978
rect 558474 112294 558530 112350
rect 558598 112294 558654 112350
rect 558722 112294 558778 112350
rect 558846 112294 558902 112350
rect 558474 112170 558530 112226
rect 558598 112170 558654 112226
rect 558722 112170 558778 112226
rect 558846 112170 558902 112226
rect 558474 112046 558530 112102
rect 558598 112046 558654 112102
rect 558722 112046 558778 112102
rect 558846 112046 558902 112102
rect 558474 111922 558530 111978
rect 558598 111922 558654 111978
rect 558722 111922 558778 111978
rect 558846 111922 558902 111978
rect 559132 162062 559188 162118
rect 562194 154294 562250 154350
rect 562318 154294 562374 154350
rect 562442 154294 562498 154350
rect 562566 154294 562622 154350
rect 562194 154170 562250 154226
rect 562318 154170 562374 154226
rect 562442 154170 562498 154226
rect 562566 154170 562622 154226
rect 562194 154046 562250 154102
rect 562318 154046 562374 154102
rect 562442 154046 562498 154102
rect 562566 154046 562622 154102
rect 562194 153922 562250 153978
rect 562318 153922 562374 153978
rect 562442 153922 562498 153978
rect 562566 153922 562622 153978
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 590492 409022 590548 409078
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 590716 409562 590772 409618
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 590828 403982 590884 404038
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 590940 402542 590996 402598
rect 591164 403262 591220 403318
rect 590604 402362 590660 402418
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 586348 398582 586404 398638
rect 584780 395342 584836 395398
rect 584668 394802 584724 394858
rect 562194 136294 562250 136350
rect 562318 136294 562374 136350
rect 562442 136294 562498 136350
rect 562566 136294 562622 136350
rect 562194 136170 562250 136226
rect 562318 136170 562374 136226
rect 562442 136170 562498 136226
rect 562566 136170 562622 136226
rect 562194 136046 562250 136102
rect 562318 136046 562374 136102
rect 562442 136046 562498 136102
rect 562566 136046 562622 136102
rect 562194 135922 562250 135978
rect 562318 135922 562374 135978
rect 562442 135922 562498 135978
rect 562566 135922 562622 135978
rect 562194 118294 562250 118350
rect 562318 118294 562374 118350
rect 562442 118294 562498 118350
rect 562566 118294 562622 118350
rect 562194 118170 562250 118226
rect 562318 118170 562374 118226
rect 562442 118170 562498 118226
rect 562566 118170 562622 118226
rect 562194 118046 562250 118102
rect 562318 118046 562374 118102
rect 562442 118046 562498 118102
rect 562566 118046 562622 118102
rect 562194 117922 562250 117978
rect 562318 117922 562374 117978
rect 562442 117922 562498 117978
rect 562566 117922 562622 117978
rect 562194 100294 562250 100350
rect 562318 100294 562374 100350
rect 562442 100294 562498 100350
rect 562566 100294 562622 100350
rect 562194 100170 562250 100226
rect 562318 100170 562374 100226
rect 562442 100170 562498 100226
rect 562566 100170 562622 100226
rect 562194 100046 562250 100102
rect 562318 100046 562374 100102
rect 562442 100046 562498 100102
rect 562566 100046 562622 100102
rect 562194 99922 562250 99978
rect 562318 99922 562374 99978
rect 562442 99922 562498 99978
rect 562566 99922 562622 99978
rect 558474 94294 558530 94350
rect 558598 94294 558654 94350
rect 558722 94294 558778 94350
rect 558846 94294 558902 94350
rect 558474 94170 558530 94226
rect 558598 94170 558654 94226
rect 558722 94170 558778 94226
rect 558846 94170 558902 94226
rect 558474 94046 558530 94102
rect 558598 94046 558654 94102
rect 558722 94046 558778 94102
rect 558846 94046 558902 94102
rect 558474 93922 558530 93978
rect 558598 93922 558654 93978
rect 558722 93922 558778 93978
rect 558846 93922 558902 93978
rect 558474 76294 558530 76350
rect 558598 76294 558654 76350
rect 558722 76294 558778 76350
rect 558846 76294 558902 76350
rect 558474 76170 558530 76226
rect 558598 76170 558654 76226
rect 558722 76170 558778 76226
rect 558846 76170 558902 76226
rect 558474 76046 558530 76102
rect 558598 76046 558654 76102
rect 558722 76046 558778 76102
rect 558846 76046 558902 76102
rect 558474 75922 558530 75978
rect 558598 75922 558654 75978
rect 558722 75922 558778 75978
rect 558846 75922 558902 75978
rect 479878 64294 479934 64350
rect 480002 64294 480058 64350
rect 479878 64170 479934 64226
rect 480002 64170 480058 64226
rect 479878 64046 479934 64102
rect 480002 64046 480058 64102
rect 479878 63922 479934 63978
rect 480002 63922 480058 63978
rect 510598 64294 510654 64350
rect 510722 64294 510778 64350
rect 510598 64170 510654 64226
rect 510722 64170 510778 64226
rect 510598 64046 510654 64102
rect 510722 64046 510778 64102
rect 510598 63922 510654 63978
rect 510722 63922 510778 63978
rect 541318 64294 541374 64350
rect 541442 64294 541498 64350
rect 541318 64170 541374 64226
rect 541442 64170 541498 64226
rect 541318 64046 541374 64102
rect 541442 64046 541498 64102
rect 541318 63922 541374 63978
rect 541442 63922 541498 63978
rect 464518 58294 464574 58350
rect 464642 58294 464698 58350
rect 464518 58170 464574 58226
rect 464642 58170 464698 58226
rect 464518 58046 464574 58102
rect 464642 58046 464698 58102
rect 464518 57922 464574 57978
rect 464642 57922 464698 57978
rect 495238 58294 495294 58350
rect 495362 58294 495418 58350
rect 495238 58170 495294 58226
rect 495362 58170 495418 58226
rect 495238 58046 495294 58102
rect 495362 58046 495418 58102
rect 495238 57922 495294 57978
rect 495362 57922 495418 57978
rect 525958 58294 526014 58350
rect 526082 58294 526138 58350
rect 525958 58170 526014 58226
rect 526082 58170 526138 58226
rect 525958 58046 526014 58102
rect 526082 58046 526138 58102
rect 525958 57922 526014 57978
rect 526082 57922 526138 57978
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 466314 40294 466370 40350
rect 466438 40294 466494 40350
rect 466562 40294 466618 40350
rect 466686 40294 466742 40350
rect 466314 40170 466370 40226
rect 466438 40170 466494 40226
rect 466562 40170 466618 40226
rect 466686 40170 466742 40226
rect 466314 40046 466370 40102
rect 466438 40046 466494 40102
rect 466562 40046 466618 40102
rect 466686 40046 466742 40102
rect 466314 39922 466370 39978
rect 466438 39922 466494 39978
rect 466562 39922 466618 39978
rect 466686 39922 466742 39978
rect 466314 22294 466370 22350
rect 466438 22294 466494 22350
rect 466562 22294 466618 22350
rect 466686 22294 466742 22350
rect 466314 22170 466370 22226
rect 466438 22170 466494 22226
rect 466562 22170 466618 22226
rect 466686 22170 466742 22226
rect 466314 22046 466370 22102
rect 466438 22046 466494 22102
rect 466562 22046 466618 22102
rect 466686 22046 466742 22102
rect 466314 21922 466370 21978
rect 466438 21922 466494 21978
rect 466562 21922 466618 21978
rect 466686 21922 466742 21978
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 470034 46294 470090 46350
rect 470158 46294 470214 46350
rect 470282 46294 470338 46350
rect 470406 46294 470462 46350
rect 470034 46170 470090 46226
rect 470158 46170 470214 46226
rect 470282 46170 470338 46226
rect 470406 46170 470462 46226
rect 470034 46046 470090 46102
rect 470158 46046 470214 46102
rect 470282 46046 470338 46102
rect 470406 46046 470462 46102
rect 470034 45922 470090 45978
rect 470158 45922 470214 45978
rect 470282 45922 470338 45978
rect 470406 45922 470462 45978
rect 470034 28294 470090 28350
rect 470158 28294 470214 28350
rect 470282 28294 470338 28350
rect 470406 28294 470462 28350
rect 470034 28170 470090 28226
rect 470158 28170 470214 28226
rect 470282 28170 470338 28226
rect 470406 28170 470462 28226
rect 470034 28046 470090 28102
rect 470158 28046 470214 28102
rect 470282 28046 470338 28102
rect 470406 28046 470462 28102
rect 470034 27922 470090 27978
rect 470158 27922 470214 27978
rect 470282 27922 470338 27978
rect 470406 27922 470462 27978
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 497034 40294 497090 40350
rect 497158 40294 497214 40350
rect 497282 40294 497338 40350
rect 497406 40294 497462 40350
rect 497034 40170 497090 40226
rect 497158 40170 497214 40226
rect 497282 40170 497338 40226
rect 497406 40170 497462 40226
rect 497034 40046 497090 40102
rect 497158 40046 497214 40102
rect 497282 40046 497338 40102
rect 497406 40046 497462 40102
rect 497034 39922 497090 39978
rect 497158 39922 497214 39978
rect 497282 39922 497338 39978
rect 497406 39922 497462 39978
rect 497034 22294 497090 22350
rect 497158 22294 497214 22350
rect 497282 22294 497338 22350
rect 497406 22294 497462 22350
rect 497034 22170 497090 22226
rect 497158 22170 497214 22226
rect 497282 22170 497338 22226
rect 497406 22170 497462 22226
rect 497034 22046 497090 22102
rect 497158 22046 497214 22102
rect 497282 22046 497338 22102
rect 497406 22046 497462 22102
rect 497034 21922 497090 21978
rect 497158 21922 497214 21978
rect 497282 21922 497338 21978
rect 497406 21922 497462 21978
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 500754 46294 500810 46350
rect 500878 46294 500934 46350
rect 501002 46294 501058 46350
rect 501126 46294 501182 46350
rect 500754 46170 500810 46226
rect 500878 46170 500934 46226
rect 501002 46170 501058 46226
rect 501126 46170 501182 46226
rect 500754 46046 500810 46102
rect 500878 46046 500934 46102
rect 501002 46046 501058 46102
rect 501126 46046 501182 46102
rect 500754 45922 500810 45978
rect 500878 45922 500934 45978
rect 501002 45922 501058 45978
rect 501126 45922 501182 45978
rect 500754 28294 500810 28350
rect 500878 28294 500934 28350
rect 501002 28294 501058 28350
rect 501126 28294 501182 28350
rect 500754 28170 500810 28226
rect 500878 28170 500934 28226
rect 501002 28170 501058 28226
rect 501126 28170 501182 28226
rect 500754 28046 500810 28102
rect 500878 28046 500934 28102
rect 501002 28046 501058 28102
rect 501126 28046 501182 28102
rect 500754 27922 500810 27978
rect 500878 27922 500934 27978
rect 501002 27922 501058 27978
rect 501126 27922 501182 27978
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 527754 40294 527810 40350
rect 527878 40294 527934 40350
rect 528002 40294 528058 40350
rect 528126 40294 528182 40350
rect 527754 40170 527810 40226
rect 527878 40170 527934 40226
rect 528002 40170 528058 40226
rect 528126 40170 528182 40226
rect 527754 40046 527810 40102
rect 527878 40046 527934 40102
rect 528002 40046 528058 40102
rect 528126 40046 528182 40102
rect 527754 39922 527810 39978
rect 527878 39922 527934 39978
rect 528002 39922 528058 39978
rect 528126 39922 528182 39978
rect 527754 22294 527810 22350
rect 527878 22294 527934 22350
rect 528002 22294 528058 22350
rect 528126 22294 528182 22350
rect 527754 22170 527810 22226
rect 527878 22170 527934 22226
rect 528002 22170 528058 22226
rect 528126 22170 528182 22226
rect 527754 22046 527810 22102
rect 527878 22046 527934 22102
rect 528002 22046 528058 22102
rect 528126 22046 528182 22102
rect 527754 21922 527810 21978
rect 527878 21922 527934 21978
rect 528002 21922 528058 21978
rect 528126 21922 528182 21978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 558474 58294 558530 58350
rect 558598 58294 558654 58350
rect 558722 58294 558778 58350
rect 558846 58294 558902 58350
rect 558474 58170 558530 58226
rect 558598 58170 558654 58226
rect 558722 58170 558778 58226
rect 558846 58170 558902 58226
rect 558474 58046 558530 58102
rect 558598 58046 558654 58102
rect 558722 58046 558778 58102
rect 558846 58046 558902 58102
rect 558474 57922 558530 57978
rect 558598 57922 558654 57978
rect 558722 57922 558778 57978
rect 558846 57922 558902 57978
rect 531474 46294 531530 46350
rect 531598 46294 531654 46350
rect 531722 46294 531778 46350
rect 531846 46294 531902 46350
rect 531474 46170 531530 46226
rect 531598 46170 531654 46226
rect 531722 46170 531778 46226
rect 531846 46170 531902 46226
rect 531474 46046 531530 46102
rect 531598 46046 531654 46102
rect 531722 46046 531778 46102
rect 531846 46046 531902 46102
rect 531474 45922 531530 45978
rect 531598 45922 531654 45978
rect 531722 45922 531778 45978
rect 531846 45922 531902 45978
rect 531474 28294 531530 28350
rect 531598 28294 531654 28350
rect 531722 28294 531778 28350
rect 531846 28294 531902 28350
rect 531474 28170 531530 28226
rect 531598 28170 531654 28226
rect 531722 28170 531778 28226
rect 531846 28170 531902 28226
rect 531474 28046 531530 28102
rect 531598 28046 531654 28102
rect 531722 28046 531778 28102
rect 531846 28046 531902 28102
rect 531474 27922 531530 27978
rect 531598 27922 531654 27978
rect 531722 27922 531778 27978
rect 531846 27922 531902 27978
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 558474 40294 558530 40350
rect 558598 40294 558654 40350
rect 558722 40294 558778 40350
rect 558846 40294 558902 40350
rect 558474 40170 558530 40226
rect 558598 40170 558654 40226
rect 558722 40170 558778 40226
rect 558846 40170 558902 40226
rect 558474 40046 558530 40102
rect 558598 40046 558654 40102
rect 558722 40046 558778 40102
rect 558846 40046 558902 40102
rect 558474 39922 558530 39978
rect 558598 39922 558654 39978
rect 558722 39922 558778 39978
rect 558846 39922 558902 39978
rect 558474 22294 558530 22350
rect 558598 22294 558654 22350
rect 558722 22294 558778 22350
rect 558846 22294 558902 22350
rect 558474 22170 558530 22226
rect 558598 22170 558654 22226
rect 558722 22170 558778 22226
rect 558846 22170 558902 22226
rect 558474 22046 558530 22102
rect 558598 22046 558654 22102
rect 558722 22046 558778 22102
rect 558846 22046 558902 22102
rect 558474 21922 558530 21978
rect 558598 21922 558654 21978
rect 558722 21922 558778 21978
rect 558846 21922 558902 21978
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 562194 82294 562250 82350
rect 562318 82294 562374 82350
rect 562442 82294 562498 82350
rect 562566 82294 562622 82350
rect 562194 82170 562250 82226
rect 562318 82170 562374 82226
rect 562442 82170 562498 82226
rect 562566 82170 562622 82226
rect 562194 82046 562250 82102
rect 562318 82046 562374 82102
rect 562442 82046 562498 82102
rect 562566 82046 562622 82102
rect 562194 81922 562250 81978
rect 562318 81922 562374 81978
rect 562442 81922 562498 81978
rect 562566 81922 562622 81978
rect 562194 64294 562250 64350
rect 562318 64294 562374 64350
rect 562442 64294 562498 64350
rect 562566 64294 562622 64350
rect 562194 64170 562250 64226
rect 562318 64170 562374 64226
rect 562442 64170 562498 64226
rect 562566 64170 562622 64226
rect 562194 64046 562250 64102
rect 562318 64046 562374 64102
rect 562442 64046 562498 64102
rect 562566 64046 562622 64102
rect 562194 63922 562250 63978
rect 562318 63922 562374 63978
rect 562442 63922 562498 63978
rect 562566 63922 562622 63978
rect 562194 46294 562250 46350
rect 562318 46294 562374 46350
rect 562442 46294 562498 46350
rect 562566 46294 562622 46350
rect 562194 46170 562250 46226
rect 562318 46170 562374 46226
rect 562442 46170 562498 46226
rect 562566 46170 562622 46226
rect 562194 46046 562250 46102
rect 562318 46046 562374 46102
rect 562442 46046 562498 46102
rect 562566 46046 562622 46102
rect 562194 45922 562250 45978
rect 562318 45922 562374 45978
rect 562442 45922 562498 45978
rect 562566 45922 562622 45978
rect 562194 28294 562250 28350
rect 562318 28294 562374 28350
rect 562442 28294 562498 28350
rect 562566 28294 562622 28350
rect 562194 28170 562250 28226
rect 562318 28170 562374 28226
rect 562442 28170 562498 28226
rect 562566 28170 562622 28226
rect 562194 28046 562250 28102
rect 562318 28046 562374 28102
rect 562442 28046 562498 28102
rect 562566 28046 562622 28102
rect 562194 27922 562250 27978
rect 562318 27922 562374 27978
rect 562442 27922 562498 27978
rect 562566 27922 562622 27978
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 585452 393902 585508 393958
rect 586460 395162 586516 395218
rect 587132 393722 587188 393778
rect 587356 393362 587412 393418
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 590492 400562 590548 400618
rect 591052 398402 591108 398458
rect 590828 398222 590884 398278
rect 590604 393542 590660 393598
rect 592172 401642 592228 401698
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 590492 164582 590548 164638
rect 590156 152740 590212 152758
rect 590156 152702 590212 152740
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 590492 151262 590548 151318
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 592284 393182 592340 393238
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580063 159114 580102
rect 98102 580046 130346 580063
rect -1916 580007 130346 580046
rect 130402 580007 130470 580063
rect 130526 580007 130594 580063
rect 130650 580007 130718 580063
rect 130774 580046 159114 580063
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect 130774 580007 597980 580046
rect -1916 579978 597980 580007
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579939 159114 579978
rect 98102 579922 130346 579939
rect -1916 579883 130346 579922
rect 130402 579883 130470 579939
rect 130526 579883 130594 579939
rect 130650 579883 130718 579939
rect 130774 579922 159114 579939
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect 130774 579883 597980 579922
rect -1916 579826 597980 579883
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 194518 562350
rect 194574 562294 194642 562350
rect 194698 562294 225238 562350
rect 225294 562294 225362 562350
rect 225418 562294 255958 562350
rect 256014 562294 256082 562350
rect 256138 562294 286678 562350
rect 286734 562294 286802 562350
rect 286858 562294 317398 562350
rect 317454 562294 317522 562350
rect 317578 562294 348118 562350
rect 348174 562294 348242 562350
rect 348298 562294 378838 562350
rect 378894 562294 378962 562350
rect 379018 562294 409558 562350
rect 409614 562294 409682 562350
rect 409738 562294 440278 562350
rect 440334 562294 440402 562350
rect 440458 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 470998 562350
rect 471054 562294 471122 562350
rect 471178 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 501718 562350
rect 501774 562294 501842 562350
rect 501898 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562272 597980 562294
rect -1916 562226 116228 562272
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562216 116228 562226
rect 116284 562216 116352 562272
rect 116408 562216 116476 562272
rect 116532 562216 116600 562272
rect 116656 562216 116724 562272
rect 116780 562216 116848 562272
rect 116904 562216 116972 562272
rect 117028 562216 117096 562272
rect 117152 562216 117220 562272
rect 117276 562216 117344 562272
rect 117400 562216 117468 562272
rect 117524 562216 117592 562272
rect 117648 562216 117716 562272
rect 117772 562216 117840 562272
rect 117896 562216 117964 562272
rect 118020 562216 118088 562272
rect 118144 562216 118212 562272
rect 118268 562216 118336 562272
rect 118392 562216 118460 562272
rect 118516 562216 118584 562272
rect 118640 562216 118708 562272
rect 118764 562216 118832 562272
rect 118888 562216 118956 562272
rect 119012 562216 119080 562272
rect 119136 562216 119204 562272
rect 119260 562216 119328 562272
rect 119384 562216 119452 562272
rect 119508 562216 119576 562272
rect 119632 562216 119700 562272
rect 119756 562216 119824 562272
rect 119880 562216 119948 562272
rect 120004 562216 120072 562272
rect 120128 562216 120196 562272
rect 120252 562216 120320 562272
rect 120376 562216 120444 562272
rect 120500 562216 120568 562272
rect 120624 562216 120692 562272
rect 120748 562216 120816 562272
rect 120872 562216 120940 562272
rect 120996 562216 121064 562272
rect 121120 562216 121188 562272
rect 121244 562216 121312 562272
rect 121368 562216 121436 562272
rect 121492 562216 121560 562272
rect 121616 562216 121684 562272
rect 121740 562216 121808 562272
rect 121864 562216 121932 562272
rect 121988 562216 122056 562272
rect 122112 562216 122180 562272
rect 122236 562216 122304 562272
rect 122360 562216 122428 562272
rect 122484 562216 122552 562272
rect 122608 562216 122676 562272
rect 122732 562216 122800 562272
rect 122856 562216 122924 562272
rect 122980 562216 123048 562272
rect 123104 562216 123172 562272
rect 123228 562216 123296 562272
rect 123352 562216 123420 562272
rect 123476 562216 123544 562272
rect 123600 562216 123668 562272
rect 123724 562216 123792 562272
rect 123848 562216 123916 562272
rect 123972 562216 124040 562272
rect 124096 562216 124164 562272
rect 124220 562216 124288 562272
rect 124344 562216 124412 562272
rect 124468 562216 124536 562272
rect 124592 562216 124660 562272
rect 124716 562216 124784 562272
rect 124840 562216 124908 562272
rect 124964 562216 125032 562272
rect 125088 562216 125156 562272
rect 125212 562216 125280 562272
rect 125336 562216 125404 562272
rect 125460 562216 125528 562272
rect 125584 562216 125652 562272
rect 125708 562216 125776 562272
rect 125832 562216 125900 562272
rect 125956 562216 126024 562272
rect 126080 562216 126148 562272
rect 126204 562216 126272 562272
rect 126328 562216 126396 562272
rect 126452 562216 126520 562272
rect 126576 562216 126644 562272
rect 126700 562216 126768 562272
rect 126824 562216 126892 562272
rect 126948 562216 127016 562272
rect 127072 562216 127140 562272
rect 127196 562216 127264 562272
rect 127320 562216 127388 562272
rect 127444 562216 127512 562272
rect 127568 562216 127636 562272
rect 127692 562216 127760 562272
rect 127816 562216 127884 562272
rect 127940 562216 128008 562272
rect 128064 562216 128132 562272
rect 128188 562216 128256 562272
rect 128312 562216 128380 562272
rect 128436 562216 128504 562272
rect 128560 562216 128628 562272
rect 128684 562216 128752 562272
rect 128808 562216 128876 562272
rect 128932 562216 129000 562272
rect 129056 562216 129124 562272
rect 129180 562216 129248 562272
rect 129304 562216 129372 562272
rect 129428 562216 129496 562272
rect 129552 562216 129620 562272
rect 129676 562216 129744 562272
rect 129800 562216 129868 562272
rect 129924 562216 129992 562272
rect 130048 562216 130116 562272
rect 130172 562216 130240 562272
rect 130296 562216 130364 562272
rect 130420 562216 130488 562272
rect 130544 562216 130612 562272
rect 130668 562216 130736 562272
rect 130792 562216 130860 562272
rect 130916 562216 130984 562272
rect 131040 562216 131108 562272
rect 131164 562216 131232 562272
rect 131288 562216 131356 562272
rect 131412 562216 131480 562272
rect 131536 562216 131604 562272
rect 131660 562216 131728 562272
rect 131784 562216 131852 562272
rect 131908 562216 131976 562272
rect 132032 562216 132100 562272
rect 132156 562216 132224 562272
rect 132280 562216 132348 562272
rect 132404 562216 132472 562272
rect 132528 562216 132596 562272
rect 132652 562226 597980 562272
rect 132652 562216 159114 562226
rect 98102 562170 159114 562216
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 194518 562226
rect 194574 562170 194642 562226
rect 194698 562170 225238 562226
rect 225294 562170 225362 562226
rect 225418 562170 255958 562226
rect 256014 562170 256082 562226
rect 256138 562170 286678 562226
rect 286734 562170 286802 562226
rect 286858 562170 317398 562226
rect 317454 562170 317522 562226
rect 317578 562170 348118 562226
rect 348174 562170 348242 562226
rect 348298 562170 378838 562226
rect 378894 562170 378962 562226
rect 379018 562170 409558 562226
rect 409614 562170 409682 562226
rect 409738 562170 440278 562226
rect 440334 562170 440402 562226
rect 440458 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 470998 562226
rect 471054 562170 471122 562226
rect 471178 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 501718 562226
rect 501774 562170 501842 562226
rect 501898 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562148 597980 562170
rect -1916 562102 116228 562148
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562092 116228 562102
rect 116284 562092 116352 562148
rect 116408 562092 116476 562148
rect 116532 562092 116600 562148
rect 116656 562092 116724 562148
rect 116780 562092 116848 562148
rect 116904 562092 116972 562148
rect 117028 562092 117096 562148
rect 117152 562092 117220 562148
rect 117276 562092 117344 562148
rect 117400 562092 117468 562148
rect 117524 562092 117592 562148
rect 117648 562092 117716 562148
rect 117772 562092 117840 562148
rect 117896 562092 117964 562148
rect 118020 562092 118088 562148
rect 118144 562092 118212 562148
rect 118268 562092 118336 562148
rect 118392 562092 118460 562148
rect 118516 562092 118584 562148
rect 118640 562092 118708 562148
rect 118764 562092 118832 562148
rect 118888 562092 118956 562148
rect 119012 562092 119080 562148
rect 119136 562092 119204 562148
rect 119260 562092 119328 562148
rect 119384 562092 119452 562148
rect 119508 562092 119576 562148
rect 119632 562092 119700 562148
rect 119756 562092 119824 562148
rect 119880 562092 119948 562148
rect 120004 562092 120072 562148
rect 120128 562092 120196 562148
rect 120252 562092 120320 562148
rect 120376 562092 120444 562148
rect 120500 562092 120568 562148
rect 120624 562092 120692 562148
rect 120748 562092 120816 562148
rect 120872 562092 120940 562148
rect 120996 562092 121064 562148
rect 121120 562092 121188 562148
rect 121244 562092 121312 562148
rect 121368 562092 121436 562148
rect 121492 562092 121560 562148
rect 121616 562092 121684 562148
rect 121740 562092 121808 562148
rect 121864 562092 121932 562148
rect 121988 562092 122056 562148
rect 122112 562092 122180 562148
rect 122236 562092 122304 562148
rect 122360 562092 122428 562148
rect 122484 562092 122552 562148
rect 122608 562092 122676 562148
rect 122732 562092 122800 562148
rect 122856 562092 122924 562148
rect 122980 562092 123048 562148
rect 123104 562092 123172 562148
rect 123228 562092 123296 562148
rect 123352 562092 123420 562148
rect 123476 562092 123544 562148
rect 123600 562092 123668 562148
rect 123724 562092 123792 562148
rect 123848 562092 123916 562148
rect 123972 562092 124040 562148
rect 124096 562092 124164 562148
rect 124220 562092 124288 562148
rect 124344 562092 124412 562148
rect 124468 562092 124536 562148
rect 124592 562092 124660 562148
rect 124716 562092 124784 562148
rect 124840 562092 124908 562148
rect 124964 562092 125032 562148
rect 125088 562092 125156 562148
rect 125212 562092 125280 562148
rect 125336 562092 125404 562148
rect 125460 562092 125528 562148
rect 125584 562092 125652 562148
rect 125708 562092 125776 562148
rect 125832 562092 125900 562148
rect 125956 562092 126024 562148
rect 126080 562092 126148 562148
rect 126204 562092 126272 562148
rect 126328 562092 126396 562148
rect 126452 562092 126520 562148
rect 126576 562092 126644 562148
rect 126700 562092 126768 562148
rect 126824 562092 126892 562148
rect 126948 562092 127016 562148
rect 127072 562092 127140 562148
rect 127196 562092 127264 562148
rect 127320 562092 127388 562148
rect 127444 562092 127512 562148
rect 127568 562092 127636 562148
rect 127692 562092 127760 562148
rect 127816 562092 127884 562148
rect 127940 562092 128008 562148
rect 128064 562092 128132 562148
rect 128188 562092 128256 562148
rect 128312 562092 128380 562148
rect 128436 562092 128504 562148
rect 128560 562092 128628 562148
rect 128684 562092 128752 562148
rect 128808 562092 128876 562148
rect 128932 562092 129000 562148
rect 129056 562092 129124 562148
rect 129180 562092 129248 562148
rect 129304 562092 129372 562148
rect 129428 562092 129496 562148
rect 129552 562092 129620 562148
rect 129676 562092 129744 562148
rect 129800 562092 129868 562148
rect 129924 562092 129992 562148
rect 130048 562092 130116 562148
rect 130172 562092 130240 562148
rect 130296 562092 130364 562148
rect 130420 562092 130488 562148
rect 130544 562092 130612 562148
rect 130668 562092 130736 562148
rect 130792 562092 130860 562148
rect 130916 562092 130984 562148
rect 131040 562092 131108 562148
rect 131164 562092 131232 562148
rect 131288 562092 131356 562148
rect 131412 562092 131480 562148
rect 131536 562092 131604 562148
rect 131660 562092 131728 562148
rect 131784 562092 131852 562148
rect 131908 562092 131976 562148
rect 132032 562092 132100 562148
rect 132156 562092 132224 562148
rect 132280 562092 132348 562148
rect 132404 562092 132472 562148
rect 132528 562092 132596 562148
rect 132652 562102 597980 562148
rect 132652 562092 159114 562102
rect 98102 562046 159114 562092
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 194518 562102
rect 194574 562046 194642 562102
rect 194698 562046 225238 562102
rect 225294 562046 225362 562102
rect 225418 562046 255958 562102
rect 256014 562046 256082 562102
rect 256138 562046 286678 562102
rect 286734 562046 286802 562102
rect 286858 562046 317398 562102
rect 317454 562046 317522 562102
rect 317578 562046 348118 562102
rect 348174 562046 348242 562102
rect 348298 562046 378838 562102
rect 378894 562046 378962 562102
rect 379018 562046 409558 562102
rect 409614 562046 409682 562102
rect 409738 562046 440278 562102
rect 440334 562046 440402 562102
rect 440458 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 470998 562102
rect 471054 562046 471122 562102
rect 471178 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 501718 562102
rect 501774 562046 501842 562102
rect 501898 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 562024 597980 562046
rect -1916 561978 116228 562024
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561968 116228 561978
rect 116284 561968 116352 562024
rect 116408 561968 116476 562024
rect 116532 561968 116600 562024
rect 116656 561968 116724 562024
rect 116780 561968 116848 562024
rect 116904 561968 116972 562024
rect 117028 561968 117096 562024
rect 117152 561968 117220 562024
rect 117276 561968 117344 562024
rect 117400 561968 117468 562024
rect 117524 561968 117592 562024
rect 117648 561968 117716 562024
rect 117772 561968 117840 562024
rect 117896 561968 117964 562024
rect 118020 561968 118088 562024
rect 118144 561968 118212 562024
rect 118268 561968 118336 562024
rect 118392 561968 118460 562024
rect 118516 561968 118584 562024
rect 118640 561968 118708 562024
rect 118764 561968 118832 562024
rect 118888 561968 118956 562024
rect 119012 561968 119080 562024
rect 119136 561968 119204 562024
rect 119260 561968 119328 562024
rect 119384 561968 119452 562024
rect 119508 561968 119576 562024
rect 119632 561968 119700 562024
rect 119756 561968 119824 562024
rect 119880 561968 119948 562024
rect 120004 561968 120072 562024
rect 120128 561968 120196 562024
rect 120252 561968 120320 562024
rect 120376 561968 120444 562024
rect 120500 561968 120568 562024
rect 120624 561968 120692 562024
rect 120748 561968 120816 562024
rect 120872 561968 120940 562024
rect 120996 561968 121064 562024
rect 121120 561968 121188 562024
rect 121244 561968 121312 562024
rect 121368 561968 121436 562024
rect 121492 561968 121560 562024
rect 121616 561968 121684 562024
rect 121740 561968 121808 562024
rect 121864 561968 121932 562024
rect 121988 561968 122056 562024
rect 122112 561968 122180 562024
rect 122236 561968 122304 562024
rect 122360 561968 122428 562024
rect 122484 561968 122552 562024
rect 122608 561968 122676 562024
rect 122732 561968 122800 562024
rect 122856 561968 122924 562024
rect 122980 561968 123048 562024
rect 123104 561968 123172 562024
rect 123228 561968 123296 562024
rect 123352 561968 123420 562024
rect 123476 561968 123544 562024
rect 123600 561968 123668 562024
rect 123724 561968 123792 562024
rect 123848 561968 123916 562024
rect 123972 561968 124040 562024
rect 124096 561968 124164 562024
rect 124220 561968 124288 562024
rect 124344 561968 124412 562024
rect 124468 561968 124536 562024
rect 124592 561968 124660 562024
rect 124716 561968 124784 562024
rect 124840 561968 124908 562024
rect 124964 561968 125032 562024
rect 125088 561968 125156 562024
rect 125212 561968 125280 562024
rect 125336 561968 125404 562024
rect 125460 561968 125528 562024
rect 125584 561968 125652 562024
rect 125708 561968 125776 562024
rect 125832 561968 125900 562024
rect 125956 561968 126024 562024
rect 126080 561968 126148 562024
rect 126204 561968 126272 562024
rect 126328 561968 126396 562024
rect 126452 561968 126520 562024
rect 126576 561968 126644 562024
rect 126700 561968 126768 562024
rect 126824 561968 126892 562024
rect 126948 561968 127016 562024
rect 127072 561968 127140 562024
rect 127196 561968 127264 562024
rect 127320 561968 127388 562024
rect 127444 561968 127512 562024
rect 127568 561968 127636 562024
rect 127692 561968 127760 562024
rect 127816 561968 127884 562024
rect 127940 561968 128008 562024
rect 128064 561968 128132 562024
rect 128188 561968 128256 562024
rect 128312 561968 128380 562024
rect 128436 561968 128504 562024
rect 128560 561968 128628 562024
rect 128684 561968 128752 562024
rect 128808 561968 128876 562024
rect 128932 561968 129000 562024
rect 129056 561968 129124 562024
rect 129180 561968 129248 562024
rect 129304 561968 129372 562024
rect 129428 561968 129496 562024
rect 129552 561968 129620 562024
rect 129676 561968 129744 562024
rect 129800 561968 129868 562024
rect 129924 561968 129992 562024
rect 130048 561968 130116 562024
rect 130172 561968 130240 562024
rect 130296 561968 130364 562024
rect 130420 561968 130488 562024
rect 130544 561968 130612 562024
rect 130668 561968 130736 562024
rect 130792 561968 130860 562024
rect 130916 561968 130984 562024
rect 131040 561968 131108 562024
rect 131164 561968 131232 562024
rect 131288 561968 131356 562024
rect 131412 561968 131480 562024
rect 131536 561968 131604 562024
rect 131660 561968 131728 562024
rect 131784 561968 131852 562024
rect 131908 561968 131976 562024
rect 132032 561968 132100 562024
rect 132156 561968 132224 562024
rect 132280 561968 132348 562024
rect 132404 561968 132472 562024
rect 132528 561968 132596 562024
rect 132652 561978 597980 562024
rect 132652 561968 159114 561978
rect 98102 561922 159114 561968
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 194518 561978
rect 194574 561922 194642 561978
rect 194698 561922 225238 561978
rect 225294 561922 225362 561978
rect 225418 561922 255958 561978
rect 256014 561922 256082 561978
rect 256138 561922 286678 561978
rect 286734 561922 286802 561978
rect 286858 561922 317398 561978
rect 317454 561922 317522 561978
rect 317578 561922 348118 561978
rect 348174 561922 348242 561978
rect 348298 561922 378838 561978
rect 378894 561922 378962 561978
rect 379018 561922 409558 561978
rect 409614 561922 409682 561978
rect 409738 561922 440278 561978
rect 440334 561922 440402 561978
rect 440458 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 470998 561978
rect 471054 561922 471122 561978
rect 471178 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 501718 561978
rect 501774 561922 501842 561978
rect 501898 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 209878 550350
rect 209934 550294 210002 550350
rect 210058 550294 240598 550350
rect 240654 550294 240722 550350
rect 240778 550294 271318 550350
rect 271374 550294 271442 550350
rect 271498 550294 302038 550350
rect 302094 550294 302162 550350
rect 302218 550294 332758 550350
rect 332814 550294 332882 550350
rect 332938 550294 363478 550350
rect 363534 550294 363602 550350
rect 363658 550294 394198 550350
rect 394254 550294 394322 550350
rect 394378 550294 424918 550350
rect 424974 550294 425042 550350
rect 425098 550294 455638 550350
rect 455694 550294 455762 550350
rect 455818 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 486358 550350
rect 486414 550294 486482 550350
rect 486538 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 517078 550350
rect 517134 550294 517202 550350
rect 517258 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 209878 550226
rect 209934 550170 210002 550226
rect 210058 550170 240598 550226
rect 240654 550170 240722 550226
rect 240778 550170 271318 550226
rect 271374 550170 271442 550226
rect 271498 550170 302038 550226
rect 302094 550170 302162 550226
rect 302218 550170 332758 550226
rect 332814 550170 332882 550226
rect 332938 550170 363478 550226
rect 363534 550170 363602 550226
rect 363658 550170 394198 550226
rect 394254 550170 394322 550226
rect 394378 550170 424918 550226
rect 424974 550170 425042 550226
rect 425098 550170 455638 550226
rect 455694 550170 455762 550226
rect 455818 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 486358 550226
rect 486414 550170 486482 550226
rect 486538 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 517078 550226
rect 517134 550170 517202 550226
rect 517258 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 209878 550102
rect 209934 550046 210002 550102
rect 210058 550046 240598 550102
rect 240654 550046 240722 550102
rect 240778 550046 271318 550102
rect 271374 550046 271442 550102
rect 271498 550046 302038 550102
rect 302094 550046 302162 550102
rect 302218 550046 332758 550102
rect 332814 550046 332882 550102
rect 332938 550046 363478 550102
rect 363534 550046 363602 550102
rect 363658 550046 394198 550102
rect 394254 550046 394322 550102
rect 394378 550046 424918 550102
rect 424974 550046 425042 550102
rect 425098 550046 455638 550102
rect 455694 550046 455762 550102
rect 455818 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 486358 550102
rect 486414 550046 486482 550102
rect 486538 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 517078 550102
rect 517134 550046 517202 550102
rect 517258 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 209878 549978
rect 209934 549922 210002 549978
rect 210058 549922 240598 549978
rect 240654 549922 240722 549978
rect 240778 549922 271318 549978
rect 271374 549922 271442 549978
rect 271498 549922 302038 549978
rect 302094 549922 302162 549978
rect 302218 549922 332758 549978
rect 332814 549922 332882 549978
rect 332938 549922 363478 549978
rect 363534 549922 363602 549978
rect 363658 549922 394198 549978
rect 394254 549922 394322 549978
rect 394378 549922 424918 549978
rect 424974 549922 425042 549978
rect 425098 549922 455638 549978
rect 455694 549922 455762 549978
rect 455818 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 486358 549978
rect 486414 549922 486482 549978
rect 486538 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 517078 549978
rect 517134 549922 517202 549978
rect 517258 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 194518 544350
rect 194574 544294 194642 544350
rect 194698 544294 225238 544350
rect 225294 544294 225362 544350
rect 225418 544294 255958 544350
rect 256014 544294 256082 544350
rect 256138 544294 286678 544350
rect 286734 544294 286802 544350
rect 286858 544294 317398 544350
rect 317454 544294 317522 544350
rect 317578 544294 348118 544350
rect 348174 544294 348242 544350
rect 348298 544294 378838 544350
rect 378894 544294 378962 544350
rect 379018 544294 409558 544350
rect 409614 544294 409682 544350
rect 409738 544294 440278 544350
rect 440334 544294 440402 544350
rect 440458 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 470998 544350
rect 471054 544294 471122 544350
rect 471178 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 501718 544350
rect 501774 544294 501842 544350
rect 501898 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 194518 544226
rect 194574 544170 194642 544226
rect 194698 544170 225238 544226
rect 225294 544170 225362 544226
rect 225418 544170 255958 544226
rect 256014 544170 256082 544226
rect 256138 544170 286678 544226
rect 286734 544170 286802 544226
rect 286858 544170 317398 544226
rect 317454 544170 317522 544226
rect 317578 544170 348118 544226
rect 348174 544170 348242 544226
rect 348298 544170 378838 544226
rect 378894 544170 378962 544226
rect 379018 544170 409558 544226
rect 409614 544170 409682 544226
rect 409738 544170 440278 544226
rect 440334 544170 440402 544226
rect 440458 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 470998 544226
rect 471054 544170 471122 544226
rect 471178 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 501718 544226
rect 501774 544170 501842 544226
rect 501898 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544058 159114 544102
rect 67382 544046 104348 544058
rect -1916 544002 104348 544046
rect 104404 544002 104472 544058
rect 104528 544002 104596 544058
rect 104652 544002 104720 544058
rect 104776 544002 104844 544058
rect 104900 544002 104968 544058
rect 105024 544002 105092 544058
rect 105148 544002 105216 544058
rect 105272 544002 105340 544058
rect 105396 544002 105464 544058
rect 105520 544002 105588 544058
rect 105644 544002 105712 544058
rect 105768 544002 105836 544058
rect 105892 544002 105960 544058
rect 106016 544002 106084 544058
rect 106140 544002 106208 544058
rect 106264 544002 106332 544058
rect 106388 544002 106456 544058
rect 106512 544002 106580 544058
rect 106636 544002 106704 544058
rect 106760 544002 106828 544058
rect 106884 544002 106952 544058
rect 107008 544002 107076 544058
rect 107132 544002 107200 544058
rect 107256 544002 107324 544058
rect 107380 544002 107448 544058
rect 107504 544002 107572 544058
rect 107628 544002 107696 544058
rect 107752 544002 107820 544058
rect 107876 544002 107944 544058
rect 108000 544002 108068 544058
rect 108124 544002 108192 544058
rect 108248 544002 108316 544058
rect 108372 544002 108440 544058
rect 108496 544002 108564 544058
rect 108620 544002 108688 544058
rect 108744 544002 108812 544058
rect 108868 544002 108936 544058
rect 108992 544002 109060 544058
rect 109116 544002 109184 544058
rect 109240 544002 109308 544058
rect 109364 544002 109432 544058
rect 109488 544002 109556 544058
rect 109612 544002 109680 544058
rect 109736 544002 109804 544058
rect 109860 544002 109928 544058
rect 109984 544002 110052 544058
rect 110108 544002 110176 544058
rect 110232 544002 110300 544058
rect 110356 544002 110424 544058
rect 110480 544002 110548 544058
rect 110604 544002 110672 544058
rect 110728 544002 110796 544058
rect 110852 544002 110920 544058
rect 110976 544002 111044 544058
rect 111100 544002 111168 544058
rect 111224 544002 111292 544058
rect 111348 544002 111416 544058
rect 111472 544002 111540 544058
rect 111596 544002 111664 544058
rect 111720 544002 111788 544058
rect 111844 544002 111912 544058
rect 111968 544002 112036 544058
rect 112092 544002 112160 544058
rect 112216 544002 112284 544058
rect 112340 544002 112408 544058
rect 112464 544002 112532 544058
rect 112588 544002 112656 544058
rect 112712 544002 112780 544058
rect 112836 544002 112904 544058
rect 112960 544002 113028 544058
rect 113084 544002 113152 544058
rect 113208 544002 113276 544058
rect 113332 544002 113400 544058
rect 113456 544002 113524 544058
rect 113580 544002 113648 544058
rect 113704 544002 113772 544058
rect 113828 544002 113896 544058
rect 113952 544002 114020 544058
rect 114076 544002 114144 544058
rect 114200 544002 114268 544058
rect 114324 544002 114392 544058
rect 114448 544002 114516 544058
rect 114572 544002 114640 544058
rect 114696 544002 114764 544058
rect 114820 544002 114888 544058
rect 114944 544002 115012 544058
rect 115068 544002 115136 544058
rect 115192 544002 115260 544058
rect 115316 544002 115384 544058
rect 115440 544002 115508 544058
rect 115564 544002 115632 544058
rect 115688 544002 115756 544058
rect 115812 544002 115880 544058
rect 115936 544002 116004 544058
rect 116060 544002 116128 544058
rect 116184 544002 116252 544058
rect 116308 544002 116376 544058
rect 116432 544002 116500 544058
rect 116556 544002 116624 544058
rect 116680 544002 116748 544058
rect 116804 544002 116872 544058
rect 116928 544002 116996 544058
rect 117052 544002 117120 544058
rect 117176 544002 117244 544058
rect 117300 544002 117368 544058
rect 117424 544002 117492 544058
rect 117548 544002 117616 544058
rect 117672 544002 117740 544058
rect 117796 544002 117864 544058
rect 117920 544002 117988 544058
rect 118044 544002 118112 544058
rect 118168 544002 118236 544058
rect 118292 544002 118360 544058
rect 118416 544002 118484 544058
rect 118540 544002 118608 544058
rect 118664 544002 118732 544058
rect 118788 544002 118856 544058
rect 118912 544002 118980 544058
rect 119036 544002 119104 544058
rect 119160 544002 119228 544058
rect 119284 544002 119352 544058
rect 119408 544002 119476 544058
rect 119532 544002 119600 544058
rect 119656 544002 119724 544058
rect 119780 544002 119848 544058
rect 119904 544002 119972 544058
rect 120028 544002 120096 544058
rect 120152 544002 120220 544058
rect 120276 544002 120344 544058
rect 120400 544002 120468 544058
rect 120524 544002 120592 544058
rect 120648 544002 120716 544058
rect 120772 544002 120840 544058
rect 120896 544002 120964 544058
rect 121020 544002 121088 544058
rect 121144 544002 121212 544058
rect 121268 544002 121336 544058
rect 121392 544002 121460 544058
rect 121516 544002 121584 544058
rect 121640 544002 121708 544058
rect 121764 544002 121832 544058
rect 121888 544002 121956 544058
rect 122012 544002 122080 544058
rect 122136 544002 122204 544058
rect 122260 544002 122328 544058
rect 122384 544002 122452 544058
rect 122508 544002 122576 544058
rect 122632 544002 122700 544058
rect 122756 544002 122824 544058
rect 122880 544002 122948 544058
rect 123004 544002 123072 544058
rect 123128 544002 123196 544058
rect 123252 544002 123320 544058
rect 123376 544002 123444 544058
rect 123500 544002 123568 544058
rect 123624 544002 123692 544058
rect 123748 544002 123816 544058
rect 123872 544002 123940 544058
rect 123996 544002 124064 544058
rect 124120 544002 124188 544058
rect 124244 544002 124312 544058
rect 124368 544002 124436 544058
rect 124492 544002 124560 544058
rect 124616 544002 124684 544058
rect 124740 544002 124808 544058
rect 124864 544002 124932 544058
rect 124988 544002 125056 544058
rect 125112 544002 125180 544058
rect 125236 544002 125304 544058
rect 125360 544002 125428 544058
rect 125484 544002 125552 544058
rect 125608 544002 125676 544058
rect 125732 544002 125800 544058
rect 125856 544002 125924 544058
rect 125980 544002 126048 544058
rect 126104 544002 126172 544058
rect 126228 544002 126296 544058
rect 126352 544046 159114 544058
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 194518 544102
rect 194574 544046 194642 544102
rect 194698 544046 225238 544102
rect 225294 544046 225362 544102
rect 225418 544046 255958 544102
rect 256014 544046 256082 544102
rect 256138 544046 286678 544102
rect 286734 544046 286802 544102
rect 286858 544046 317398 544102
rect 317454 544046 317522 544102
rect 317578 544046 348118 544102
rect 348174 544046 348242 544102
rect 348298 544046 378838 544102
rect 378894 544046 378962 544102
rect 379018 544046 409558 544102
rect 409614 544046 409682 544102
rect 409738 544046 440278 544102
rect 440334 544046 440402 544102
rect 440458 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 470998 544102
rect 471054 544046 471122 544102
rect 471178 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 501718 544102
rect 501774 544046 501842 544102
rect 501898 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect 126352 544002 597980 544046
rect -1916 543978 597980 544002
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 194518 543978
rect 194574 543922 194642 543978
rect 194698 543922 225238 543978
rect 225294 543922 225362 543978
rect 225418 543922 255958 543978
rect 256014 543922 256082 543978
rect 256138 543922 286678 543978
rect 286734 543922 286802 543978
rect 286858 543922 317398 543978
rect 317454 543922 317522 543978
rect 317578 543922 348118 543978
rect 348174 543922 348242 543978
rect 348298 543922 378838 543978
rect 378894 543922 378962 543978
rect 379018 543922 409558 543978
rect 409614 543922 409682 543978
rect 409738 543922 440278 543978
rect 440334 543922 440402 543978
rect 440458 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 470998 543978
rect 471054 543922 471122 543978
rect 471178 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 501718 543978
rect 501774 543922 501842 543978
rect 501898 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532358 597980 532446
rect -1916 532350 66714 532358
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532302 66714 532350
rect 66770 532302 66838 532358
rect 66894 532302 66962 532358
rect 67018 532302 67086 532358
rect 67142 532302 67210 532358
rect 67266 532302 67334 532358
rect 67390 532302 67458 532358
rect 67514 532302 67582 532358
rect 67638 532302 67706 532358
rect 67762 532302 67830 532358
rect 67886 532302 67954 532358
rect 68010 532302 68078 532358
rect 68134 532302 68202 532358
rect 68258 532302 68326 532358
rect 68382 532302 68450 532358
rect 68506 532302 68574 532358
rect 68630 532302 68698 532358
rect 68754 532302 68822 532358
rect 68878 532302 68946 532358
rect 69002 532302 69070 532358
rect 69126 532302 69194 532358
rect 69250 532302 69318 532358
rect 69374 532302 69442 532358
rect 69498 532302 69566 532358
rect 69622 532302 69690 532358
rect 69746 532302 69814 532358
rect 69870 532302 69938 532358
rect 69994 532302 70062 532358
rect 70118 532302 70186 532358
rect 70242 532302 70310 532358
rect 70366 532302 70434 532358
rect 70490 532302 70558 532358
rect 70614 532302 70682 532358
rect 70738 532302 70806 532358
rect 70862 532302 70930 532358
rect 70986 532302 71054 532358
rect 71110 532302 71178 532358
rect 71234 532302 71302 532358
rect 71358 532302 71426 532358
rect 71482 532302 71550 532358
rect 71606 532302 71674 532358
rect 71730 532302 71798 532358
rect 71854 532302 71922 532358
rect 71978 532302 72046 532358
rect 72102 532302 72170 532358
rect 72226 532302 72294 532358
rect 72350 532302 72418 532358
rect 72474 532302 72542 532358
rect 72598 532302 72666 532358
rect 72722 532302 72790 532358
rect 72846 532302 72914 532358
rect 72970 532302 73038 532358
rect 73094 532302 73162 532358
rect 73218 532302 73286 532358
rect 73342 532302 73410 532358
rect 73466 532302 73534 532358
rect 73590 532302 73658 532358
rect 73714 532302 73782 532358
rect 73838 532302 73906 532358
rect 73962 532302 74030 532358
rect 74086 532302 74154 532358
rect 74210 532302 74278 532358
rect 74334 532302 74402 532358
rect 74458 532302 74526 532358
rect 74582 532302 74650 532358
rect 74706 532350 597980 532358
rect 74706 532302 162834 532350
rect 40382 532294 162834 532302
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 209878 532350
rect 209934 532294 210002 532350
rect 210058 532294 240598 532350
rect 240654 532294 240722 532350
rect 240778 532294 271318 532350
rect 271374 532294 271442 532350
rect 271498 532294 302038 532350
rect 302094 532294 302162 532350
rect 302218 532294 332758 532350
rect 332814 532294 332882 532350
rect 332938 532294 363478 532350
rect 363534 532294 363602 532350
rect 363658 532294 394198 532350
rect 394254 532294 394322 532350
rect 394378 532294 424918 532350
rect 424974 532294 425042 532350
rect 425098 532294 455638 532350
rect 455694 532294 455762 532350
rect 455818 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 486358 532350
rect 486414 532294 486482 532350
rect 486538 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 517078 532350
rect 517134 532294 517202 532350
rect 517258 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 209878 532226
rect 209934 532170 210002 532226
rect 210058 532170 240598 532226
rect 240654 532170 240722 532226
rect 240778 532170 271318 532226
rect 271374 532170 271442 532226
rect 271498 532170 302038 532226
rect 302094 532170 302162 532226
rect 302218 532170 332758 532226
rect 332814 532170 332882 532226
rect 332938 532170 363478 532226
rect 363534 532170 363602 532226
rect 363658 532170 394198 532226
rect 394254 532170 394322 532226
rect 394378 532170 424918 532226
rect 424974 532170 425042 532226
rect 425098 532170 455638 532226
rect 455694 532170 455762 532226
rect 455818 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 486358 532226
rect 486414 532170 486482 532226
rect 486538 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 517078 532226
rect 517134 532170 517202 532226
rect 517258 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 209878 532102
rect 209934 532046 210002 532102
rect 210058 532046 240598 532102
rect 240654 532046 240722 532102
rect 240778 532046 271318 532102
rect 271374 532046 271442 532102
rect 271498 532046 302038 532102
rect 302094 532046 302162 532102
rect 302218 532046 332758 532102
rect 332814 532046 332882 532102
rect 332938 532046 363478 532102
rect 363534 532046 363602 532102
rect 363658 532046 394198 532102
rect 394254 532046 394322 532102
rect 394378 532046 424918 532102
rect 424974 532046 425042 532102
rect 425098 532046 455638 532102
rect 455694 532046 455762 532102
rect 455818 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 486358 532102
rect 486414 532046 486482 532102
rect 486538 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 517078 532102
rect 517134 532046 517202 532102
rect 517258 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531998 597980 532046
rect -1916 531978 66506 531998
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531942 66506 531978
rect 66562 531942 66630 531998
rect 66686 531942 66754 531998
rect 66810 531942 66878 531998
rect 66934 531942 67002 531998
rect 67058 531942 67126 531998
rect 67182 531942 67250 531998
rect 67306 531942 67374 531998
rect 67430 531942 67498 531998
rect 67554 531942 67622 531998
rect 67678 531942 67746 531998
rect 67802 531942 67870 531998
rect 67926 531942 67994 531998
rect 68050 531942 68118 531998
rect 68174 531942 68242 531998
rect 68298 531942 68366 531998
rect 68422 531942 68490 531998
rect 68546 531942 68614 531998
rect 68670 531942 68738 531998
rect 68794 531942 68862 531998
rect 68918 531942 68986 531998
rect 69042 531942 69110 531998
rect 69166 531942 69234 531998
rect 69290 531942 69358 531998
rect 69414 531942 69482 531998
rect 69538 531942 69606 531998
rect 69662 531942 69730 531998
rect 69786 531942 69854 531998
rect 69910 531942 69978 531998
rect 70034 531942 70102 531998
rect 70158 531942 70226 531998
rect 70282 531942 70350 531998
rect 70406 531942 70474 531998
rect 70530 531942 70598 531998
rect 70654 531942 70722 531998
rect 70778 531942 70846 531998
rect 70902 531942 70970 531998
rect 71026 531942 71094 531998
rect 71150 531942 71218 531998
rect 71274 531942 71342 531998
rect 71398 531942 71466 531998
rect 71522 531942 71590 531998
rect 71646 531942 71714 531998
rect 71770 531942 71838 531998
rect 71894 531942 71962 531998
rect 72018 531942 72086 531998
rect 72142 531942 72210 531998
rect 72266 531942 72334 531998
rect 72390 531942 72458 531998
rect 72514 531942 72582 531998
rect 72638 531942 72706 531998
rect 72762 531942 72830 531998
rect 72886 531942 72954 531998
rect 73010 531942 73078 531998
rect 73134 531942 73202 531998
rect 73258 531942 73326 531998
rect 73382 531942 73450 531998
rect 73506 531942 73574 531998
rect 73630 531942 73698 531998
rect 73754 531942 73822 531998
rect 73878 531942 73946 531998
rect 74002 531942 74070 531998
rect 74126 531942 74194 531998
rect 74250 531942 74318 531998
rect 74374 531978 597980 531998
rect 74374 531942 162834 531978
rect 40382 531922 162834 531942
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 209878 531978
rect 209934 531922 210002 531978
rect 210058 531922 240598 531978
rect 240654 531922 240722 531978
rect 240778 531922 271318 531978
rect 271374 531922 271442 531978
rect 271498 531922 302038 531978
rect 302094 531922 302162 531978
rect 302218 531922 332758 531978
rect 332814 531922 332882 531978
rect 332938 531922 363478 531978
rect 363534 531922 363602 531978
rect 363658 531922 394198 531978
rect 394254 531922 394322 531978
rect 394378 531922 424918 531978
rect 424974 531922 425042 531978
rect 425098 531922 455638 531978
rect 455694 531922 455762 531978
rect 455818 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 486358 531978
rect 486414 531922 486482 531978
rect 486538 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 517078 531978
rect 517134 531922 517202 531978
rect 517258 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 194518 526350
rect 194574 526294 194642 526350
rect 194698 526294 225238 526350
rect 225294 526294 225362 526350
rect 225418 526294 255958 526350
rect 256014 526294 256082 526350
rect 256138 526294 286678 526350
rect 286734 526294 286802 526350
rect 286858 526294 317398 526350
rect 317454 526294 317522 526350
rect 317578 526294 348118 526350
rect 348174 526294 348242 526350
rect 348298 526294 378838 526350
rect 378894 526294 378962 526350
rect 379018 526294 409558 526350
rect 409614 526294 409682 526350
rect 409738 526294 440278 526350
rect 440334 526294 440402 526350
rect 440458 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 470998 526350
rect 471054 526294 471122 526350
rect 471178 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 501718 526350
rect 501774 526294 501842 526350
rect 501898 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526238 597980 526294
rect -1916 526226 96026 526238
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526182 96026 526226
rect 96082 526182 96150 526238
rect 96206 526182 96274 526238
rect 96330 526182 96398 526238
rect 96454 526182 96522 526238
rect 96578 526182 96646 526238
rect 96702 526182 96770 526238
rect 96826 526182 96894 526238
rect 96950 526182 97018 526238
rect 97074 526182 97142 526238
rect 97198 526182 97266 526238
rect 97322 526182 97390 526238
rect 97446 526182 97514 526238
rect 97570 526182 97638 526238
rect 97694 526182 97762 526238
rect 97818 526182 97886 526238
rect 97942 526182 98010 526238
rect 98066 526182 98134 526238
rect 98190 526182 98258 526238
rect 98314 526182 98382 526238
rect 98438 526182 98506 526238
rect 98562 526182 98630 526238
rect 98686 526182 98754 526238
rect 98810 526182 98878 526238
rect 98934 526182 99002 526238
rect 99058 526182 99126 526238
rect 99182 526182 99250 526238
rect 99306 526182 99374 526238
rect 99430 526182 99498 526238
rect 99554 526182 99622 526238
rect 99678 526182 99746 526238
rect 99802 526182 99870 526238
rect 99926 526182 99994 526238
rect 100050 526182 100118 526238
rect 100174 526182 100242 526238
rect 100298 526182 100366 526238
rect 100422 526182 100490 526238
rect 100546 526182 100614 526238
rect 100670 526182 100738 526238
rect 100794 526182 100862 526238
rect 100918 526182 100986 526238
rect 101042 526182 101110 526238
rect 101166 526182 101234 526238
rect 101290 526182 101358 526238
rect 101414 526182 101482 526238
rect 101538 526182 101606 526238
rect 101662 526182 101730 526238
rect 101786 526182 101854 526238
rect 101910 526182 101978 526238
rect 102034 526182 102102 526238
rect 102158 526182 102226 526238
rect 102282 526182 102350 526238
rect 102406 526182 102474 526238
rect 102530 526182 102598 526238
rect 102654 526182 102722 526238
rect 102778 526182 102846 526238
rect 102902 526182 102970 526238
rect 103026 526182 103094 526238
rect 103150 526182 103218 526238
rect 103274 526182 103342 526238
rect 103398 526182 103466 526238
rect 103522 526182 103590 526238
rect 103646 526182 103714 526238
rect 103770 526182 103838 526238
rect 103894 526182 103962 526238
rect 104018 526182 104086 526238
rect 104142 526182 104210 526238
rect 104266 526182 104334 526238
rect 104390 526182 104458 526238
rect 104514 526182 104582 526238
rect 104638 526182 104706 526238
rect 104762 526182 104830 526238
rect 104886 526182 104954 526238
rect 105010 526182 105078 526238
rect 105134 526182 105202 526238
rect 105258 526182 105326 526238
rect 105382 526182 105450 526238
rect 105506 526182 105574 526238
rect 105630 526182 105698 526238
rect 105754 526182 105822 526238
rect 105878 526182 105946 526238
rect 106002 526182 106070 526238
rect 106126 526182 106194 526238
rect 106250 526182 106318 526238
rect 106374 526182 106442 526238
rect 106498 526182 106566 526238
rect 106622 526182 106690 526238
rect 106746 526182 106814 526238
rect 106870 526182 106938 526238
rect 106994 526182 107062 526238
rect 107118 526182 107186 526238
rect 107242 526182 107310 526238
rect 107366 526182 107434 526238
rect 107490 526182 107558 526238
rect 107614 526182 107682 526238
rect 107738 526182 107806 526238
rect 107862 526182 107930 526238
rect 107986 526182 108054 526238
rect 108110 526182 108178 526238
rect 108234 526182 108302 526238
rect 108358 526182 108426 526238
rect 108482 526182 108550 526238
rect 108606 526182 108674 526238
rect 108730 526182 108798 526238
rect 108854 526182 108922 526238
rect 108978 526182 109046 526238
rect 109102 526182 109170 526238
rect 109226 526182 109294 526238
rect 109350 526182 109418 526238
rect 109474 526182 109542 526238
rect 109598 526182 109666 526238
rect 109722 526182 109790 526238
rect 109846 526182 109914 526238
rect 109970 526182 110038 526238
rect 110094 526182 110162 526238
rect 110218 526182 110286 526238
rect 110342 526182 110410 526238
rect 110466 526182 110534 526238
rect 110590 526182 110658 526238
rect 110714 526182 110782 526238
rect 110838 526182 110906 526238
rect 110962 526182 111030 526238
rect 111086 526182 111154 526238
rect 111210 526182 111278 526238
rect 111334 526182 111402 526238
rect 111458 526182 111526 526238
rect 111582 526182 111650 526238
rect 111706 526182 111774 526238
rect 111830 526182 111898 526238
rect 111954 526182 112022 526238
rect 112078 526182 112146 526238
rect 112202 526182 112270 526238
rect 112326 526182 112394 526238
rect 112450 526182 112518 526238
rect 112574 526182 112642 526238
rect 112698 526182 112766 526238
rect 112822 526182 112890 526238
rect 112946 526182 113014 526238
rect 113070 526182 113138 526238
rect 113194 526182 113262 526238
rect 113318 526182 113386 526238
rect 113442 526182 113510 526238
rect 113566 526182 113634 526238
rect 113690 526182 113758 526238
rect 113814 526182 113882 526238
rect 113938 526182 114006 526238
rect 114062 526182 114130 526238
rect 114186 526182 114254 526238
rect 114310 526182 114378 526238
rect 114434 526182 114502 526238
rect 114558 526182 114626 526238
rect 114682 526182 114750 526238
rect 114806 526182 114874 526238
rect 114930 526182 114998 526238
rect 115054 526226 597980 526238
rect 115054 526182 159114 526226
rect 36662 526170 159114 526182
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 194518 526226
rect 194574 526170 194642 526226
rect 194698 526170 225238 526226
rect 225294 526170 225362 526226
rect 225418 526170 255958 526226
rect 256014 526170 256082 526226
rect 256138 526170 286678 526226
rect 286734 526170 286802 526226
rect 286858 526170 317398 526226
rect 317454 526170 317522 526226
rect 317578 526170 348118 526226
rect 348174 526170 348242 526226
rect 348298 526170 378838 526226
rect 378894 526170 378962 526226
rect 379018 526170 409558 526226
rect 409614 526170 409682 526226
rect 409738 526170 440278 526226
rect 440334 526170 440402 526226
rect 440458 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 470998 526226
rect 471054 526170 471122 526226
rect 471178 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 501718 526226
rect 501774 526170 501842 526226
rect 501898 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 194518 526102
rect 194574 526046 194642 526102
rect 194698 526046 225238 526102
rect 225294 526046 225362 526102
rect 225418 526046 255958 526102
rect 256014 526046 256082 526102
rect 256138 526046 286678 526102
rect 286734 526046 286802 526102
rect 286858 526046 317398 526102
rect 317454 526046 317522 526102
rect 317578 526046 348118 526102
rect 348174 526046 348242 526102
rect 348298 526046 378838 526102
rect 378894 526046 378962 526102
rect 379018 526046 409558 526102
rect 409614 526046 409682 526102
rect 409738 526046 440278 526102
rect 440334 526046 440402 526102
rect 440458 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 470998 526102
rect 471054 526046 471122 526102
rect 471178 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 501718 526102
rect 501774 526046 501842 526102
rect 501898 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 194518 525978
rect 194574 525922 194642 525978
rect 194698 525922 225238 525978
rect 225294 525922 225362 525978
rect 225418 525922 255958 525978
rect 256014 525922 256082 525978
rect 256138 525922 286678 525978
rect 286734 525922 286802 525978
rect 286858 525922 317398 525978
rect 317454 525922 317522 525978
rect 317578 525922 348118 525978
rect 348174 525922 348242 525978
rect 348298 525922 378838 525978
rect 378894 525922 378962 525978
rect 379018 525922 409558 525978
rect 409614 525922 409682 525978
rect 409738 525922 440278 525978
rect 440334 525922 440402 525978
rect 440458 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 470998 525978
rect 471054 525922 471122 525978
rect 471178 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 501718 525978
rect 501774 525922 501842 525978
rect 501898 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525911 597980 525922
rect -1916 525855 95880 525911
rect 95936 525855 96004 525911
rect 96060 525855 96128 525911
rect 96184 525855 96252 525911
rect 96308 525855 96376 525911
rect 96432 525855 96500 525911
rect 96556 525855 96624 525911
rect 96680 525855 96748 525911
rect 96804 525855 96872 525911
rect 96928 525855 96996 525911
rect 97052 525855 97120 525911
rect 97176 525855 97244 525911
rect 97300 525855 97368 525911
rect 97424 525855 97492 525911
rect 97548 525855 97616 525911
rect 97672 525855 97740 525911
rect 97796 525855 97864 525911
rect 97920 525855 97988 525911
rect 98044 525855 98112 525911
rect 98168 525855 98236 525911
rect 98292 525855 98360 525911
rect 98416 525855 98484 525911
rect 98540 525855 98608 525911
rect 98664 525855 98732 525911
rect 98788 525855 98856 525911
rect 98912 525855 98980 525911
rect 99036 525855 99104 525911
rect 99160 525855 99228 525911
rect 99284 525855 99352 525911
rect 99408 525855 99476 525911
rect 99532 525855 99600 525911
rect 99656 525855 99724 525911
rect 99780 525855 99848 525911
rect 99904 525855 99972 525911
rect 100028 525855 100096 525911
rect 100152 525855 100220 525911
rect 100276 525855 100344 525911
rect 100400 525855 100468 525911
rect 100524 525855 100592 525911
rect 100648 525855 100716 525911
rect 100772 525855 100840 525911
rect 100896 525855 100964 525911
rect 101020 525855 101088 525911
rect 101144 525855 101212 525911
rect 101268 525855 101336 525911
rect 101392 525855 101460 525911
rect 101516 525855 101584 525911
rect 101640 525855 101708 525911
rect 101764 525855 101832 525911
rect 101888 525855 101956 525911
rect 102012 525855 102080 525911
rect 102136 525855 102204 525911
rect 102260 525855 102328 525911
rect 102384 525855 102452 525911
rect 102508 525855 102576 525911
rect 102632 525855 102700 525911
rect 102756 525855 102824 525911
rect 102880 525855 102948 525911
rect 103004 525855 103072 525911
rect 103128 525855 103196 525911
rect 103252 525855 103320 525911
rect 103376 525855 103444 525911
rect 103500 525855 103568 525911
rect 103624 525855 103692 525911
rect 103748 525855 103816 525911
rect 103872 525855 103940 525911
rect 103996 525855 104064 525911
rect 104120 525855 104188 525911
rect 104244 525855 104312 525911
rect 104368 525855 104436 525911
rect 104492 525855 104560 525911
rect 104616 525855 104684 525911
rect 104740 525855 104808 525911
rect 104864 525855 104932 525911
rect 104988 525855 105056 525911
rect 105112 525855 105180 525911
rect 105236 525855 105304 525911
rect 105360 525855 105428 525911
rect 105484 525855 105552 525911
rect 105608 525855 105676 525911
rect 105732 525855 105800 525911
rect 105856 525855 105924 525911
rect 105980 525855 106048 525911
rect 106104 525855 106172 525911
rect 106228 525855 106296 525911
rect 106352 525855 106420 525911
rect 106476 525855 106544 525911
rect 106600 525855 106668 525911
rect 106724 525855 106792 525911
rect 106848 525855 106916 525911
rect 106972 525855 107040 525911
rect 107096 525855 107164 525911
rect 107220 525855 107288 525911
rect 107344 525855 107412 525911
rect 107468 525855 107536 525911
rect 107592 525855 107660 525911
rect 107716 525855 107784 525911
rect 107840 525855 107908 525911
rect 107964 525855 108032 525911
rect 108088 525855 108156 525911
rect 108212 525855 108280 525911
rect 108336 525855 108404 525911
rect 108460 525855 108528 525911
rect 108584 525855 108652 525911
rect 108708 525855 108776 525911
rect 108832 525855 108900 525911
rect 108956 525855 109024 525911
rect 109080 525855 109148 525911
rect 109204 525855 109272 525911
rect 109328 525855 109396 525911
rect 109452 525855 109520 525911
rect 109576 525855 109644 525911
rect 109700 525855 109768 525911
rect 109824 525855 109892 525911
rect 109948 525855 110016 525911
rect 110072 525855 110140 525911
rect 110196 525855 110264 525911
rect 110320 525855 110388 525911
rect 110444 525855 110512 525911
rect 110568 525855 110636 525911
rect 110692 525855 110760 525911
rect 110816 525855 110884 525911
rect 110940 525855 111008 525911
rect 111064 525855 111132 525911
rect 111188 525855 111256 525911
rect 111312 525855 111380 525911
rect 111436 525855 111504 525911
rect 111560 525855 111628 525911
rect 111684 525855 111752 525911
rect 111808 525855 111876 525911
rect 111932 525855 112000 525911
rect 112056 525855 112124 525911
rect 112180 525855 112248 525911
rect 112304 525855 112372 525911
rect 112428 525855 112496 525911
rect 112552 525855 112620 525911
rect 112676 525855 112744 525911
rect 112800 525855 112868 525911
rect 112924 525855 112992 525911
rect 113048 525855 113116 525911
rect 113172 525855 113240 525911
rect 113296 525855 113364 525911
rect 113420 525855 113488 525911
rect 113544 525855 113612 525911
rect 113668 525855 113736 525911
rect 113792 525855 113860 525911
rect 113916 525855 113984 525911
rect 114040 525855 114108 525911
rect 114164 525855 114232 525911
rect 114288 525855 114356 525911
rect 114412 525855 114480 525911
rect 114536 525855 114604 525911
rect 114660 525855 597980 525911
rect -1916 525826 597980 525855
rect -1916 514412 597980 514446
rect -1916 514356 60202 514412
rect 60258 514356 60326 514412
rect 60382 514356 60450 514412
rect 60506 514356 60574 514412
rect 60630 514356 60698 514412
rect 60754 514356 60822 514412
rect 60878 514356 60946 514412
rect 61002 514356 61070 514412
rect 61126 514356 61194 514412
rect 61250 514356 61318 514412
rect 61374 514356 61442 514412
rect 61498 514356 61566 514412
rect 61622 514356 61690 514412
rect 61746 514356 61814 514412
rect 61870 514356 61938 514412
rect 61994 514356 62062 514412
rect 62118 514356 62186 514412
rect 62242 514356 62310 514412
rect 62366 514356 62434 514412
rect 62490 514356 62558 514412
rect 62614 514356 62682 514412
rect 62738 514356 62806 514412
rect 62862 514356 62930 514412
rect 62986 514356 63054 514412
rect 63110 514356 63178 514412
rect 63234 514356 63302 514412
rect 63358 514356 63426 514412
rect 63482 514356 63550 514412
rect 63606 514356 63674 514412
rect 63730 514356 63798 514412
rect 63854 514356 63922 514412
rect 63978 514356 64046 514412
rect 64102 514356 64170 514412
rect 64226 514356 64294 514412
rect 64350 514356 64418 514412
rect 64474 514356 64542 514412
rect 64598 514356 64666 514412
rect 64722 514356 64790 514412
rect 64846 514356 64914 514412
rect 64970 514356 65038 514412
rect 65094 514356 65162 514412
rect 65218 514356 65286 514412
rect 65342 514356 65410 514412
rect 65466 514356 65534 514412
rect 65590 514356 65658 514412
rect 65714 514356 65782 514412
rect 65838 514356 65906 514412
rect 65962 514356 66030 514412
rect 66086 514356 66154 514412
rect 66210 514356 66278 514412
rect 66334 514356 66402 514412
rect 66458 514356 597980 514412
rect -1916 514350 597980 514356
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 209878 514350
rect 209934 514294 210002 514350
rect 210058 514294 240598 514350
rect 240654 514294 240722 514350
rect 240778 514294 271318 514350
rect 271374 514294 271442 514350
rect 271498 514294 302038 514350
rect 302094 514294 302162 514350
rect 302218 514294 332758 514350
rect 332814 514294 332882 514350
rect 332938 514294 363478 514350
rect 363534 514294 363602 514350
rect 363658 514294 394198 514350
rect 394254 514294 394322 514350
rect 394378 514294 424918 514350
rect 424974 514294 425042 514350
rect 425098 514294 455638 514350
rect 455694 514294 455762 514350
rect 455818 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 486358 514350
rect 486414 514294 486482 514350
rect 486538 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 517078 514350
rect 517134 514294 517202 514350
rect 517258 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514288 597980 514294
rect -1916 514232 60202 514288
rect 60258 514232 60326 514288
rect 60382 514232 60450 514288
rect 60506 514232 60574 514288
rect 60630 514232 60698 514288
rect 60754 514232 60822 514288
rect 60878 514232 60946 514288
rect 61002 514232 61070 514288
rect 61126 514232 61194 514288
rect 61250 514232 61318 514288
rect 61374 514232 61442 514288
rect 61498 514232 61566 514288
rect 61622 514232 61690 514288
rect 61746 514232 61814 514288
rect 61870 514232 61938 514288
rect 61994 514232 62062 514288
rect 62118 514232 62186 514288
rect 62242 514232 62310 514288
rect 62366 514232 62434 514288
rect 62490 514232 62558 514288
rect 62614 514232 62682 514288
rect 62738 514232 62806 514288
rect 62862 514232 62930 514288
rect 62986 514232 63054 514288
rect 63110 514232 63178 514288
rect 63234 514232 63302 514288
rect 63358 514232 63426 514288
rect 63482 514232 63550 514288
rect 63606 514232 63674 514288
rect 63730 514232 63798 514288
rect 63854 514232 63922 514288
rect 63978 514232 64046 514288
rect 64102 514232 64170 514288
rect 64226 514232 64294 514288
rect 64350 514232 64418 514288
rect 64474 514232 64542 514288
rect 64598 514232 64666 514288
rect 64722 514232 64790 514288
rect 64846 514232 64914 514288
rect 64970 514232 65038 514288
rect 65094 514232 65162 514288
rect 65218 514232 65286 514288
rect 65342 514232 65410 514288
rect 65466 514232 65534 514288
rect 65590 514232 65658 514288
rect 65714 514232 65782 514288
rect 65838 514232 65906 514288
rect 65962 514232 66030 514288
rect 66086 514232 66154 514288
rect 66210 514232 66278 514288
rect 66334 514232 66402 514288
rect 66458 514232 597980 514288
rect -1916 514226 597980 514232
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 209878 514226
rect 209934 514170 210002 514226
rect 210058 514170 240598 514226
rect 240654 514170 240722 514226
rect 240778 514170 271318 514226
rect 271374 514170 271442 514226
rect 271498 514170 302038 514226
rect 302094 514170 302162 514226
rect 302218 514170 332758 514226
rect 332814 514170 332882 514226
rect 332938 514170 363478 514226
rect 363534 514170 363602 514226
rect 363658 514170 394198 514226
rect 394254 514170 394322 514226
rect 394378 514170 424918 514226
rect 424974 514170 425042 514226
rect 425098 514170 455638 514226
rect 455694 514170 455762 514226
rect 455818 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 486358 514226
rect 486414 514170 486482 514226
rect 486538 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 517078 514226
rect 517134 514170 517202 514226
rect 517258 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514164 597980 514170
rect -1916 514108 60202 514164
rect 60258 514108 60326 514164
rect 60382 514108 60450 514164
rect 60506 514108 60574 514164
rect 60630 514108 60698 514164
rect 60754 514108 60822 514164
rect 60878 514108 60946 514164
rect 61002 514108 61070 514164
rect 61126 514108 61194 514164
rect 61250 514108 61318 514164
rect 61374 514108 61442 514164
rect 61498 514108 61566 514164
rect 61622 514108 61690 514164
rect 61746 514108 61814 514164
rect 61870 514108 61938 514164
rect 61994 514108 62062 514164
rect 62118 514108 62186 514164
rect 62242 514108 62310 514164
rect 62366 514108 62434 514164
rect 62490 514108 62558 514164
rect 62614 514108 62682 514164
rect 62738 514108 62806 514164
rect 62862 514108 62930 514164
rect 62986 514108 63054 514164
rect 63110 514108 63178 514164
rect 63234 514108 63302 514164
rect 63358 514108 63426 514164
rect 63482 514108 63550 514164
rect 63606 514108 63674 514164
rect 63730 514108 63798 514164
rect 63854 514108 63922 514164
rect 63978 514108 64046 514164
rect 64102 514108 64170 514164
rect 64226 514108 64294 514164
rect 64350 514108 64418 514164
rect 64474 514108 64542 514164
rect 64598 514108 64666 514164
rect 64722 514108 64790 514164
rect 64846 514108 64914 514164
rect 64970 514108 65038 514164
rect 65094 514108 65162 514164
rect 65218 514108 65286 514164
rect 65342 514108 65410 514164
rect 65466 514108 65534 514164
rect 65590 514108 65658 514164
rect 65714 514108 65782 514164
rect 65838 514108 65906 514164
rect 65962 514108 66030 514164
rect 66086 514108 66154 514164
rect 66210 514108 66278 514164
rect 66334 514108 66402 514164
rect 66458 514108 597980 514164
rect -1916 514102 597980 514108
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 209878 514102
rect 209934 514046 210002 514102
rect 210058 514046 240598 514102
rect 240654 514046 240722 514102
rect 240778 514046 271318 514102
rect 271374 514046 271442 514102
rect 271498 514046 302038 514102
rect 302094 514046 302162 514102
rect 302218 514046 332758 514102
rect 332814 514046 332882 514102
rect 332938 514046 363478 514102
rect 363534 514046 363602 514102
rect 363658 514046 394198 514102
rect 394254 514046 394322 514102
rect 394378 514046 424918 514102
rect 424974 514046 425042 514102
rect 425098 514046 455638 514102
rect 455694 514046 455762 514102
rect 455818 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 486358 514102
rect 486414 514046 486482 514102
rect 486538 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 517078 514102
rect 517134 514046 517202 514102
rect 517258 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 514040 597980 514046
rect -1916 513984 60202 514040
rect 60258 513984 60326 514040
rect 60382 513984 60450 514040
rect 60506 513984 60574 514040
rect 60630 513984 60698 514040
rect 60754 513984 60822 514040
rect 60878 513984 60946 514040
rect 61002 513984 61070 514040
rect 61126 513984 61194 514040
rect 61250 513984 61318 514040
rect 61374 513984 61442 514040
rect 61498 513984 61566 514040
rect 61622 513984 61690 514040
rect 61746 513984 61814 514040
rect 61870 513984 61938 514040
rect 61994 513984 62062 514040
rect 62118 513984 62186 514040
rect 62242 513984 62310 514040
rect 62366 513984 62434 514040
rect 62490 513984 62558 514040
rect 62614 513984 62682 514040
rect 62738 513984 62806 514040
rect 62862 513984 62930 514040
rect 62986 513984 63054 514040
rect 63110 513984 63178 514040
rect 63234 513984 63302 514040
rect 63358 513984 63426 514040
rect 63482 513984 63550 514040
rect 63606 513984 63674 514040
rect 63730 513984 63798 514040
rect 63854 513984 63922 514040
rect 63978 513984 64046 514040
rect 64102 513984 64170 514040
rect 64226 513984 64294 514040
rect 64350 513984 64418 514040
rect 64474 513984 64542 514040
rect 64598 513984 64666 514040
rect 64722 513984 64790 514040
rect 64846 513984 64914 514040
rect 64970 513984 65038 514040
rect 65094 513984 65162 514040
rect 65218 513984 65286 514040
rect 65342 513984 65410 514040
rect 65466 513984 65534 514040
rect 65590 513984 65658 514040
rect 65714 513984 65782 514040
rect 65838 513984 65906 514040
rect 65962 513984 66030 514040
rect 66086 513984 66154 514040
rect 66210 513984 66278 514040
rect 66334 513984 66402 514040
rect 66458 513984 597980 514040
rect -1916 513978 597980 513984
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 209878 513978
rect 209934 513922 210002 513978
rect 210058 513922 240598 513978
rect 240654 513922 240722 513978
rect 240778 513922 271318 513978
rect 271374 513922 271442 513978
rect 271498 513922 302038 513978
rect 302094 513922 302162 513978
rect 302218 513922 332758 513978
rect 332814 513922 332882 513978
rect 332938 513922 363478 513978
rect 363534 513922 363602 513978
rect 363658 513922 394198 513978
rect 394254 513922 394322 513978
rect 394378 513922 424918 513978
rect 424974 513922 425042 513978
rect 425098 513922 455638 513978
rect 455694 513922 455762 513978
rect 455818 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 486358 513978
rect 486414 513922 486482 513978
rect 486538 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 517078 513978
rect 517134 513922 517202 513978
rect 517258 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513916 597980 513922
rect -1916 513860 60202 513916
rect 60258 513860 60326 513916
rect 60382 513860 60450 513916
rect 60506 513860 60574 513916
rect 60630 513860 60698 513916
rect 60754 513860 60822 513916
rect 60878 513860 60946 513916
rect 61002 513860 61070 513916
rect 61126 513860 61194 513916
rect 61250 513860 61318 513916
rect 61374 513860 61442 513916
rect 61498 513860 61566 513916
rect 61622 513860 61690 513916
rect 61746 513860 61814 513916
rect 61870 513860 61938 513916
rect 61994 513860 62062 513916
rect 62118 513860 62186 513916
rect 62242 513860 62310 513916
rect 62366 513860 62434 513916
rect 62490 513860 62558 513916
rect 62614 513860 62682 513916
rect 62738 513860 62806 513916
rect 62862 513860 62930 513916
rect 62986 513860 63054 513916
rect 63110 513860 63178 513916
rect 63234 513860 63302 513916
rect 63358 513860 63426 513916
rect 63482 513860 63550 513916
rect 63606 513860 63674 513916
rect 63730 513860 63798 513916
rect 63854 513860 63922 513916
rect 63978 513860 64046 513916
rect 64102 513860 64170 513916
rect 64226 513860 64294 513916
rect 64350 513860 64418 513916
rect 64474 513860 64542 513916
rect 64598 513860 64666 513916
rect 64722 513860 64790 513916
rect 64846 513860 64914 513916
rect 64970 513860 65038 513916
rect 65094 513860 65162 513916
rect 65218 513860 65286 513916
rect 65342 513860 65410 513916
rect 65466 513860 65534 513916
rect 65590 513860 65658 513916
rect 65714 513860 65782 513916
rect 65838 513860 65906 513916
rect 65962 513860 66030 513916
rect 66086 513860 66154 513916
rect 66210 513860 66278 513916
rect 66334 513860 66402 513916
rect 66458 513860 597980 513916
rect -1916 513826 597980 513860
rect -1916 508435 597980 508446
rect -1916 508379 90112 508435
rect 90168 508379 90236 508435
rect 90292 508379 90360 508435
rect 90416 508379 90484 508435
rect 90540 508379 90608 508435
rect 90664 508379 90732 508435
rect 90788 508379 90856 508435
rect 90912 508379 90980 508435
rect 91036 508379 91104 508435
rect 91160 508379 91228 508435
rect 91284 508379 91352 508435
rect 91408 508379 91476 508435
rect 91532 508379 91600 508435
rect 91656 508379 91724 508435
rect 91780 508379 91848 508435
rect 91904 508379 91972 508435
rect 92028 508379 92096 508435
rect 92152 508379 92220 508435
rect 92276 508379 92344 508435
rect 92400 508379 92468 508435
rect 92524 508379 92592 508435
rect 92648 508379 92716 508435
rect 92772 508379 92840 508435
rect 92896 508379 92964 508435
rect 93020 508379 93088 508435
rect 93144 508379 93212 508435
rect 93268 508379 93336 508435
rect 93392 508379 93460 508435
rect 93516 508379 93584 508435
rect 93640 508379 93708 508435
rect 93764 508379 93832 508435
rect 93888 508379 93956 508435
rect 94012 508379 94080 508435
rect 94136 508379 94204 508435
rect 94260 508379 94328 508435
rect 94384 508379 94452 508435
rect 94508 508379 94576 508435
rect 94632 508379 94700 508435
rect 94756 508379 94824 508435
rect 94880 508379 94948 508435
rect 95004 508379 95072 508435
rect 95128 508379 95196 508435
rect 95252 508379 95320 508435
rect 95376 508379 95444 508435
rect 95500 508379 95568 508435
rect 95624 508379 95692 508435
rect 95748 508379 95816 508435
rect 95872 508379 95940 508435
rect 95996 508379 96064 508435
rect 96120 508379 96188 508435
rect 96244 508379 96312 508435
rect 96368 508379 96436 508435
rect 96492 508379 96560 508435
rect 96616 508379 96684 508435
rect 96740 508379 96808 508435
rect 96864 508379 96932 508435
rect 96988 508379 97056 508435
rect 97112 508379 97180 508435
rect 97236 508379 97304 508435
rect 97360 508379 97428 508435
rect 97484 508379 97552 508435
rect 97608 508379 97676 508435
rect 97732 508379 97800 508435
rect 97856 508379 97924 508435
rect 97980 508379 98048 508435
rect 98104 508379 98172 508435
rect 98228 508379 98296 508435
rect 98352 508379 98420 508435
rect 98476 508379 98544 508435
rect 98600 508379 98668 508435
rect 98724 508379 98792 508435
rect 98848 508379 98916 508435
rect 98972 508379 99040 508435
rect 99096 508379 99164 508435
rect 99220 508379 99288 508435
rect 99344 508379 99412 508435
rect 99468 508379 99536 508435
rect 99592 508379 99660 508435
rect 99716 508379 99784 508435
rect 99840 508379 99908 508435
rect 99964 508379 100032 508435
rect 100088 508379 597980 508435
rect -1916 508350 597980 508379
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508311 159114 508350
rect 36662 508294 90112 508311
rect -1916 508255 90112 508294
rect 90168 508255 90236 508311
rect 90292 508255 90360 508311
rect 90416 508255 90484 508311
rect 90540 508255 90608 508311
rect 90664 508255 90732 508311
rect 90788 508255 90856 508311
rect 90912 508255 90980 508311
rect 91036 508255 91104 508311
rect 91160 508255 91228 508311
rect 91284 508255 91352 508311
rect 91408 508255 91476 508311
rect 91532 508255 91600 508311
rect 91656 508255 91724 508311
rect 91780 508255 91848 508311
rect 91904 508255 91972 508311
rect 92028 508255 92096 508311
rect 92152 508255 92220 508311
rect 92276 508255 92344 508311
rect 92400 508255 92468 508311
rect 92524 508255 92592 508311
rect 92648 508255 92716 508311
rect 92772 508255 92840 508311
rect 92896 508255 92964 508311
rect 93020 508255 93088 508311
rect 93144 508255 93212 508311
rect 93268 508255 93336 508311
rect 93392 508255 93460 508311
rect 93516 508255 93584 508311
rect 93640 508255 93708 508311
rect 93764 508255 93832 508311
rect 93888 508255 93956 508311
rect 94012 508255 94080 508311
rect 94136 508255 94204 508311
rect 94260 508255 94328 508311
rect 94384 508255 94452 508311
rect 94508 508255 94576 508311
rect 94632 508255 94700 508311
rect 94756 508255 94824 508311
rect 94880 508255 94948 508311
rect 95004 508255 95072 508311
rect 95128 508255 95196 508311
rect 95252 508255 95320 508311
rect 95376 508255 95444 508311
rect 95500 508255 95568 508311
rect 95624 508255 95692 508311
rect 95748 508255 95816 508311
rect 95872 508255 95940 508311
rect 95996 508255 96064 508311
rect 96120 508255 96188 508311
rect 96244 508255 96312 508311
rect 96368 508255 96436 508311
rect 96492 508255 96560 508311
rect 96616 508255 96684 508311
rect 96740 508255 96808 508311
rect 96864 508255 96932 508311
rect 96988 508255 97056 508311
rect 97112 508255 97180 508311
rect 97236 508255 97304 508311
rect 97360 508255 97428 508311
rect 97484 508255 97552 508311
rect 97608 508255 97676 508311
rect 97732 508255 97800 508311
rect 97856 508255 97924 508311
rect 97980 508255 98048 508311
rect 98104 508255 98172 508311
rect 98228 508255 98296 508311
rect 98352 508255 98420 508311
rect 98476 508255 98544 508311
rect 98600 508255 98668 508311
rect 98724 508255 98792 508311
rect 98848 508255 98916 508311
rect 98972 508255 99040 508311
rect 99096 508255 99164 508311
rect 99220 508255 99288 508311
rect 99344 508255 99412 508311
rect 99468 508255 99536 508311
rect 99592 508255 99660 508311
rect 99716 508255 99784 508311
rect 99840 508255 99908 508311
rect 99964 508255 100032 508311
rect 100088 508294 159114 508311
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 194518 508350
rect 194574 508294 194642 508350
rect 194698 508294 225238 508350
rect 225294 508294 225362 508350
rect 225418 508294 255958 508350
rect 256014 508294 256082 508350
rect 256138 508294 286678 508350
rect 286734 508294 286802 508350
rect 286858 508294 317398 508350
rect 317454 508294 317522 508350
rect 317578 508294 348118 508350
rect 348174 508294 348242 508350
rect 348298 508294 378838 508350
rect 378894 508294 378962 508350
rect 379018 508294 409558 508350
rect 409614 508294 409682 508350
rect 409738 508294 440278 508350
rect 440334 508294 440402 508350
rect 440458 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 470998 508350
rect 471054 508294 471122 508350
rect 471178 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 501718 508350
rect 501774 508294 501842 508350
rect 501898 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect 100088 508255 597980 508294
rect -1916 508226 597980 508255
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508187 159114 508226
rect 36662 508170 90112 508187
rect -1916 508131 90112 508170
rect 90168 508131 90236 508187
rect 90292 508131 90360 508187
rect 90416 508131 90484 508187
rect 90540 508131 90608 508187
rect 90664 508131 90732 508187
rect 90788 508131 90856 508187
rect 90912 508131 90980 508187
rect 91036 508131 91104 508187
rect 91160 508131 91228 508187
rect 91284 508131 91352 508187
rect 91408 508131 91476 508187
rect 91532 508131 91600 508187
rect 91656 508131 91724 508187
rect 91780 508131 91848 508187
rect 91904 508131 91972 508187
rect 92028 508131 92096 508187
rect 92152 508131 92220 508187
rect 92276 508131 92344 508187
rect 92400 508131 92468 508187
rect 92524 508131 92592 508187
rect 92648 508131 92716 508187
rect 92772 508131 92840 508187
rect 92896 508131 92964 508187
rect 93020 508131 93088 508187
rect 93144 508131 93212 508187
rect 93268 508131 93336 508187
rect 93392 508131 93460 508187
rect 93516 508131 93584 508187
rect 93640 508131 93708 508187
rect 93764 508131 93832 508187
rect 93888 508131 93956 508187
rect 94012 508131 94080 508187
rect 94136 508131 94204 508187
rect 94260 508131 94328 508187
rect 94384 508131 94452 508187
rect 94508 508131 94576 508187
rect 94632 508131 94700 508187
rect 94756 508131 94824 508187
rect 94880 508131 94948 508187
rect 95004 508131 95072 508187
rect 95128 508131 95196 508187
rect 95252 508131 95320 508187
rect 95376 508131 95444 508187
rect 95500 508131 95568 508187
rect 95624 508131 95692 508187
rect 95748 508131 95816 508187
rect 95872 508131 95940 508187
rect 95996 508131 96064 508187
rect 96120 508131 96188 508187
rect 96244 508131 96312 508187
rect 96368 508131 96436 508187
rect 96492 508131 96560 508187
rect 96616 508131 96684 508187
rect 96740 508131 96808 508187
rect 96864 508131 96932 508187
rect 96988 508131 97056 508187
rect 97112 508131 97180 508187
rect 97236 508131 97304 508187
rect 97360 508131 97428 508187
rect 97484 508131 97552 508187
rect 97608 508131 97676 508187
rect 97732 508131 97800 508187
rect 97856 508131 97924 508187
rect 97980 508131 98048 508187
rect 98104 508131 98172 508187
rect 98228 508131 98296 508187
rect 98352 508131 98420 508187
rect 98476 508131 98544 508187
rect 98600 508131 98668 508187
rect 98724 508131 98792 508187
rect 98848 508131 98916 508187
rect 98972 508131 99040 508187
rect 99096 508131 99164 508187
rect 99220 508131 99288 508187
rect 99344 508131 99412 508187
rect 99468 508131 99536 508187
rect 99592 508131 99660 508187
rect 99716 508131 99784 508187
rect 99840 508131 99908 508187
rect 99964 508131 100032 508187
rect 100088 508170 159114 508187
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 194518 508226
rect 194574 508170 194642 508226
rect 194698 508170 225238 508226
rect 225294 508170 225362 508226
rect 225418 508170 255958 508226
rect 256014 508170 256082 508226
rect 256138 508170 286678 508226
rect 286734 508170 286802 508226
rect 286858 508170 317398 508226
rect 317454 508170 317522 508226
rect 317578 508170 348118 508226
rect 348174 508170 348242 508226
rect 348298 508170 378838 508226
rect 378894 508170 378962 508226
rect 379018 508170 409558 508226
rect 409614 508170 409682 508226
rect 409738 508170 440278 508226
rect 440334 508170 440402 508226
rect 440458 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 470998 508226
rect 471054 508170 471122 508226
rect 471178 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 501718 508226
rect 501774 508170 501842 508226
rect 501898 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect 100088 508131 597980 508170
rect -1916 508102 597980 508131
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 194518 508102
rect 194574 508046 194642 508102
rect 194698 508046 225238 508102
rect 225294 508046 225362 508102
rect 225418 508046 255958 508102
rect 256014 508046 256082 508102
rect 256138 508046 286678 508102
rect 286734 508046 286802 508102
rect 286858 508046 317398 508102
rect 317454 508046 317522 508102
rect 317578 508046 348118 508102
rect 348174 508046 348242 508102
rect 348298 508046 378838 508102
rect 378894 508046 378962 508102
rect 379018 508046 409558 508102
rect 409614 508046 409682 508102
rect 409738 508046 440278 508102
rect 440334 508046 440402 508102
rect 440458 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 470998 508102
rect 471054 508046 471122 508102
rect 471178 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 501718 508102
rect 501774 508046 501842 508102
rect 501898 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 194518 507978
rect 194574 507922 194642 507978
rect 194698 507922 225238 507978
rect 225294 507922 225362 507978
rect 225418 507922 255958 507978
rect 256014 507922 256082 507978
rect 256138 507922 286678 507978
rect 286734 507922 286802 507978
rect 286858 507922 317398 507978
rect 317454 507922 317522 507978
rect 317578 507922 348118 507978
rect 348174 507922 348242 507978
rect 348298 507922 378838 507978
rect 378894 507922 378962 507978
rect 379018 507922 409558 507978
rect 409614 507922 409682 507978
rect 409738 507922 440278 507978
rect 440334 507922 440402 507978
rect 440458 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 470998 507978
rect 471054 507922 471122 507978
rect 471178 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 501718 507978
rect 501774 507922 501842 507978
rect 501898 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 209878 496350
rect 209934 496294 210002 496350
rect 210058 496294 240598 496350
rect 240654 496294 240722 496350
rect 240778 496294 271318 496350
rect 271374 496294 271442 496350
rect 271498 496294 302038 496350
rect 302094 496294 302162 496350
rect 302218 496294 332758 496350
rect 332814 496294 332882 496350
rect 332938 496294 363478 496350
rect 363534 496294 363602 496350
rect 363658 496294 394198 496350
rect 394254 496294 394322 496350
rect 394378 496294 424918 496350
rect 424974 496294 425042 496350
rect 425098 496294 455638 496350
rect 455694 496294 455762 496350
rect 455818 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 486358 496350
rect 486414 496294 486482 496350
rect 486538 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 517078 496350
rect 517134 496294 517202 496350
rect 517258 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496212 162834 496226
rect 40382 496170 63430 496212
rect -1916 496156 63430 496170
rect 63486 496156 63554 496212
rect 63610 496156 63678 496212
rect 63734 496156 63802 496212
rect 63858 496156 63926 496212
rect 63982 496156 64050 496212
rect 64106 496156 64174 496212
rect 64230 496156 64298 496212
rect 64354 496156 64422 496212
rect 64478 496156 64546 496212
rect 64602 496156 64670 496212
rect 64726 496156 64794 496212
rect 64850 496156 64918 496212
rect 64974 496156 65042 496212
rect 65098 496156 65166 496212
rect 65222 496156 65290 496212
rect 65346 496156 65414 496212
rect 65470 496156 65538 496212
rect 65594 496156 65662 496212
rect 65718 496156 65786 496212
rect 65842 496156 65910 496212
rect 65966 496156 66034 496212
rect 66090 496156 66158 496212
rect 66214 496156 66282 496212
rect 66338 496156 66406 496212
rect 66462 496156 66530 496212
rect 66586 496156 66654 496212
rect 66710 496156 66778 496212
rect 66834 496156 66902 496212
rect 66958 496156 67026 496212
rect 67082 496156 67150 496212
rect 67206 496156 67274 496212
rect 67330 496156 67398 496212
rect 67454 496156 67522 496212
rect 67578 496156 67646 496212
rect 67702 496156 67770 496212
rect 67826 496156 67894 496212
rect 67950 496156 68018 496212
rect 68074 496156 68142 496212
rect 68198 496156 68266 496212
rect 68322 496156 68390 496212
rect 68446 496156 68514 496212
rect 68570 496156 68638 496212
rect 68694 496156 68762 496212
rect 68818 496156 68886 496212
rect 68942 496156 69010 496212
rect 69066 496156 69134 496212
rect 69190 496156 69258 496212
rect 69314 496156 69382 496212
rect 69438 496156 69506 496212
rect 69562 496156 69630 496212
rect 69686 496156 69754 496212
rect 69810 496156 69878 496212
rect 69934 496156 70002 496212
rect 70058 496156 70126 496212
rect 70182 496156 70250 496212
rect 70306 496156 70374 496212
rect 70430 496170 162834 496212
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 209878 496226
rect 209934 496170 210002 496226
rect 210058 496170 240598 496226
rect 240654 496170 240722 496226
rect 240778 496170 271318 496226
rect 271374 496170 271442 496226
rect 271498 496170 302038 496226
rect 302094 496170 302162 496226
rect 302218 496170 332758 496226
rect 332814 496170 332882 496226
rect 332938 496170 363478 496226
rect 363534 496170 363602 496226
rect 363658 496170 394198 496226
rect 394254 496170 394322 496226
rect 394378 496170 424918 496226
rect 424974 496170 425042 496226
rect 425098 496170 455638 496226
rect 455694 496170 455762 496226
rect 455818 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 486358 496226
rect 486414 496170 486482 496226
rect 486538 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 517078 496226
rect 517134 496170 517202 496226
rect 517258 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 70430 496156 597980 496170
rect -1916 496102 597980 496156
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496088 162834 496102
rect 40382 496046 63430 496088
rect -1916 496032 63430 496046
rect 63486 496032 63554 496088
rect 63610 496032 63678 496088
rect 63734 496032 63802 496088
rect 63858 496032 63926 496088
rect 63982 496032 64050 496088
rect 64106 496032 64174 496088
rect 64230 496032 64298 496088
rect 64354 496032 64422 496088
rect 64478 496032 64546 496088
rect 64602 496032 64670 496088
rect 64726 496032 64794 496088
rect 64850 496032 64918 496088
rect 64974 496032 65042 496088
rect 65098 496032 65166 496088
rect 65222 496032 65290 496088
rect 65346 496032 65414 496088
rect 65470 496032 65538 496088
rect 65594 496032 65662 496088
rect 65718 496032 65786 496088
rect 65842 496032 65910 496088
rect 65966 496032 66034 496088
rect 66090 496032 66158 496088
rect 66214 496032 66282 496088
rect 66338 496032 66406 496088
rect 66462 496032 66530 496088
rect 66586 496032 66654 496088
rect 66710 496032 66778 496088
rect 66834 496032 66902 496088
rect 66958 496032 67026 496088
rect 67082 496032 67150 496088
rect 67206 496032 67274 496088
rect 67330 496032 67398 496088
rect 67454 496032 67522 496088
rect 67578 496032 67646 496088
rect 67702 496032 67770 496088
rect 67826 496032 67894 496088
rect 67950 496032 68018 496088
rect 68074 496032 68142 496088
rect 68198 496032 68266 496088
rect 68322 496032 68390 496088
rect 68446 496032 68514 496088
rect 68570 496032 68638 496088
rect 68694 496032 68762 496088
rect 68818 496032 68886 496088
rect 68942 496032 69010 496088
rect 69066 496032 69134 496088
rect 69190 496032 69258 496088
rect 69314 496032 69382 496088
rect 69438 496032 69506 496088
rect 69562 496032 69630 496088
rect 69686 496032 69754 496088
rect 69810 496032 69878 496088
rect 69934 496032 70002 496088
rect 70058 496032 70126 496088
rect 70182 496032 70250 496088
rect 70306 496032 70374 496088
rect 70430 496046 162834 496088
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 209878 496102
rect 209934 496046 210002 496102
rect 210058 496046 240598 496102
rect 240654 496046 240722 496102
rect 240778 496046 271318 496102
rect 271374 496046 271442 496102
rect 271498 496046 302038 496102
rect 302094 496046 302162 496102
rect 302218 496046 332758 496102
rect 332814 496046 332882 496102
rect 332938 496046 363478 496102
rect 363534 496046 363602 496102
rect 363658 496046 394198 496102
rect 394254 496046 394322 496102
rect 394378 496046 424918 496102
rect 424974 496046 425042 496102
rect 425098 496046 455638 496102
rect 455694 496046 455762 496102
rect 455818 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 486358 496102
rect 486414 496046 486482 496102
rect 486538 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 517078 496102
rect 517134 496046 517202 496102
rect 517258 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 70430 496032 597980 496046
rect -1916 495978 597980 496032
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495964 162834 495978
rect 40382 495922 63430 495964
rect -1916 495908 63430 495922
rect 63486 495908 63554 495964
rect 63610 495908 63678 495964
rect 63734 495908 63802 495964
rect 63858 495908 63926 495964
rect 63982 495908 64050 495964
rect 64106 495908 64174 495964
rect 64230 495908 64298 495964
rect 64354 495908 64422 495964
rect 64478 495908 64546 495964
rect 64602 495908 64670 495964
rect 64726 495908 64794 495964
rect 64850 495908 64918 495964
rect 64974 495908 65042 495964
rect 65098 495908 65166 495964
rect 65222 495908 65290 495964
rect 65346 495908 65414 495964
rect 65470 495908 65538 495964
rect 65594 495908 65662 495964
rect 65718 495908 65786 495964
rect 65842 495908 65910 495964
rect 65966 495908 66034 495964
rect 66090 495908 66158 495964
rect 66214 495908 66282 495964
rect 66338 495908 66406 495964
rect 66462 495908 66530 495964
rect 66586 495908 66654 495964
rect 66710 495908 66778 495964
rect 66834 495908 66902 495964
rect 66958 495908 67026 495964
rect 67082 495908 67150 495964
rect 67206 495908 67274 495964
rect 67330 495908 67398 495964
rect 67454 495908 67522 495964
rect 67578 495908 67646 495964
rect 67702 495908 67770 495964
rect 67826 495908 67894 495964
rect 67950 495908 68018 495964
rect 68074 495908 68142 495964
rect 68198 495908 68266 495964
rect 68322 495908 68390 495964
rect 68446 495908 68514 495964
rect 68570 495908 68638 495964
rect 68694 495908 68762 495964
rect 68818 495908 68886 495964
rect 68942 495908 69010 495964
rect 69066 495908 69134 495964
rect 69190 495908 69258 495964
rect 69314 495908 69382 495964
rect 69438 495908 69506 495964
rect 69562 495908 69630 495964
rect 69686 495908 69754 495964
rect 69810 495908 69878 495964
rect 69934 495908 70002 495964
rect 70058 495908 70126 495964
rect 70182 495908 70250 495964
rect 70306 495908 70374 495964
rect 70430 495922 162834 495964
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 209878 495978
rect 209934 495922 210002 495978
rect 210058 495922 240598 495978
rect 240654 495922 240722 495978
rect 240778 495922 271318 495978
rect 271374 495922 271442 495978
rect 271498 495922 302038 495978
rect 302094 495922 302162 495978
rect 302218 495922 332758 495978
rect 332814 495922 332882 495978
rect 332938 495922 363478 495978
rect 363534 495922 363602 495978
rect 363658 495922 394198 495978
rect 394254 495922 394322 495978
rect 394378 495922 424918 495978
rect 424974 495922 425042 495978
rect 425098 495922 455638 495978
rect 455694 495922 455762 495978
rect 455818 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 486358 495978
rect 486414 495922 486482 495978
rect 486538 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 517078 495978
rect 517134 495922 517202 495978
rect 517258 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 70430 495908 597980 495922
rect -1916 495826 597980 495908
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 194518 490350
rect 194574 490294 194642 490350
rect 194698 490294 225238 490350
rect 225294 490294 225362 490350
rect 225418 490294 255958 490350
rect 256014 490294 256082 490350
rect 256138 490294 286678 490350
rect 286734 490294 286802 490350
rect 286858 490294 317398 490350
rect 317454 490294 317522 490350
rect 317578 490294 348118 490350
rect 348174 490294 348242 490350
rect 348298 490294 378838 490350
rect 378894 490294 378962 490350
rect 379018 490294 409558 490350
rect 409614 490294 409682 490350
rect 409738 490294 440278 490350
rect 440334 490294 440402 490350
rect 440458 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 470998 490350
rect 471054 490294 471122 490350
rect 471178 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 501718 490350
rect 501774 490294 501842 490350
rect 501898 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490272 597980 490294
rect -1916 490226 85236 490272
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490216 85236 490226
rect 85292 490216 85360 490272
rect 85416 490216 85484 490272
rect 85540 490216 85608 490272
rect 85664 490216 85732 490272
rect 85788 490216 85856 490272
rect 85912 490216 85980 490272
rect 86036 490216 86104 490272
rect 86160 490216 86228 490272
rect 86284 490216 86352 490272
rect 86408 490216 86476 490272
rect 86532 490216 86600 490272
rect 86656 490216 86724 490272
rect 86780 490216 86848 490272
rect 86904 490216 86972 490272
rect 87028 490216 87096 490272
rect 87152 490216 87220 490272
rect 87276 490216 87344 490272
rect 87400 490216 87468 490272
rect 87524 490216 87592 490272
rect 87648 490216 87716 490272
rect 87772 490216 87840 490272
rect 87896 490216 87964 490272
rect 88020 490216 88088 490272
rect 88144 490216 88212 490272
rect 88268 490216 88336 490272
rect 88392 490216 88460 490272
rect 88516 490216 88584 490272
rect 88640 490216 88708 490272
rect 88764 490226 597980 490272
rect 88764 490216 159114 490226
rect 36662 490170 159114 490216
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 194518 490226
rect 194574 490170 194642 490226
rect 194698 490170 225238 490226
rect 225294 490170 225362 490226
rect 225418 490170 255958 490226
rect 256014 490170 256082 490226
rect 256138 490170 286678 490226
rect 286734 490170 286802 490226
rect 286858 490170 317398 490226
rect 317454 490170 317522 490226
rect 317578 490170 348118 490226
rect 348174 490170 348242 490226
rect 348298 490170 378838 490226
rect 378894 490170 378962 490226
rect 379018 490170 409558 490226
rect 409614 490170 409682 490226
rect 409738 490170 440278 490226
rect 440334 490170 440402 490226
rect 440458 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 470998 490226
rect 471054 490170 471122 490226
rect 471178 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 501718 490226
rect 501774 490170 501842 490226
rect 501898 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490148 597980 490170
rect -1916 490102 85236 490148
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490092 85236 490102
rect 85292 490092 85360 490148
rect 85416 490092 85484 490148
rect 85540 490092 85608 490148
rect 85664 490092 85732 490148
rect 85788 490092 85856 490148
rect 85912 490092 85980 490148
rect 86036 490092 86104 490148
rect 86160 490092 86228 490148
rect 86284 490092 86352 490148
rect 86408 490092 86476 490148
rect 86532 490092 86600 490148
rect 86656 490092 86724 490148
rect 86780 490092 86848 490148
rect 86904 490092 86972 490148
rect 87028 490092 87096 490148
rect 87152 490092 87220 490148
rect 87276 490092 87344 490148
rect 87400 490092 87468 490148
rect 87524 490092 87592 490148
rect 87648 490092 87716 490148
rect 87772 490092 87840 490148
rect 87896 490092 87964 490148
rect 88020 490092 88088 490148
rect 88144 490092 88212 490148
rect 88268 490092 88336 490148
rect 88392 490092 88460 490148
rect 88516 490092 88584 490148
rect 88640 490092 88708 490148
rect 88764 490102 597980 490148
rect 88764 490092 159114 490102
rect 36662 490046 159114 490092
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 194518 490102
rect 194574 490046 194642 490102
rect 194698 490046 225238 490102
rect 225294 490046 225362 490102
rect 225418 490046 255958 490102
rect 256014 490046 256082 490102
rect 256138 490046 286678 490102
rect 286734 490046 286802 490102
rect 286858 490046 317398 490102
rect 317454 490046 317522 490102
rect 317578 490046 348118 490102
rect 348174 490046 348242 490102
rect 348298 490046 378838 490102
rect 378894 490046 378962 490102
rect 379018 490046 409558 490102
rect 409614 490046 409682 490102
rect 409738 490046 440278 490102
rect 440334 490046 440402 490102
rect 440458 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 470998 490102
rect 471054 490046 471122 490102
rect 471178 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 501718 490102
rect 501774 490046 501842 490102
rect 501898 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 490024 597980 490046
rect -1916 489978 85236 490024
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489968 85236 489978
rect 85292 489968 85360 490024
rect 85416 489968 85484 490024
rect 85540 489968 85608 490024
rect 85664 489968 85732 490024
rect 85788 489968 85856 490024
rect 85912 489968 85980 490024
rect 86036 489968 86104 490024
rect 86160 489968 86228 490024
rect 86284 489968 86352 490024
rect 86408 489968 86476 490024
rect 86532 489968 86600 490024
rect 86656 489968 86724 490024
rect 86780 489968 86848 490024
rect 86904 489968 86972 490024
rect 87028 489968 87096 490024
rect 87152 489968 87220 490024
rect 87276 489968 87344 490024
rect 87400 489968 87468 490024
rect 87524 489968 87592 490024
rect 87648 489968 87716 490024
rect 87772 489968 87840 490024
rect 87896 489968 87964 490024
rect 88020 489968 88088 490024
rect 88144 489968 88212 490024
rect 88268 489968 88336 490024
rect 88392 489968 88460 490024
rect 88516 489968 88584 490024
rect 88640 489968 88708 490024
rect 88764 489978 597980 490024
rect 88764 489968 159114 489978
rect 36662 489922 159114 489968
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 194518 489978
rect 194574 489922 194642 489978
rect 194698 489922 225238 489978
rect 225294 489922 225362 489978
rect 225418 489922 255958 489978
rect 256014 489922 256082 489978
rect 256138 489922 286678 489978
rect 286734 489922 286802 489978
rect 286858 489922 317398 489978
rect 317454 489922 317522 489978
rect 317578 489922 348118 489978
rect 348174 489922 348242 489978
rect 348298 489922 378838 489978
rect 378894 489922 378962 489978
rect 379018 489922 409558 489978
rect 409614 489922 409682 489978
rect 409738 489922 440278 489978
rect 440334 489922 440402 489978
rect 440458 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 470998 489978
rect 471054 489922 471122 489978
rect 471178 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 501718 489978
rect 501774 489922 501842 489978
rect 501898 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478358 597980 478446
rect -1916 478350 80936 478358
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478302 80936 478350
rect 80992 478302 81060 478358
rect 81116 478302 81184 478358
rect 81240 478302 81308 478358
rect 81364 478350 597980 478358
rect 81364 478302 132114 478350
rect 71102 478294 132114 478302
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 209878 478350
rect 209934 478294 210002 478350
rect 210058 478294 240598 478350
rect 240654 478294 240722 478350
rect 240778 478294 271318 478350
rect 271374 478294 271442 478350
rect 271498 478294 302038 478350
rect 302094 478294 302162 478350
rect 302218 478294 332758 478350
rect 332814 478294 332882 478350
rect 332938 478294 363478 478350
rect 363534 478294 363602 478350
rect 363658 478294 394198 478350
rect 394254 478294 394322 478350
rect 394378 478294 424918 478350
rect 424974 478294 425042 478350
rect 425098 478294 455638 478350
rect 455694 478294 455762 478350
rect 455818 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 486358 478350
rect 486414 478294 486482 478350
rect 486538 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 517078 478350
rect 517134 478294 517202 478350
rect 517258 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 209878 478226
rect 209934 478170 210002 478226
rect 210058 478170 240598 478226
rect 240654 478170 240722 478226
rect 240778 478170 271318 478226
rect 271374 478170 271442 478226
rect 271498 478170 302038 478226
rect 302094 478170 302162 478226
rect 302218 478170 332758 478226
rect 332814 478170 332882 478226
rect 332938 478170 363478 478226
rect 363534 478170 363602 478226
rect 363658 478170 394198 478226
rect 394254 478170 394322 478226
rect 394378 478170 424918 478226
rect 424974 478170 425042 478226
rect 425098 478170 455638 478226
rect 455694 478170 455762 478226
rect 455818 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 486358 478226
rect 486414 478170 486482 478226
rect 486538 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 517078 478226
rect 517134 478170 517202 478226
rect 517258 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 209878 478102
rect 209934 478046 210002 478102
rect 210058 478046 240598 478102
rect 240654 478046 240722 478102
rect 240778 478046 271318 478102
rect 271374 478046 271442 478102
rect 271498 478046 302038 478102
rect 302094 478046 302162 478102
rect 302218 478046 332758 478102
rect 332814 478046 332882 478102
rect 332938 478046 363478 478102
rect 363534 478046 363602 478102
rect 363658 478046 394198 478102
rect 394254 478046 394322 478102
rect 394378 478046 424918 478102
rect 424974 478046 425042 478102
rect 425098 478046 455638 478102
rect 455694 478046 455762 478102
rect 455818 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 486358 478102
rect 486414 478046 486482 478102
rect 486538 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 517078 478102
rect 517134 478046 517202 478102
rect 517258 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 209878 477978
rect 209934 477922 210002 477978
rect 210058 477922 240598 477978
rect 240654 477922 240722 477978
rect 240778 477922 271318 477978
rect 271374 477922 271442 477978
rect 271498 477922 302038 477978
rect 302094 477922 302162 477978
rect 302218 477922 332758 477978
rect 332814 477922 332882 477978
rect 332938 477922 363478 477978
rect 363534 477922 363602 477978
rect 363658 477922 394198 477978
rect 394254 477922 394322 477978
rect 394378 477922 424918 477978
rect 424974 477922 425042 477978
rect 425098 477922 455638 477978
rect 455694 477922 455762 477978
rect 455818 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 486358 477978
rect 486414 477922 486482 477978
rect 486538 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 517078 477978
rect 517134 477922 517202 477978
rect 517258 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 194518 472350
rect 194574 472294 194642 472350
rect 194698 472294 225238 472350
rect 225294 472294 225362 472350
rect 225418 472294 255958 472350
rect 256014 472294 256082 472350
rect 256138 472294 286678 472350
rect 286734 472294 286802 472350
rect 286858 472294 317398 472350
rect 317454 472294 317522 472350
rect 317578 472294 348118 472350
rect 348174 472294 348242 472350
rect 348298 472294 378838 472350
rect 378894 472294 378962 472350
rect 379018 472294 409558 472350
rect 409614 472294 409682 472350
rect 409738 472294 440278 472350
rect 440334 472294 440402 472350
rect 440458 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 470998 472350
rect 471054 472294 471122 472350
rect 471178 472294 497034 472350
rect 497090 472294 497158 472350
rect 497214 472294 497282 472350
rect 497338 472294 497406 472350
rect 497462 472294 501718 472350
rect 501774 472294 501842 472350
rect 501898 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 194518 472226
rect 194574 472170 194642 472226
rect 194698 472170 225238 472226
rect 225294 472170 225362 472226
rect 225418 472170 255958 472226
rect 256014 472170 256082 472226
rect 256138 472170 286678 472226
rect 286734 472170 286802 472226
rect 286858 472170 317398 472226
rect 317454 472170 317522 472226
rect 317578 472170 348118 472226
rect 348174 472170 348242 472226
rect 348298 472170 378838 472226
rect 378894 472170 378962 472226
rect 379018 472170 409558 472226
rect 409614 472170 409682 472226
rect 409738 472170 440278 472226
rect 440334 472170 440402 472226
rect 440458 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 470998 472226
rect 471054 472170 471122 472226
rect 471178 472170 497034 472226
rect 497090 472170 497158 472226
rect 497214 472170 497282 472226
rect 497338 472170 497406 472226
rect 497462 472170 501718 472226
rect 501774 472170 501842 472226
rect 501898 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 194518 472102
rect 194574 472046 194642 472102
rect 194698 472046 225238 472102
rect 225294 472046 225362 472102
rect 225418 472046 255958 472102
rect 256014 472046 256082 472102
rect 256138 472046 286678 472102
rect 286734 472046 286802 472102
rect 286858 472046 317398 472102
rect 317454 472046 317522 472102
rect 317578 472046 348118 472102
rect 348174 472046 348242 472102
rect 348298 472046 378838 472102
rect 378894 472046 378962 472102
rect 379018 472046 409558 472102
rect 409614 472046 409682 472102
rect 409738 472046 440278 472102
rect 440334 472046 440402 472102
rect 440458 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 470998 472102
rect 471054 472046 471122 472102
rect 471178 472046 497034 472102
rect 497090 472046 497158 472102
rect 497214 472046 497282 472102
rect 497338 472046 497406 472102
rect 497462 472046 501718 472102
rect 501774 472046 501842 472102
rect 501898 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 194518 471978
rect 194574 471922 194642 471978
rect 194698 471922 225238 471978
rect 225294 471922 225362 471978
rect 225418 471922 255958 471978
rect 256014 471922 256082 471978
rect 256138 471922 286678 471978
rect 286734 471922 286802 471978
rect 286858 471922 317398 471978
rect 317454 471922 317522 471978
rect 317578 471922 348118 471978
rect 348174 471922 348242 471978
rect 348298 471922 378838 471978
rect 378894 471922 378962 471978
rect 379018 471922 409558 471978
rect 409614 471922 409682 471978
rect 409738 471922 440278 471978
rect 440334 471922 440402 471978
rect 440458 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 470998 471978
rect 471054 471922 471122 471978
rect 471178 471922 497034 471978
rect 497090 471922 497158 471978
rect 497214 471922 497282 471978
rect 497338 471922 497406 471978
rect 497462 471922 501718 471978
rect 501774 471922 501842 471978
rect 501898 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 209878 460350
rect 209934 460294 210002 460350
rect 210058 460294 240598 460350
rect 240654 460294 240722 460350
rect 240778 460294 271318 460350
rect 271374 460294 271442 460350
rect 271498 460294 302038 460350
rect 302094 460294 302162 460350
rect 302218 460294 332758 460350
rect 332814 460294 332882 460350
rect 332938 460294 363478 460350
rect 363534 460294 363602 460350
rect 363658 460294 394198 460350
rect 394254 460294 394322 460350
rect 394378 460294 424918 460350
rect 424974 460294 425042 460350
rect 425098 460294 455638 460350
rect 455694 460294 455762 460350
rect 455818 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 486358 460350
rect 486414 460294 486482 460350
rect 486538 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 517078 460350
rect 517134 460294 517202 460350
rect 517258 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 209878 460226
rect 209934 460170 210002 460226
rect 210058 460170 240598 460226
rect 240654 460170 240722 460226
rect 240778 460170 271318 460226
rect 271374 460170 271442 460226
rect 271498 460170 302038 460226
rect 302094 460170 302162 460226
rect 302218 460170 332758 460226
rect 332814 460170 332882 460226
rect 332938 460170 363478 460226
rect 363534 460170 363602 460226
rect 363658 460170 394198 460226
rect 394254 460170 394322 460226
rect 394378 460170 424918 460226
rect 424974 460170 425042 460226
rect 425098 460170 455638 460226
rect 455694 460170 455762 460226
rect 455818 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 486358 460226
rect 486414 460170 486482 460226
rect 486538 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 517078 460226
rect 517134 460170 517202 460226
rect 517258 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 209878 460102
rect 209934 460046 210002 460102
rect 210058 460046 240598 460102
rect 240654 460046 240722 460102
rect 240778 460046 271318 460102
rect 271374 460046 271442 460102
rect 271498 460046 302038 460102
rect 302094 460046 302162 460102
rect 302218 460046 332758 460102
rect 332814 460046 332882 460102
rect 332938 460046 363478 460102
rect 363534 460046 363602 460102
rect 363658 460046 394198 460102
rect 394254 460046 394322 460102
rect 394378 460046 424918 460102
rect 424974 460046 425042 460102
rect 425098 460046 455638 460102
rect 455694 460046 455762 460102
rect 455818 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 486358 460102
rect 486414 460046 486482 460102
rect 486538 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 517078 460102
rect 517134 460046 517202 460102
rect 517258 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 209878 459978
rect 209934 459922 210002 459978
rect 210058 459922 240598 459978
rect 240654 459922 240722 459978
rect 240778 459922 271318 459978
rect 271374 459922 271442 459978
rect 271498 459922 302038 459978
rect 302094 459922 302162 459978
rect 302218 459922 332758 459978
rect 332814 459922 332882 459978
rect 332938 459922 363478 459978
rect 363534 459922 363602 459978
rect 363658 459922 394198 459978
rect 394254 459922 394322 459978
rect 394378 459922 424918 459978
rect 424974 459922 425042 459978
rect 425098 459922 455638 459978
rect 455694 459922 455762 459978
rect 455818 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 486358 459978
rect 486414 459922 486482 459978
rect 486538 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 517078 459978
rect 517134 459922 517202 459978
rect 517258 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 194518 454350
rect 194574 454294 194642 454350
rect 194698 454294 225238 454350
rect 225294 454294 225362 454350
rect 225418 454294 255958 454350
rect 256014 454294 256082 454350
rect 256138 454294 286678 454350
rect 286734 454294 286802 454350
rect 286858 454294 317398 454350
rect 317454 454294 317522 454350
rect 317578 454294 348118 454350
rect 348174 454294 348242 454350
rect 348298 454294 378838 454350
rect 378894 454294 378962 454350
rect 379018 454294 409558 454350
rect 409614 454294 409682 454350
rect 409738 454294 440278 454350
rect 440334 454294 440402 454350
rect 440458 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 470998 454350
rect 471054 454294 471122 454350
rect 471178 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 501718 454350
rect 501774 454294 501842 454350
rect 501898 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 194518 454226
rect 194574 454170 194642 454226
rect 194698 454170 225238 454226
rect 225294 454170 225362 454226
rect 225418 454170 255958 454226
rect 256014 454170 256082 454226
rect 256138 454170 286678 454226
rect 286734 454170 286802 454226
rect 286858 454170 317398 454226
rect 317454 454170 317522 454226
rect 317578 454170 348118 454226
rect 348174 454170 348242 454226
rect 348298 454170 378838 454226
rect 378894 454170 378962 454226
rect 379018 454170 409558 454226
rect 409614 454170 409682 454226
rect 409738 454170 440278 454226
rect 440334 454170 440402 454226
rect 440458 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 470998 454226
rect 471054 454170 471122 454226
rect 471178 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 501718 454226
rect 501774 454170 501842 454226
rect 501898 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 194518 454102
rect 194574 454046 194642 454102
rect 194698 454046 225238 454102
rect 225294 454046 225362 454102
rect 225418 454046 255958 454102
rect 256014 454046 256082 454102
rect 256138 454046 286678 454102
rect 286734 454046 286802 454102
rect 286858 454046 317398 454102
rect 317454 454046 317522 454102
rect 317578 454046 348118 454102
rect 348174 454046 348242 454102
rect 348298 454046 378838 454102
rect 378894 454046 378962 454102
rect 379018 454046 409558 454102
rect 409614 454046 409682 454102
rect 409738 454046 440278 454102
rect 440334 454046 440402 454102
rect 440458 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 470998 454102
rect 471054 454046 471122 454102
rect 471178 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 501718 454102
rect 501774 454046 501842 454102
rect 501898 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 194518 453978
rect 194574 453922 194642 453978
rect 194698 453922 225238 453978
rect 225294 453922 225362 453978
rect 225418 453922 255958 453978
rect 256014 453922 256082 453978
rect 256138 453922 286678 453978
rect 286734 453922 286802 453978
rect 286858 453922 317398 453978
rect 317454 453922 317522 453978
rect 317578 453922 348118 453978
rect 348174 453922 348242 453978
rect 348298 453922 378838 453978
rect 378894 453922 378962 453978
rect 379018 453922 409558 453978
rect 409614 453922 409682 453978
rect 409738 453922 440278 453978
rect 440334 453922 440402 453978
rect 440458 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 470998 453978
rect 471054 453922 471122 453978
rect 471178 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 501718 453978
rect 501774 453922 501842 453978
rect 501898 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 209878 442350
rect 209934 442294 210002 442350
rect 210058 442294 240598 442350
rect 240654 442294 240722 442350
rect 240778 442294 271318 442350
rect 271374 442294 271442 442350
rect 271498 442294 302038 442350
rect 302094 442294 302162 442350
rect 302218 442294 332758 442350
rect 332814 442294 332882 442350
rect 332938 442294 363478 442350
rect 363534 442294 363602 442350
rect 363658 442294 394198 442350
rect 394254 442294 394322 442350
rect 394378 442294 424918 442350
rect 424974 442294 425042 442350
rect 425098 442294 455638 442350
rect 455694 442294 455762 442350
rect 455818 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 486358 442350
rect 486414 442294 486482 442350
rect 486538 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 517078 442350
rect 517134 442294 517202 442350
rect 517258 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 209878 442226
rect 209934 442170 210002 442226
rect 210058 442170 240598 442226
rect 240654 442170 240722 442226
rect 240778 442170 271318 442226
rect 271374 442170 271442 442226
rect 271498 442170 302038 442226
rect 302094 442170 302162 442226
rect 302218 442170 332758 442226
rect 332814 442170 332882 442226
rect 332938 442170 363478 442226
rect 363534 442170 363602 442226
rect 363658 442170 394198 442226
rect 394254 442170 394322 442226
rect 394378 442170 424918 442226
rect 424974 442170 425042 442226
rect 425098 442170 455638 442226
rect 455694 442170 455762 442226
rect 455818 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 486358 442226
rect 486414 442170 486482 442226
rect 486538 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 517078 442226
rect 517134 442170 517202 442226
rect 517258 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 209878 442102
rect 209934 442046 210002 442102
rect 210058 442046 240598 442102
rect 240654 442046 240722 442102
rect 240778 442046 271318 442102
rect 271374 442046 271442 442102
rect 271498 442046 302038 442102
rect 302094 442046 302162 442102
rect 302218 442046 332758 442102
rect 332814 442046 332882 442102
rect 332938 442046 363478 442102
rect 363534 442046 363602 442102
rect 363658 442046 394198 442102
rect 394254 442046 394322 442102
rect 394378 442046 424918 442102
rect 424974 442046 425042 442102
rect 425098 442046 455638 442102
rect 455694 442046 455762 442102
rect 455818 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 486358 442102
rect 486414 442046 486482 442102
rect 486538 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 517078 442102
rect 517134 442046 517202 442102
rect 517258 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 209878 441978
rect 209934 441922 210002 441978
rect 210058 441922 240598 441978
rect 240654 441922 240722 441978
rect 240778 441922 271318 441978
rect 271374 441922 271442 441978
rect 271498 441922 302038 441978
rect 302094 441922 302162 441978
rect 302218 441922 332758 441978
rect 332814 441922 332882 441978
rect 332938 441922 363478 441978
rect 363534 441922 363602 441978
rect 363658 441922 394198 441978
rect 394254 441922 394322 441978
rect 394378 441922 424918 441978
rect 424974 441922 425042 441978
rect 425098 441922 455638 441978
rect 455694 441922 455762 441978
rect 455818 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 486358 441978
rect 486414 441922 486482 441978
rect 486538 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 517078 441978
rect 517134 441922 517202 441978
rect 517258 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 194518 436350
rect 194574 436294 194642 436350
rect 194698 436294 225238 436350
rect 225294 436294 225362 436350
rect 225418 436294 255958 436350
rect 256014 436294 256082 436350
rect 256138 436294 286678 436350
rect 286734 436294 286802 436350
rect 286858 436294 317398 436350
rect 317454 436294 317522 436350
rect 317578 436294 348118 436350
rect 348174 436294 348242 436350
rect 348298 436294 378838 436350
rect 378894 436294 378962 436350
rect 379018 436294 409558 436350
rect 409614 436294 409682 436350
rect 409738 436294 440278 436350
rect 440334 436294 440402 436350
rect 440458 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 470998 436350
rect 471054 436294 471122 436350
rect 471178 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 501718 436350
rect 501774 436294 501842 436350
rect 501898 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 194518 436226
rect 194574 436170 194642 436226
rect 194698 436170 225238 436226
rect 225294 436170 225362 436226
rect 225418 436170 255958 436226
rect 256014 436170 256082 436226
rect 256138 436170 286678 436226
rect 286734 436170 286802 436226
rect 286858 436170 317398 436226
rect 317454 436170 317522 436226
rect 317578 436170 348118 436226
rect 348174 436170 348242 436226
rect 348298 436170 378838 436226
rect 378894 436170 378962 436226
rect 379018 436170 409558 436226
rect 409614 436170 409682 436226
rect 409738 436170 440278 436226
rect 440334 436170 440402 436226
rect 440458 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 470998 436226
rect 471054 436170 471122 436226
rect 471178 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 501718 436226
rect 501774 436170 501842 436226
rect 501898 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 194518 436102
rect 194574 436046 194642 436102
rect 194698 436046 225238 436102
rect 225294 436046 225362 436102
rect 225418 436046 255958 436102
rect 256014 436046 256082 436102
rect 256138 436046 286678 436102
rect 286734 436046 286802 436102
rect 286858 436046 317398 436102
rect 317454 436046 317522 436102
rect 317578 436046 348118 436102
rect 348174 436046 348242 436102
rect 348298 436046 378838 436102
rect 378894 436046 378962 436102
rect 379018 436046 409558 436102
rect 409614 436046 409682 436102
rect 409738 436046 440278 436102
rect 440334 436046 440402 436102
rect 440458 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 470998 436102
rect 471054 436046 471122 436102
rect 471178 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 501718 436102
rect 501774 436046 501842 436102
rect 501898 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 194518 435978
rect 194574 435922 194642 435978
rect 194698 435922 225238 435978
rect 225294 435922 225362 435978
rect 225418 435922 255958 435978
rect 256014 435922 256082 435978
rect 256138 435922 286678 435978
rect 286734 435922 286802 435978
rect 286858 435922 317398 435978
rect 317454 435922 317522 435978
rect 317578 435922 348118 435978
rect 348174 435922 348242 435978
rect 348298 435922 378838 435978
rect 378894 435922 378962 435978
rect 379018 435922 409558 435978
rect 409614 435922 409682 435978
rect 409738 435922 440278 435978
rect 440334 435922 440402 435978
rect 440458 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 470998 435978
rect 471054 435922 471122 435978
rect 471178 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 501718 435978
rect 501774 435922 501842 435978
rect 501898 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect 525796 428698 529300 428714
rect 525796 428642 529228 428698
rect 529284 428642 529300 428698
rect 525796 428626 529300 428642
rect 525796 428534 525884 428626
rect 445996 428518 525884 428534
rect 445996 428462 446012 428518
rect 446068 428462 525884 428518
rect 445996 428446 525884 428462
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 209878 424350
rect 209934 424294 210002 424350
rect 210058 424294 240598 424350
rect 240654 424294 240722 424350
rect 240778 424294 271318 424350
rect 271374 424294 271442 424350
rect 271498 424294 302038 424350
rect 302094 424294 302162 424350
rect 302218 424294 332758 424350
rect 332814 424294 332882 424350
rect 332938 424294 363478 424350
rect 363534 424294 363602 424350
rect 363658 424294 394198 424350
rect 394254 424294 394322 424350
rect 394378 424294 424918 424350
rect 424974 424294 425042 424350
rect 425098 424294 455638 424350
rect 455694 424294 455762 424350
rect 455818 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 486358 424350
rect 486414 424294 486482 424350
rect 486538 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 517078 424350
rect 517134 424294 517202 424350
rect 517258 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 209878 424226
rect 209934 424170 210002 424226
rect 210058 424170 240598 424226
rect 240654 424170 240722 424226
rect 240778 424170 271318 424226
rect 271374 424170 271442 424226
rect 271498 424170 302038 424226
rect 302094 424170 302162 424226
rect 302218 424170 332758 424226
rect 332814 424170 332882 424226
rect 332938 424170 363478 424226
rect 363534 424170 363602 424226
rect 363658 424170 394198 424226
rect 394254 424170 394322 424226
rect 394378 424170 424918 424226
rect 424974 424170 425042 424226
rect 425098 424170 455638 424226
rect 455694 424170 455762 424226
rect 455818 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 486358 424226
rect 486414 424170 486482 424226
rect 486538 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 517078 424226
rect 517134 424170 517202 424226
rect 517258 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 209878 424102
rect 209934 424046 210002 424102
rect 210058 424046 240598 424102
rect 240654 424046 240722 424102
rect 240778 424046 271318 424102
rect 271374 424046 271442 424102
rect 271498 424046 302038 424102
rect 302094 424046 302162 424102
rect 302218 424046 332758 424102
rect 332814 424046 332882 424102
rect 332938 424046 363478 424102
rect 363534 424046 363602 424102
rect 363658 424046 394198 424102
rect 394254 424046 394322 424102
rect 394378 424046 424918 424102
rect 424974 424046 425042 424102
rect 425098 424046 455638 424102
rect 455694 424046 455762 424102
rect 455818 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 486358 424102
rect 486414 424046 486482 424102
rect 486538 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 517078 424102
rect 517134 424046 517202 424102
rect 517258 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 209878 423978
rect 209934 423922 210002 423978
rect 210058 423922 240598 423978
rect 240654 423922 240722 423978
rect 240778 423922 271318 423978
rect 271374 423922 271442 423978
rect 271498 423922 302038 423978
rect 302094 423922 302162 423978
rect 302218 423922 332758 423978
rect 332814 423922 332882 423978
rect 332938 423922 363478 423978
rect 363534 423922 363602 423978
rect 363658 423922 394198 423978
rect 394254 423922 394322 423978
rect 394378 423922 424918 423978
rect 424974 423922 425042 423978
rect 425098 423922 455638 423978
rect 455694 423922 455762 423978
rect 455818 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 486358 423978
rect 486414 423922 486482 423978
rect 486538 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 517078 423978
rect 517134 423922 517202 423978
rect 517258 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 194518 418350
rect 194574 418294 194642 418350
rect 194698 418294 225238 418350
rect 225294 418294 225362 418350
rect 225418 418294 255958 418350
rect 256014 418294 256082 418350
rect 256138 418294 286678 418350
rect 286734 418294 286802 418350
rect 286858 418294 317398 418350
rect 317454 418294 317522 418350
rect 317578 418294 348118 418350
rect 348174 418294 348242 418350
rect 348298 418294 378838 418350
rect 378894 418294 378962 418350
rect 379018 418294 409558 418350
rect 409614 418294 409682 418350
rect 409738 418294 440278 418350
rect 440334 418294 440402 418350
rect 440458 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 470998 418350
rect 471054 418294 471122 418350
rect 471178 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 501718 418350
rect 501774 418294 501842 418350
rect 501898 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 194518 418226
rect 194574 418170 194642 418226
rect 194698 418170 225238 418226
rect 225294 418170 225362 418226
rect 225418 418170 255958 418226
rect 256014 418170 256082 418226
rect 256138 418170 286678 418226
rect 286734 418170 286802 418226
rect 286858 418170 317398 418226
rect 317454 418170 317522 418226
rect 317578 418170 348118 418226
rect 348174 418170 348242 418226
rect 348298 418170 378838 418226
rect 378894 418170 378962 418226
rect 379018 418170 409558 418226
rect 409614 418170 409682 418226
rect 409738 418170 440278 418226
rect 440334 418170 440402 418226
rect 440458 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 470998 418226
rect 471054 418170 471122 418226
rect 471178 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 501718 418226
rect 501774 418170 501842 418226
rect 501898 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 194518 418102
rect 194574 418046 194642 418102
rect 194698 418046 225238 418102
rect 225294 418046 225362 418102
rect 225418 418046 255958 418102
rect 256014 418046 256082 418102
rect 256138 418046 286678 418102
rect 286734 418046 286802 418102
rect 286858 418046 317398 418102
rect 317454 418046 317522 418102
rect 317578 418046 348118 418102
rect 348174 418046 348242 418102
rect 348298 418046 378838 418102
rect 378894 418046 378962 418102
rect 379018 418046 409558 418102
rect 409614 418046 409682 418102
rect 409738 418046 440278 418102
rect 440334 418046 440402 418102
rect 440458 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 470998 418102
rect 471054 418046 471122 418102
rect 471178 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 501718 418102
rect 501774 418046 501842 418102
rect 501898 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 194518 417978
rect 194574 417922 194642 417978
rect 194698 417922 225238 417978
rect 225294 417922 225362 417978
rect 225418 417922 255958 417978
rect 256014 417922 256082 417978
rect 256138 417922 286678 417978
rect 286734 417922 286802 417978
rect 286858 417922 317398 417978
rect 317454 417922 317522 417978
rect 317578 417922 348118 417978
rect 348174 417922 348242 417978
rect 348298 417922 378838 417978
rect 378894 417922 378962 417978
rect 379018 417922 409558 417978
rect 409614 417922 409682 417978
rect 409738 417922 440278 417978
rect 440334 417922 440402 417978
rect 440458 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 470998 417978
rect 471054 417922 471122 417978
rect 471178 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 501718 417978
rect 501774 417922 501842 417978
rect 501898 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect 4156 416818 83988 416834
rect 4156 416762 4172 416818
rect 4228 416762 83916 416818
rect 83972 416762 83988 416818
rect 4156 416746 83988 416762
rect 354380 409798 584740 409814
rect 354380 409742 354396 409798
rect 354452 409742 584668 409798
rect 584724 409742 584740 409798
rect 354380 409726 584740 409742
rect 357740 409618 590788 409634
rect 357740 409562 357756 409618
rect 357812 409562 590716 409618
rect 590772 409562 590788 409618
rect 357740 409546 590788 409562
rect 157036 409438 289844 409454
rect 157036 409382 157052 409438
rect 157108 409382 289772 409438
rect 289828 409382 289844 409438
rect 157036 409366 289844 409382
rect 291436 409438 532772 409454
rect 291436 409382 291452 409438
rect 291508 409382 532700 409438
rect 532756 409382 532772 409438
rect 291436 409366 532772 409382
rect 288860 409258 537700 409274
rect 288860 409202 288876 409258
rect 288932 409202 537628 409258
rect 537684 409202 537700 409258
rect 288860 409186 537700 409202
rect 7516 409078 295668 409094
rect 7516 409022 7532 409078
rect 7588 409022 295596 409078
rect 295652 409022 295668 409078
rect 7516 409006 295668 409022
rect 356060 409078 590564 409094
rect 356060 409022 356076 409078
rect 356132 409022 590492 409078
rect 590548 409022 590564 409078
rect 356060 409006 590564 409022
rect 150316 407998 300708 408014
rect 150316 407942 150332 407998
rect 150388 407942 299852 407998
rect 299908 407942 300636 407998
rect 300692 407942 300708 407998
rect 150316 407926 300708 407942
rect 187836 407818 339684 407834
rect 187836 407762 187852 407818
rect 187908 407762 339612 407818
rect 339668 407762 339684 407818
rect 187836 407746 339684 407762
rect 187724 407638 339796 407654
rect 187724 407582 187740 407638
rect 187796 407582 339724 407638
rect 339780 407582 339796 407638
rect 187724 407566 339796 407582
rect 288076 407458 532884 407474
rect 288076 407402 288092 407458
rect 288148 407402 532812 407458
rect 532868 407402 532884 407458
rect 288076 407386 532884 407402
rect 348556 407278 444964 407294
rect 348556 407222 348572 407278
rect 348628 407222 444892 407278
rect 444948 407222 444964 407278
rect 348556 407206 444964 407222
rect 355276 407098 496484 407114
rect 355276 407042 355292 407098
rect 355348 407042 496412 407098
rect 496468 407042 496484 407098
rect 355276 407026 496484 407042
rect 353820 406918 522244 406934
rect 353820 406862 353836 406918
rect 353892 406862 522172 406918
rect 522228 406862 522244 406918
rect 353820 406846 522244 406862
rect 353596 406738 527396 406754
rect 353596 406682 353612 406738
rect 353668 406682 527324 406738
rect 527380 406682 527396 406738
rect 353596 406666 527396 406682
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 66574 406350
rect 66630 406294 66698 406350
rect 66754 406294 71894 406350
rect 71950 406294 72018 406350
rect 72074 406294 77214 406350
rect 77270 406294 77338 406350
rect 77394 406294 82534 406350
rect 82590 406294 82658 406350
rect 82714 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 66574 406226
rect 66630 406170 66698 406226
rect 66754 406170 71894 406226
rect 71950 406170 72018 406226
rect 72074 406170 77214 406226
rect 77270 406170 77338 406226
rect 77394 406170 82534 406226
rect 82590 406170 82658 406226
rect 82714 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 66574 406102
rect 66630 406046 66698 406102
rect 66754 406046 71894 406102
rect 71950 406046 72018 406102
rect 72074 406046 77214 406102
rect 77270 406046 77338 406102
rect 77394 406046 82534 406102
rect 82590 406046 82658 406102
rect 82714 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 66574 405978
rect 66630 405922 66698 405978
rect 66754 405922 71894 405978
rect 71950 405922 72018 405978
rect 72074 405922 77214 405978
rect 77270 405922 77338 405978
rect 77394 405922 82534 405978
rect 82590 405922 82658 405978
rect 82714 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect 290540 405658 536020 405674
rect 290540 405602 290556 405658
rect 290612 405602 535948 405658
rect 536004 405602 536020 405658
rect 290540 405586 536020 405602
rect 301516 405478 532996 405494
rect 301516 405422 301532 405478
rect 301588 405422 532924 405478
rect 532980 405422 532996 405478
rect 301516 405406 532996 405422
rect 209900 404398 541844 404414
rect 209900 404342 209916 404398
rect 209972 404342 541772 404398
rect 541828 404342 541844 404398
rect 209900 404326 541844 404342
rect 208108 404218 540164 404234
rect 208108 404162 208124 404218
rect 208180 404162 540092 404218
rect 540148 404162 540164 404218
rect 208108 404146 540164 404162
rect 184588 404038 590900 404054
rect 184588 403982 184604 404038
rect 184660 403982 590828 404038
rect 590884 403982 590900 404038
rect 184588 403966 590900 403982
rect 184700 403318 591236 403334
rect 184700 403262 184716 403318
rect 184772 403262 591164 403318
rect 591220 403262 591236 403318
rect 184700 403246 591236 403262
rect 209788 402778 543524 402794
rect 209788 402722 209804 402778
rect 209860 402722 543452 402778
rect 543508 402722 543524 402778
rect 209788 402706 543524 402722
rect 186268 402598 591012 402614
rect 186268 402542 186284 402598
rect 186340 402542 590940 402598
rect 590996 402542 591012 402598
rect 186268 402526 591012 402542
rect 182908 402418 590676 402434
rect 182908 402362 182924 402418
rect 182980 402362 590604 402418
rect 590660 402362 590676 402418
rect 182908 402346 590676 402362
rect 201388 401698 592244 401714
rect 201388 401642 201404 401698
rect 201460 401642 592172 401698
rect 592228 401642 592244 401698
rect 201388 401626 592244 401642
rect 355724 400618 590564 400634
rect 355724 400562 355740 400618
rect 355796 400562 590492 400618
rect 590548 400562 590564 400618
rect 355724 400546 590564 400562
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 63914 400350
rect 63970 400294 64038 400350
rect 64094 400294 69234 400350
rect 69290 400294 69358 400350
rect 69414 400294 74554 400350
rect 74610 400294 74678 400350
rect 74734 400294 79874 400350
rect 79930 400294 79998 400350
rect 80054 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 63914 400226
rect 63970 400170 64038 400226
rect 64094 400170 69234 400226
rect 69290 400170 69358 400226
rect 69414 400170 74554 400226
rect 74610 400170 74678 400226
rect 74734 400170 79874 400226
rect 79930 400170 79998 400226
rect 80054 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 63914 400102
rect 63970 400046 64038 400102
rect 64094 400046 69234 400102
rect 69290 400046 69358 400102
rect 69414 400046 74554 400102
rect 74610 400046 74678 400102
rect 74734 400046 79874 400102
rect 79930 400046 79998 400102
rect 80054 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 63914 399978
rect 63970 399922 64038 399978
rect 64094 399922 69234 399978
rect 69290 399922 69358 399978
rect 69414 399922 74554 399978
rect 74610 399922 74678 399978
rect 74734 399922 79874 399978
rect 79930 399922 79998 399978
rect 80054 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect 267020 398998 534340 399014
rect 267020 398942 267036 398998
rect 267092 398942 534268 398998
rect 534324 398942 534340 398998
rect 267020 398926 534340 398942
rect 344076 398638 586420 398654
rect 344076 398582 344092 398638
rect 344148 398582 586348 398638
rect 586404 398582 586420 398638
rect 344076 398566 586420 398582
rect 239468 398458 591124 398474
rect 239468 398402 239484 398458
rect 239540 398402 591052 398458
rect 591108 398402 591124 398458
rect 239468 398386 591124 398402
rect 206428 398278 590900 398294
rect 206428 398222 206444 398278
rect 206500 398222 590828 398278
rect 590884 398222 590900 398278
rect 206428 398206 590900 398222
rect 187948 397378 340020 397394
rect 187948 397322 187964 397378
rect 188020 397322 339948 397378
rect 340004 397322 340020 397378
rect 187948 397306 340020 397322
rect 355164 397378 546324 397394
rect 355164 397322 355180 397378
rect 355236 397322 546252 397378
rect 546308 397322 546324 397378
rect 355164 397306 546324 397322
rect 355052 397198 574100 397214
rect 355052 397142 355068 397198
rect 355124 397142 574028 397198
rect 574084 397142 574100 397198
rect 355052 397126 574100 397142
rect 356060 397018 581044 397034
rect 356060 396962 356076 397018
rect 356132 396962 580972 397018
rect 581028 396962 581044 397018
rect 356060 396946 581044 396962
rect 312380 396838 553268 396854
rect 312380 396782 312396 396838
rect 312452 396782 553196 396838
rect 553252 396782 553268 396838
rect 312380 396766 553268 396782
rect 314060 396658 567156 396674
rect 314060 396602 314076 396658
rect 314132 396602 567084 396658
rect 567140 396602 567156 396658
rect 314060 396586 567156 396602
rect 281692 395578 490660 395594
rect 281692 395522 281708 395578
rect 281764 395522 490588 395578
rect 490644 395522 490660 395578
rect 281692 395506 490660 395522
rect 344188 395398 584852 395414
rect 344188 395342 344204 395398
rect 344260 395342 584780 395398
rect 584836 395342 584852 395398
rect 344188 395326 584852 395342
rect 343180 395218 586532 395234
rect 343180 395162 343196 395218
rect 343252 395162 586460 395218
rect 586516 395162 586532 395218
rect 343180 395146 586532 395162
rect 355276 395038 525604 395054
rect 355276 394982 355292 395038
rect 355348 394982 525532 395038
rect 525588 394982 525604 395038
rect 355276 394966 525604 394982
rect 226700 394858 584740 394874
rect 226700 394802 226716 394858
rect 226772 394802 584668 394858
rect 584724 394802 584740 394858
rect 226700 394786 584740 394802
rect 204748 393958 585524 393974
rect 204748 393902 204764 393958
rect 204820 393902 585452 393958
rect 585508 393902 585524 393958
rect 204748 393886 585524 393902
rect 203180 393778 587204 393794
rect 203180 393722 203196 393778
rect 203252 393722 587132 393778
rect 587188 393722 587204 393778
rect 203180 393706 587204 393722
rect 206540 393598 590676 393614
rect 206540 393542 206556 393598
rect 206612 393542 590604 393598
rect 590660 393542 590676 393598
rect 206540 393526 590676 393542
rect 203068 393418 587428 393434
rect 203068 393362 203084 393418
rect 203140 393362 587356 393418
rect 587412 393362 587428 393418
rect 203068 393346 587428 393362
rect 204860 393238 592356 393254
rect 204860 393182 204876 393238
rect 204932 393182 592284 393238
rect 592340 393182 592356 393238
rect 204860 393166 592356 393182
rect 239356 392698 364548 392714
rect 239356 392642 239372 392698
rect 239428 392642 364476 392698
rect 364532 392642 364548 392698
rect 239356 392626 364548 392642
rect 260300 392518 356484 392534
rect 260300 392462 260316 392518
rect 260372 392462 356412 392518
rect 356468 392462 356484 392518
rect 260300 392446 356484 392462
rect 250220 392338 356596 392354
rect 250220 392282 250236 392338
rect 250292 392282 356524 392338
rect 356580 392282 356596 392338
rect 250220 392266 356596 392282
rect 315740 391078 356148 391094
rect 315740 391022 315756 391078
rect 315812 391022 356076 391078
rect 356132 391022 356148 391078
rect 315740 391006 356148 391022
rect 293900 390898 356708 390914
rect 293900 390842 293916 390898
rect 293972 390842 356636 390898
rect 356692 390842 356708 390898
rect 293900 390826 356708 390842
rect 189516 390718 342820 390734
rect 189516 390662 189532 390718
rect 189588 390662 342748 390718
rect 342804 390662 342820 390718
rect 189516 390646 342820 390662
rect 62060 390538 322660 390554
rect 62060 390482 62076 390538
rect 62132 390482 322588 390538
rect 322644 390482 322660 390538
rect 62060 390466 322660 390482
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 374878 388350
rect 374934 388294 375002 388350
rect 375058 388294 405598 388350
rect 405654 388294 405722 388350
rect 405778 388294 436318 388350
rect 436374 388294 436442 388350
rect 436498 388294 467038 388350
rect 467094 388294 467162 388350
rect 467218 388294 497758 388350
rect 497814 388294 497882 388350
rect 497938 388294 528478 388350
rect 528534 388294 528602 388350
rect 528658 388294 559198 388350
rect 559254 388294 559322 388350
rect 559378 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 374878 388226
rect 374934 388170 375002 388226
rect 375058 388170 405598 388226
rect 405654 388170 405722 388226
rect 405778 388170 436318 388226
rect 436374 388170 436442 388226
rect 436498 388170 467038 388226
rect 467094 388170 467162 388226
rect 467218 388170 497758 388226
rect 497814 388170 497882 388226
rect 497938 388170 528478 388226
rect 528534 388170 528602 388226
rect 528658 388170 559198 388226
rect 559254 388170 559322 388226
rect 559378 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 374878 388102
rect 374934 388046 375002 388102
rect 375058 388046 405598 388102
rect 405654 388046 405722 388102
rect 405778 388046 436318 388102
rect 436374 388046 436442 388102
rect 436498 388046 467038 388102
rect 467094 388046 467162 388102
rect 467218 388046 497758 388102
rect 497814 388046 497882 388102
rect 497938 388046 528478 388102
rect 528534 388046 528602 388102
rect 528658 388046 559198 388102
rect 559254 388046 559322 388102
rect 559378 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 374878 387978
rect 374934 387922 375002 387978
rect 375058 387922 405598 387978
rect 405654 387922 405722 387978
rect 405778 387922 436318 387978
rect 436374 387922 436442 387978
rect 436498 387922 467038 387978
rect 467094 387922 467162 387978
rect 467218 387922 497758 387978
rect 497814 387922 497882 387978
rect 497938 387922 528478 387978
rect 528534 387922 528602 387978
rect 528658 387922 559198 387978
rect 559254 387922 559322 387978
rect 559378 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 359518 382350
rect 359574 382294 359642 382350
rect 359698 382294 390238 382350
rect 390294 382294 390362 382350
rect 390418 382294 420958 382350
rect 421014 382294 421082 382350
rect 421138 382294 451678 382350
rect 451734 382294 451802 382350
rect 451858 382294 482398 382350
rect 482454 382294 482522 382350
rect 482578 382294 513118 382350
rect 513174 382294 513242 382350
rect 513298 382294 543838 382350
rect 543894 382294 543962 382350
rect 544018 382294 574558 382350
rect 574614 382294 574682 382350
rect 574738 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 359518 382226
rect 359574 382170 359642 382226
rect 359698 382170 390238 382226
rect 390294 382170 390362 382226
rect 390418 382170 420958 382226
rect 421014 382170 421082 382226
rect 421138 382170 451678 382226
rect 451734 382170 451802 382226
rect 451858 382170 482398 382226
rect 482454 382170 482522 382226
rect 482578 382170 513118 382226
rect 513174 382170 513242 382226
rect 513298 382170 543838 382226
rect 543894 382170 543962 382226
rect 544018 382170 574558 382226
rect 574614 382170 574682 382226
rect 574738 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 359518 382102
rect 359574 382046 359642 382102
rect 359698 382046 390238 382102
rect 390294 382046 390362 382102
rect 390418 382046 420958 382102
rect 421014 382046 421082 382102
rect 421138 382046 451678 382102
rect 451734 382046 451802 382102
rect 451858 382046 482398 382102
rect 482454 382046 482522 382102
rect 482578 382046 513118 382102
rect 513174 382046 513242 382102
rect 513298 382046 543838 382102
rect 543894 382046 543962 382102
rect 544018 382046 574558 382102
rect 574614 382046 574682 382102
rect 574738 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 359518 381978
rect 359574 381922 359642 381978
rect 359698 381922 390238 381978
rect 390294 381922 390362 381978
rect 390418 381922 420958 381978
rect 421014 381922 421082 381978
rect 421138 381922 451678 381978
rect 451734 381922 451802 381978
rect 451858 381922 482398 381978
rect 482454 381922 482522 381978
rect 482578 381922 513118 381978
rect 513174 381922 513242 381978
rect 513298 381922 543838 381978
rect 543894 381922 543962 381978
rect 544018 381922 574558 381978
rect 574614 381922 574682 381978
rect 574738 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect 186380 381358 315828 381374
rect 186380 381302 186396 381358
rect 186452 381302 315756 381358
rect 315812 381302 315828 381358
rect 186380 381286 315828 381302
rect 299836 380818 341924 380834
rect 299836 380762 299852 380818
rect 299908 380762 341852 380818
rect 341908 380762 341924 380818
rect 299836 380746 341924 380762
rect 295580 380638 338676 380654
rect 295580 380582 295596 380638
rect 295652 380582 338604 380638
rect 338660 380582 338676 380638
rect 295580 380566 338676 380582
rect 280460 380458 338564 380474
rect 280460 380402 280476 380458
rect 280532 380402 338492 380458
rect 338548 380402 338564 380458
rect 280460 380386 338564 380402
rect 31036 378838 224100 378854
rect 31036 378782 31052 378838
rect 31108 378782 224028 378838
rect 224084 378782 224100 378838
rect 31036 378766 224100 378782
rect 29356 377398 225220 377414
rect 29356 377342 29372 377398
rect 29428 377342 225148 377398
rect 225204 377342 225220 377398
rect 29356 377326 225220 377342
rect 4156 377218 225892 377234
rect 4156 377162 4172 377218
rect 4228 377162 225820 377218
rect 225876 377162 225892 377218
rect 4156 377146 225892 377162
rect 4156 376318 238660 376334
rect 4156 376262 4172 376318
rect 4228 376262 238588 376318
rect 238644 376262 238660 376318
rect 4156 376246 238660 376262
rect 39660 373798 232612 373814
rect 39660 373742 39676 373798
rect 39732 373742 232540 373798
rect 232596 373742 232612 373798
rect 39660 373726 232612 373742
rect 12556 372178 222084 372194
rect 12556 372122 12572 372178
rect 12628 372122 222012 372178
rect 222068 372122 222084 372178
rect 12556 372106 222084 372122
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 209878 370350
rect 209934 370294 210002 370350
rect 210058 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 240598 370350
rect 240654 370294 240722 370350
rect 240778 370294 271318 370350
rect 271374 370294 271442 370350
rect 271498 370294 302038 370350
rect 302094 370294 302162 370350
rect 302218 370294 332758 370350
rect 332814 370294 332882 370350
rect 332938 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 374878 370350
rect 374934 370294 375002 370350
rect 375058 370294 405598 370350
rect 405654 370294 405722 370350
rect 405778 370294 436318 370350
rect 436374 370294 436442 370350
rect 436498 370294 467038 370350
rect 467094 370294 467162 370350
rect 467218 370294 497758 370350
rect 497814 370294 497882 370350
rect 497938 370294 528478 370350
rect 528534 370294 528602 370350
rect 528658 370294 559198 370350
rect 559254 370294 559322 370350
rect 559378 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 209878 370226
rect 209934 370170 210002 370226
rect 210058 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 240598 370226
rect 240654 370170 240722 370226
rect 240778 370170 271318 370226
rect 271374 370170 271442 370226
rect 271498 370170 302038 370226
rect 302094 370170 302162 370226
rect 302218 370170 332758 370226
rect 332814 370170 332882 370226
rect 332938 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 374878 370226
rect 374934 370170 375002 370226
rect 375058 370170 405598 370226
rect 405654 370170 405722 370226
rect 405778 370170 436318 370226
rect 436374 370170 436442 370226
rect 436498 370170 467038 370226
rect 467094 370170 467162 370226
rect 467218 370170 497758 370226
rect 497814 370170 497882 370226
rect 497938 370170 528478 370226
rect 528534 370170 528602 370226
rect 528658 370170 559198 370226
rect 559254 370170 559322 370226
rect 559378 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 209878 370102
rect 209934 370046 210002 370102
rect 210058 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 240598 370102
rect 240654 370046 240722 370102
rect 240778 370046 271318 370102
rect 271374 370046 271442 370102
rect 271498 370046 302038 370102
rect 302094 370046 302162 370102
rect 302218 370046 332758 370102
rect 332814 370046 332882 370102
rect 332938 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 374878 370102
rect 374934 370046 375002 370102
rect 375058 370046 405598 370102
rect 405654 370046 405722 370102
rect 405778 370046 436318 370102
rect 436374 370046 436442 370102
rect 436498 370046 467038 370102
rect 467094 370046 467162 370102
rect 467218 370046 497758 370102
rect 497814 370046 497882 370102
rect 497938 370046 528478 370102
rect 528534 370046 528602 370102
rect 528658 370046 559198 370102
rect 559254 370046 559322 370102
rect 559378 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 209878 369978
rect 209934 369922 210002 369978
rect 210058 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 240598 369978
rect 240654 369922 240722 369978
rect 240778 369922 271318 369978
rect 271374 369922 271442 369978
rect 271498 369922 302038 369978
rect 302094 369922 302162 369978
rect 302218 369922 332758 369978
rect 332814 369922 332882 369978
rect 332938 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 374878 369978
rect 374934 369922 375002 369978
rect 375058 369922 405598 369978
rect 405654 369922 405722 369978
rect 405778 369922 436318 369978
rect 436374 369922 436442 369978
rect 436498 369922 467038 369978
rect 467094 369922 467162 369978
rect 467218 369922 497758 369978
rect 497814 369922 497882 369978
rect 497938 369922 528478 369978
rect 528534 369922 528602 369978
rect 528658 369922 559198 369978
rect 559254 369922 559322 369978
rect 559378 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect 190636 368038 210884 368054
rect 190636 367982 190652 368038
rect 190708 367982 210812 368038
rect 210868 367982 210884 368038
rect 190636 367966 210884 367982
rect 190636 366598 214244 366614
rect 190636 366542 190652 366598
rect 190708 366542 214172 366598
rect 214228 366542 214244 366598
rect 190636 366526 214244 366542
rect 190636 366418 217604 366434
rect 190636 366362 190652 366418
rect 190708 366362 217532 366418
rect 217588 366362 217604 366418
rect 190636 366346 217604 366362
rect 190636 364618 214356 364634
rect 190636 364562 190652 364618
rect 190708 364562 214284 364618
rect 214340 364562 214356 364618
rect 190636 364546 214356 364562
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 194518 364350
rect 194574 364294 194642 364350
rect 194698 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 225238 364350
rect 225294 364294 225362 364350
rect 225418 364294 255958 364350
rect 256014 364294 256082 364350
rect 256138 364294 286678 364350
rect 286734 364294 286802 364350
rect 286858 364294 317398 364350
rect 317454 364294 317522 364350
rect 317578 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 359518 364350
rect 359574 364294 359642 364350
rect 359698 364294 390238 364350
rect 390294 364294 390362 364350
rect 390418 364294 420958 364350
rect 421014 364294 421082 364350
rect 421138 364294 451678 364350
rect 451734 364294 451802 364350
rect 451858 364294 482398 364350
rect 482454 364294 482522 364350
rect 482578 364294 513118 364350
rect 513174 364294 513242 364350
rect 513298 364294 543838 364350
rect 543894 364294 543962 364350
rect 544018 364294 574558 364350
rect 574614 364294 574682 364350
rect 574738 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 194518 364226
rect 194574 364170 194642 364226
rect 194698 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 225238 364226
rect 225294 364170 225362 364226
rect 225418 364170 255958 364226
rect 256014 364170 256082 364226
rect 256138 364170 286678 364226
rect 286734 364170 286802 364226
rect 286858 364170 317398 364226
rect 317454 364170 317522 364226
rect 317578 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 359518 364226
rect 359574 364170 359642 364226
rect 359698 364170 390238 364226
rect 390294 364170 390362 364226
rect 390418 364170 420958 364226
rect 421014 364170 421082 364226
rect 421138 364170 451678 364226
rect 451734 364170 451802 364226
rect 451858 364170 482398 364226
rect 482454 364170 482522 364226
rect 482578 364170 513118 364226
rect 513174 364170 513242 364226
rect 513298 364170 543838 364226
rect 543894 364170 543962 364226
rect 544018 364170 574558 364226
rect 574614 364170 574682 364226
rect 574738 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 194518 364102
rect 194574 364046 194642 364102
rect 194698 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 225238 364102
rect 225294 364046 225362 364102
rect 225418 364046 255958 364102
rect 256014 364046 256082 364102
rect 256138 364046 286678 364102
rect 286734 364046 286802 364102
rect 286858 364046 317398 364102
rect 317454 364046 317522 364102
rect 317578 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 359518 364102
rect 359574 364046 359642 364102
rect 359698 364046 390238 364102
rect 390294 364046 390362 364102
rect 390418 364046 420958 364102
rect 421014 364046 421082 364102
rect 421138 364046 451678 364102
rect 451734 364046 451802 364102
rect 451858 364046 482398 364102
rect 482454 364046 482522 364102
rect 482578 364046 513118 364102
rect 513174 364046 513242 364102
rect 513298 364046 543838 364102
rect 543894 364046 543962 364102
rect 544018 364046 574558 364102
rect 574614 364046 574682 364102
rect 574738 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 194518 363978
rect 194574 363922 194642 363978
rect 194698 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 225238 363978
rect 225294 363922 225362 363978
rect 225418 363922 255958 363978
rect 256014 363922 256082 363978
rect 256138 363922 286678 363978
rect 286734 363922 286802 363978
rect 286858 363922 317398 363978
rect 317454 363922 317522 363978
rect 317578 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 359518 363978
rect 359574 363922 359642 363978
rect 359698 363922 390238 363978
rect 390294 363922 390362 363978
rect 390418 363922 420958 363978
rect 421014 363922 421082 363978
rect 421138 363922 451678 363978
rect 451734 363922 451802 363978
rect 451858 363922 482398 363978
rect 482454 363922 482522 363978
rect 482578 363922 513118 363978
rect 513174 363922 513242 363978
rect 513298 363922 543838 363978
rect 543894 363922 543962 363978
rect 544018 363922 574558 363978
rect 574614 363922 574682 363978
rect 574738 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect 86476 356158 91716 356174
rect 86476 356102 86492 356158
rect 86548 356102 91644 356158
rect 91700 356102 91716 356158
rect 86476 356086 91716 356102
rect 89836 354358 93732 354374
rect 89836 354302 89852 354358
rect 89908 354302 93660 354358
rect 93716 354302 93732 354358
rect 89836 354286 93732 354302
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 69878 352350
rect 69934 352294 70002 352350
rect 70058 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 139878 352350
rect 139934 352294 140002 352350
rect 140058 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 209878 352350
rect 209934 352294 210002 352350
rect 210058 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 240598 352350
rect 240654 352294 240722 352350
rect 240778 352294 271318 352350
rect 271374 352294 271442 352350
rect 271498 352294 302038 352350
rect 302094 352294 302162 352350
rect 302218 352294 332758 352350
rect 332814 352294 332882 352350
rect 332938 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 374878 352350
rect 374934 352294 375002 352350
rect 375058 352294 405598 352350
rect 405654 352294 405722 352350
rect 405778 352294 436318 352350
rect 436374 352294 436442 352350
rect 436498 352294 467038 352350
rect 467094 352294 467162 352350
rect 467218 352294 497758 352350
rect 497814 352294 497882 352350
rect 497938 352294 528478 352350
rect 528534 352294 528602 352350
rect 528658 352294 559198 352350
rect 559254 352294 559322 352350
rect 559378 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 69878 352226
rect 69934 352170 70002 352226
rect 70058 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 139878 352226
rect 139934 352170 140002 352226
rect 140058 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 209878 352226
rect 209934 352170 210002 352226
rect 210058 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 240598 352226
rect 240654 352170 240722 352226
rect 240778 352170 271318 352226
rect 271374 352170 271442 352226
rect 271498 352170 302038 352226
rect 302094 352170 302162 352226
rect 302218 352170 332758 352226
rect 332814 352170 332882 352226
rect 332938 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 374878 352226
rect 374934 352170 375002 352226
rect 375058 352170 405598 352226
rect 405654 352170 405722 352226
rect 405778 352170 436318 352226
rect 436374 352170 436442 352226
rect 436498 352170 467038 352226
rect 467094 352170 467162 352226
rect 467218 352170 497758 352226
rect 497814 352170 497882 352226
rect 497938 352170 528478 352226
rect 528534 352170 528602 352226
rect 528658 352170 559198 352226
rect 559254 352170 559322 352226
rect 559378 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 69878 352102
rect 69934 352046 70002 352102
rect 70058 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 139878 352102
rect 139934 352046 140002 352102
rect 140058 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 209878 352102
rect 209934 352046 210002 352102
rect 210058 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 240598 352102
rect 240654 352046 240722 352102
rect 240778 352046 271318 352102
rect 271374 352046 271442 352102
rect 271498 352046 302038 352102
rect 302094 352046 302162 352102
rect 302218 352046 332758 352102
rect 332814 352046 332882 352102
rect 332938 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 374878 352102
rect 374934 352046 375002 352102
rect 375058 352046 405598 352102
rect 405654 352046 405722 352102
rect 405778 352046 436318 352102
rect 436374 352046 436442 352102
rect 436498 352046 467038 352102
rect 467094 352046 467162 352102
rect 467218 352046 497758 352102
rect 497814 352046 497882 352102
rect 497938 352046 528478 352102
rect 528534 352046 528602 352102
rect 528658 352046 559198 352102
rect 559254 352046 559322 352102
rect 559378 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 69878 351978
rect 69934 351922 70002 351978
rect 70058 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 139878 351978
rect 139934 351922 140002 351978
rect 140058 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 209878 351978
rect 209934 351922 210002 351978
rect 210058 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 240598 351978
rect 240654 351922 240722 351978
rect 240778 351922 271318 351978
rect 271374 351922 271442 351978
rect 271498 351922 302038 351978
rect 302094 351922 302162 351978
rect 302218 351922 332758 351978
rect 332814 351922 332882 351978
rect 332938 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 374878 351978
rect 374934 351922 375002 351978
rect 375058 351922 405598 351978
rect 405654 351922 405722 351978
rect 405778 351922 436318 351978
rect 436374 351922 436442 351978
rect 436498 351922 467038 351978
rect 467094 351922 467162 351978
rect 467218 351922 497758 351978
rect 497814 351922 497882 351978
rect 497938 351922 528478 351978
rect 528534 351922 528602 351978
rect 528658 351922 559198 351978
rect 559254 351922 559322 351978
rect 559378 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 54518 346350
rect 54574 346294 54642 346350
rect 54698 346294 85238 346350
rect 85294 346294 85362 346350
rect 85418 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 124518 346350
rect 124574 346294 124642 346350
rect 124698 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 155238 346350
rect 155294 346294 155362 346350
rect 155418 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 194518 346350
rect 194574 346294 194642 346350
rect 194698 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 225238 346350
rect 225294 346294 225362 346350
rect 225418 346294 255958 346350
rect 256014 346294 256082 346350
rect 256138 346294 286678 346350
rect 286734 346294 286802 346350
rect 286858 346294 317398 346350
rect 317454 346294 317522 346350
rect 317578 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 359518 346350
rect 359574 346294 359642 346350
rect 359698 346294 390238 346350
rect 390294 346294 390362 346350
rect 390418 346294 420958 346350
rect 421014 346294 421082 346350
rect 421138 346294 451678 346350
rect 451734 346294 451802 346350
rect 451858 346294 482398 346350
rect 482454 346294 482522 346350
rect 482578 346294 513118 346350
rect 513174 346294 513242 346350
rect 513298 346294 543838 346350
rect 543894 346294 543962 346350
rect 544018 346294 574558 346350
rect 574614 346294 574682 346350
rect 574738 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 54518 346226
rect 54574 346170 54642 346226
rect 54698 346170 85238 346226
rect 85294 346170 85362 346226
rect 85418 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 124518 346226
rect 124574 346170 124642 346226
rect 124698 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 155238 346226
rect 155294 346170 155362 346226
rect 155418 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 194518 346226
rect 194574 346170 194642 346226
rect 194698 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 225238 346226
rect 225294 346170 225362 346226
rect 225418 346170 255958 346226
rect 256014 346170 256082 346226
rect 256138 346170 286678 346226
rect 286734 346170 286802 346226
rect 286858 346170 317398 346226
rect 317454 346170 317522 346226
rect 317578 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 359518 346226
rect 359574 346170 359642 346226
rect 359698 346170 390238 346226
rect 390294 346170 390362 346226
rect 390418 346170 420958 346226
rect 421014 346170 421082 346226
rect 421138 346170 451678 346226
rect 451734 346170 451802 346226
rect 451858 346170 482398 346226
rect 482454 346170 482522 346226
rect 482578 346170 513118 346226
rect 513174 346170 513242 346226
rect 513298 346170 543838 346226
rect 543894 346170 543962 346226
rect 544018 346170 574558 346226
rect 574614 346170 574682 346226
rect 574738 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 54518 346102
rect 54574 346046 54642 346102
rect 54698 346046 85238 346102
rect 85294 346046 85362 346102
rect 85418 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 124518 346102
rect 124574 346046 124642 346102
rect 124698 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 155238 346102
rect 155294 346046 155362 346102
rect 155418 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 194518 346102
rect 194574 346046 194642 346102
rect 194698 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 225238 346102
rect 225294 346046 225362 346102
rect 225418 346046 255958 346102
rect 256014 346046 256082 346102
rect 256138 346046 286678 346102
rect 286734 346046 286802 346102
rect 286858 346046 317398 346102
rect 317454 346046 317522 346102
rect 317578 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 359518 346102
rect 359574 346046 359642 346102
rect 359698 346046 390238 346102
rect 390294 346046 390362 346102
rect 390418 346046 420958 346102
rect 421014 346046 421082 346102
rect 421138 346046 451678 346102
rect 451734 346046 451802 346102
rect 451858 346046 482398 346102
rect 482454 346046 482522 346102
rect 482578 346046 513118 346102
rect 513174 346046 513242 346102
rect 513298 346046 543838 346102
rect 543894 346046 543962 346102
rect 544018 346046 574558 346102
rect 574614 346046 574682 346102
rect 574738 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 54518 345978
rect 54574 345922 54642 345978
rect 54698 345922 85238 345978
rect 85294 345922 85362 345978
rect 85418 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 124518 345978
rect 124574 345922 124642 345978
rect 124698 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 155238 345978
rect 155294 345922 155362 345978
rect 155418 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 194518 345978
rect 194574 345922 194642 345978
rect 194698 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 225238 345978
rect 225294 345922 225362 345978
rect 225418 345922 255958 345978
rect 256014 345922 256082 345978
rect 256138 345922 286678 345978
rect 286734 345922 286802 345978
rect 286858 345922 317398 345978
rect 317454 345922 317522 345978
rect 317578 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 359518 345978
rect 359574 345922 359642 345978
rect 359698 345922 390238 345978
rect 390294 345922 390362 345978
rect 390418 345922 420958 345978
rect 421014 345922 421082 345978
rect 421138 345922 451678 345978
rect 451734 345922 451802 345978
rect 451858 345922 482398 345978
rect 482454 345922 482522 345978
rect 482578 345922 513118 345978
rect 513174 345922 513242 345978
rect 513298 345922 543838 345978
rect 543894 345922 543962 345978
rect 544018 345922 574558 345978
rect 574614 345922 574682 345978
rect 574738 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect 338140 342478 339348 342494
rect 338140 342422 338156 342478
rect 338212 342422 339276 342478
rect 339332 342422 339348 342478
rect 338140 342406 339348 342422
rect 168012 340138 206740 340154
rect 168012 340082 168028 340138
rect 168084 340082 206668 340138
rect 206724 340082 206740 340138
rect 168012 340066 206740 340082
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 69878 334350
rect 69934 334294 70002 334350
rect 70058 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 139878 334350
rect 139934 334294 140002 334350
rect 140058 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 209878 334350
rect 209934 334294 210002 334350
rect 210058 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 240598 334350
rect 240654 334294 240722 334350
rect 240778 334294 271318 334350
rect 271374 334294 271442 334350
rect 271498 334294 302038 334350
rect 302094 334294 302162 334350
rect 302218 334294 332758 334350
rect 332814 334294 332882 334350
rect 332938 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 374878 334350
rect 374934 334294 375002 334350
rect 375058 334294 405598 334350
rect 405654 334294 405722 334350
rect 405778 334294 436318 334350
rect 436374 334294 436442 334350
rect 436498 334294 467038 334350
rect 467094 334294 467162 334350
rect 467218 334294 497758 334350
rect 497814 334294 497882 334350
rect 497938 334294 528478 334350
rect 528534 334294 528602 334350
rect 528658 334294 559198 334350
rect 559254 334294 559322 334350
rect 559378 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 69878 334226
rect 69934 334170 70002 334226
rect 70058 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 139878 334226
rect 139934 334170 140002 334226
rect 140058 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 209878 334226
rect 209934 334170 210002 334226
rect 210058 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 240598 334226
rect 240654 334170 240722 334226
rect 240778 334170 271318 334226
rect 271374 334170 271442 334226
rect 271498 334170 302038 334226
rect 302094 334170 302162 334226
rect 302218 334170 332758 334226
rect 332814 334170 332882 334226
rect 332938 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 374878 334226
rect 374934 334170 375002 334226
rect 375058 334170 405598 334226
rect 405654 334170 405722 334226
rect 405778 334170 436318 334226
rect 436374 334170 436442 334226
rect 436498 334170 467038 334226
rect 467094 334170 467162 334226
rect 467218 334170 497758 334226
rect 497814 334170 497882 334226
rect 497938 334170 528478 334226
rect 528534 334170 528602 334226
rect 528658 334170 559198 334226
rect 559254 334170 559322 334226
rect 559378 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 69878 334102
rect 69934 334046 70002 334102
rect 70058 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 139878 334102
rect 139934 334046 140002 334102
rect 140058 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 209878 334102
rect 209934 334046 210002 334102
rect 210058 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 240598 334102
rect 240654 334046 240722 334102
rect 240778 334046 271318 334102
rect 271374 334046 271442 334102
rect 271498 334046 302038 334102
rect 302094 334046 302162 334102
rect 302218 334046 332758 334102
rect 332814 334046 332882 334102
rect 332938 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 374878 334102
rect 374934 334046 375002 334102
rect 375058 334046 405598 334102
rect 405654 334046 405722 334102
rect 405778 334046 436318 334102
rect 436374 334046 436442 334102
rect 436498 334046 467038 334102
rect 467094 334046 467162 334102
rect 467218 334046 497758 334102
rect 497814 334046 497882 334102
rect 497938 334046 528478 334102
rect 528534 334046 528602 334102
rect 528658 334046 559198 334102
rect 559254 334046 559322 334102
rect 559378 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 69878 333978
rect 69934 333922 70002 333978
rect 70058 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 139878 333978
rect 139934 333922 140002 333978
rect 140058 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 209878 333978
rect 209934 333922 210002 333978
rect 210058 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 240598 333978
rect 240654 333922 240722 333978
rect 240778 333922 271318 333978
rect 271374 333922 271442 333978
rect 271498 333922 302038 333978
rect 302094 333922 302162 333978
rect 302218 333922 332758 333978
rect 332814 333922 332882 333978
rect 332938 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 374878 333978
rect 374934 333922 375002 333978
rect 375058 333922 405598 333978
rect 405654 333922 405722 333978
rect 405778 333922 436318 333978
rect 436374 333922 436442 333978
rect 436498 333922 467038 333978
rect 467094 333922 467162 333978
rect 467218 333922 497758 333978
rect 497814 333922 497882 333978
rect 497938 333922 528478 333978
rect 528534 333922 528602 333978
rect 528658 333922 559198 333978
rect 559254 333922 559322 333978
rect 559378 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect 91628 332758 93508 332774
rect 91628 332702 91644 332758
rect 91700 332702 93436 332758
rect 93492 332702 93508 332758
rect 91628 332686 93508 332702
rect 91516 330958 93284 330974
rect 91516 330902 91532 330958
rect 91588 330902 93212 330958
rect 93268 330902 93284 330958
rect 91516 330886 93284 330902
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 54518 328350
rect 54574 328294 54642 328350
rect 54698 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 85238 328350
rect 85294 328294 85362 328350
rect 85418 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 124518 328350
rect 124574 328294 124642 328350
rect 124698 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 155238 328350
rect 155294 328294 155362 328350
rect 155418 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 194518 328350
rect 194574 328294 194642 328350
rect 194698 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 225238 328350
rect 225294 328294 225362 328350
rect 225418 328294 255958 328350
rect 256014 328294 256082 328350
rect 256138 328294 286678 328350
rect 286734 328294 286802 328350
rect 286858 328294 317398 328350
rect 317454 328294 317522 328350
rect 317578 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 359518 328350
rect 359574 328294 359642 328350
rect 359698 328294 390238 328350
rect 390294 328294 390362 328350
rect 390418 328294 420958 328350
rect 421014 328294 421082 328350
rect 421138 328294 451678 328350
rect 451734 328294 451802 328350
rect 451858 328294 482398 328350
rect 482454 328294 482522 328350
rect 482578 328294 513118 328350
rect 513174 328294 513242 328350
rect 513298 328294 543838 328350
rect 543894 328294 543962 328350
rect 544018 328294 574558 328350
rect 574614 328294 574682 328350
rect 574738 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 54518 328226
rect 54574 328170 54642 328226
rect 54698 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 85238 328226
rect 85294 328170 85362 328226
rect 85418 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 124518 328226
rect 124574 328170 124642 328226
rect 124698 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 155238 328226
rect 155294 328170 155362 328226
rect 155418 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 194518 328226
rect 194574 328170 194642 328226
rect 194698 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 225238 328226
rect 225294 328170 225362 328226
rect 225418 328170 255958 328226
rect 256014 328170 256082 328226
rect 256138 328170 286678 328226
rect 286734 328170 286802 328226
rect 286858 328170 317398 328226
rect 317454 328170 317522 328226
rect 317578 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 359518 328226
rect 359574 328170 359642 328226
rect 359698 328170 390238 328226
rect 390294 328170 390362 328226
rect 390418 328170 420958 328226
rect 421014 328170 421082 328226
rect 421138 328170 451678 328226
rect 451734 328170 451802 328226
rect 451858 328170 482398 328226
rect 482454 328170 482522 328226
rect 482578 328170 513118 328226
rect 513174 328170 513242 328226
rect 513298 328170 543838 328226
rect 543894 328170 543962 328226
rect 544018 328170 574558 328226
rect 574614 328170 574682 328226
rect 574738 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 54518 328102
rect 54574 328046 54642 328102
rect 54698 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 85238 328102
rect 85294 328046 85362 328102
rect 85418 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 124518 328102
rect 124574 328046 124642 328102
rect 124698 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 155238 328102
rect 155294 328046 155362 328102
rect 155418 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 194518 328102
rect 194574 328046 194642 328102
rect 194698 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 225238 328102
rect 225294 328046 225362 328102
rect 225418 328046 255958 328102
rect 256014 328046 256082 328102
rect 256138 328046 286678 328102
rect 286734 328046 286802 328102
rect 286858 328046 317398 328102
rect 317454 328046 317522 328102
rect 317578 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 359518 328102
rect 359574 328046 359642 328102
rect 359698 328046 390238 328102
rect 390294 328046 390362 328102
rect 390418 328046 420958 328102
rect 421014 328046 421082 328102
rect 421138 328046 451678 328102
rect 451734 328046 451802 328102
rect 451858 328046 482398 328102
rect 482454 328046 482522 328102
rect 482578 328046 513118 328102
rect 513174 328046 513242 328102
rect 513298 328046 543838 328102
rect 543894 328046 543962 328102
rect 544018 328046 574558 328102
rect 574614 328046 574682 328102
rect 574738 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 54518 327978
rect 54574 327922 54642 327978
rect 54698 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 85238 327978
rect 85294 327922 85362 327978
rect 85418 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 124518 327978
rect 124574 327922 124642 327978
rect 124698 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 155238 327978
rect 155294 327922 155362 327978
rect 155418 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 194518 327978
rect 194574 327922 194642 327978
rect 194698 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 225238 327978
rect 225294 327922 225362 327978
rect 225418 327922 255958 327978
rect 256014 327922 256082 327978
rect 256138 327922 286678 327978
rect 286734 327922 286802 327978
rect 286858 327922 317398 327978
rect 317454 327922 317522 327978
rect 317578 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 359518 327978
rect 359574 327922 359642 327978
rect 359698 327922 390238 327978
rect 390294 327922 390362 327978
rect 390418 327922 420958 327978
rect 421014 327922 421082 327978
rect 421138 327922 451678 327978
rect 451734 327922 451802 327978
rect 451858 327922 482398 327978
rect 482454 327922 482522 327978
rect 482578 327922 513118 327978
rect 513174 327922 513242 327978
rect 513298 327922 543838 327978
rect 543894 327922 543962 327978
rect 544018 327922 574558 327978
rect 574614 327922 574682 327978
rect 574738 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect 93308 322498 168100 322514
rect 93308 322442 93324 322498
rect 93380 322442 168028 322498
rect 168084 322442 168100 322498
rect 93308 322426 168100 322442
rect 93196 320878 168436 320894
rect 93196 320822 93212 320878
rect 93268 320822 168364 320878
rect 168420 320822 168436 320878
rect 93196 320806 168436 320822
rect 93420 320698 168324 320714
rect 93420 320642 93436 320698
rect 93492 320642 168252 320698
rect 168308 320642 168324 320698
rect 93420 320626 168324 320642
rect 93644 320518 168212 320534
rect 93644 320462 93660 320518
rect 93716 320462 168140 320518
rect 168196 320462 168212 320518
rect 93644 320446 168212 320462
rect 190636 319258 217716 319274
rect 190636 319202 190652 319258
rect 190708 319202 217644 319258
rect 217700 319202 217716 319258
rect 190636 319186 217716 319202
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 209878 316350
rect 209934 316294 210002 316350
rect 210058 316294 224274 316350
rect 224330 316294 224398 316350
rect 224454 316294 224522 316350
rect 224578 316294 224646 316350
rect 224702 316294 240598 316350
rect 240654 316294 240722 316350
rect 240778 316294 271318 316350
rect 271374 316294 271442 316350
rect 271498 316294 302038 316350
rect 302094 316294 302162 316350
rect 302218 316294 332758 316350
rect 332814 316294 332882 316350
rect 332938 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 374878 316350
rect 374934 316294 375002 316350
rect 375058 316294 405598 316350
rect 405654 316294 405722 316350
rect 405778 316294 436318 316350
rect 436374 316294 436442 316350
rect 436498 316294 467038 316350
rect 467094 316294 467162 316350
rect 467218 316294 497758 316350
rect 497814 316294 497882 316350
rect 497938 316294 528478 316350
rect 528534 316294 528602 316350
rect 528658 316294 559198 316350
rect 559254 316294 559322 316350
rect 559378 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 209878 316226
rect 209934 316170 210002 316226
rect 210058 316170 224274 316226
rect 224330 316170 224398 316226
rect 224454 316170 224522 316226
rect 224578 316170 224646 316226
rect 224702 316170 240598 316226
rect 240654 316170 240722 316226
rect 240778 316170 271318 316226
rect 271374 316170 271442 316226
rect 271498 316170 302038 316226
rect 302094 316170 302162 316226
rect 302218 316170 332758 316226
rect 332814 316170 332882 316226
rect 332938 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 374878 316226
rect 374934 316170 375002 316226
rect 375058 316170 405598 316226
rect 405654 316170 405722 316226
rect 405778 316170 436318 316226
rect 436374 316170 436442 316226
rect 436498 316170 467038 316226
rect 467094 316170 467162 316226
rect 467218 316170 497758 316226
rect 497814 316170 497882 316226
rect 497938 316170 528478 316226
rect 528534 316170 528602 316226
rect 528658 316170 559198 316226
rect 559254 316170 559322 316226
rect 559378 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 209878 316102
rect 209934 316046 210002 316102
rect 210058 316046 224274 316102
rect 224330 316046 224398 316102
rect 224454 316046 224522 316102
rect 224578 316046 224646 316102
rect 224702 316046 240598 316102
rect 240654 316046 240722 316102
rect 240778 316046 271318 316102
rect 271374 316046 271442 316102
rect 271498 316046 302038 316102
rect 302094 316046 302162 316102
rect 302218 316046 332758 316102
rect 332814 316046 332882 316102
rect 332938 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 374878 316102
rect 374934 316046 375002 316102
rect 375058 316046 405598 316102
rect 405654 316046 405722 316102
rect 405778 316046 436318 316102
rect 436374 316046 436442 316102
rect 436498 316046 467038 316102
rect 467094 316046 467162 316102
rect 467218 316046 497758 316102
rect 497814 316046 497882 316102
rect 497938 316046 528478 316102
rect 528534 316046 528602 316102
rect 528658 316046 559198 316102
rect 559254 316046 559322 316102
rect 559378 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 209878 315978
rect 209934 315922 210002 315978
rect 210058 315922 224274 315978
rect 224330 315922 224398 315978
rect 224454 315922 224522 315978
rect 224578 315922 224646 315978
rect 224702 315922 240598 315978
rect 240654 315922 240722 315978
rect 240778 315922 271318 315978
rect 271374 315922 271442 315978
rect 271498 315922 302038 315978
rect 302094 315922 302162 315978
rect 302218 315922 332758 315978
rect 332814 315922 332882 315978
rect 332938 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 374878 315978
rect 374934 315922 375002 315978
rect 375058 315922 405598 315978
rect 405654 315922 405722 315978
rect 405778 315922 436318 315978
rect 436374 315922 436442 315978
rect 436498 315922 467038 315978
rect 467094 315922 467162 315978
rect 467218 315922 497758 315978
rect 497814 315922 497882 315978
rect 497938 315922 528478 315978
rect 528534 315922 528602 315978
rect 528658 315922 559198 315978
rect 559254 315922 559322 315978
rect 559378 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect 60380 311698 237876 311714
rect 60380 311642 60396 311698
rect 60452 311642 237804 311698
rect 237860 311642 237876 311698
rect 60380 311626 237876 311642
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 194518 310350
rect 194574 310294 194642 310350
rect 194698 310294 220554 310350
rect 220610 310294 220678 310350
rect 220734 310294 220802 310350
rect 220858 310294 220926 310350
rect 220982 310294 225238 310350
rect 225294 310294 225362 310350
rect 225418 310294 255958 310350
rect 256014 310294 256082 310350
rect 256138 310294 286678 310350
rect 286734 310294 286802 310350
rect 286858 310294 317398 310350
rect 317454 310294 317522 310350
rect 317578 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 359518 310350
rect 359574 310294 359642 310350
rect 359698 310294 390238 310350
rect 390294 310294 390362 310350
rect 390418 310294 420958 310350
rect 421014 310294 421082 310350
rect 421138 310294 451678 310350
rect 451734 310294 451802 310350
rect 451858 310294 482398 310350
rect 482454 310294 482522 310350
rect 482578 310294 513118 310350
rect 513174 310294 513242 310350
rect 513298 310294 543838 310350
rect 543894 310294 543962 310350
rect 544018 310294 574558 310350
rect 574614 310294 574682 310350
rect 574738 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 194518 310226
rect 194574 310170 194642 310226
rect 194698 310170 220554 310226
rect 220610 310170 220678 310226
rect 220734 310170 220802 310226
rect 220858 310170 220926 310226
rect 220982 310170 225238 310226
rect 225294 310170 225362 310226
rect 225418 310170 255958 310226
rect 256014 310170 256082 310226
rect 256138 310170 286678 310226
rect 286734 310170 286802 310226
rect 286858 310170 317398 310226
rect 317454 310170 317522 310226
rect 317578 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 359518 310226
rect 359574 310170 359642 310226
rect 359698 310170 390238 310226
rect 390294 310170 390362 310226
rect 390418 310170 420958 310226
rect 421014 310170 421082 310226
rect 421138 310170 451678 310226
rect 451734 310170 451802 310226
rect 451858 310170 482398 310226
rect 482454 310170 482522 310226
rect 482578 310170 513118 310226
rect 513174 310170 513242 310226
rect 513298 310170 543838 310226
rect 543894 310170 543962 310226
rect 544018 310170 574558 310226
rect 574614 310170 574682 310226
rect 574738 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 194518 310102
rect 194574 310046 194642 310102
rect 194698 310046 220554 310102
rect 220610 310046 220678 310102
rect 220734 310046 220802 310102
rect 220858 310046 220926 310102
rect 220982 310046 225238 310102
rect 225294 310046 225362 310102
rect 225418 310046 255958 310102
rect 256014 310046 256082 310102
rect 256138 310046 286678 310102
rect 286734 310046 286802 310102
rect 286858 310046 317398 310102
rect 317454 310046 317522 310102
rect 317578 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 359518 310102
rect 359574 310046 359642 310102
rect 359698 310046 390238 310102
rect 390294 310046 390362 310102
rect 390418 310046 420958 310102
rect 421014 310046 421082 310102
rect 421138 310046 451678 310102
rect 451734 310046 451802 310102
rect 451858 310046 482398 310102
rect 482454 310046 482522 310102
rect 482578 310046 513118 310102
rect 513174 310046 513242 310102
rect 513298 310046 543838 310102
rect 543894 310046 543962 310102
rect 544018 310046 574558 310102
rect 574614 310046 574682 310102
rect 574738 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 194518 309978
rect 194574 309922 194642 309978
rect 194698 309922 220554 309978
rect 220610 309922 220678 309978
rect 220734 309922 220802 309978
rect 220858 309922 220926 309978
rect 220982 309922 225238 309978
rect 225294 309922 225362 309978
rect 225418 309922 255958 309978
rect 256014 309922 256082 309978
rect 256138 309922 286678 309978
rect 286734 309922 286802 309978
rect 286858 309922 317398 309978
rect 317454 309922 317522 309978
rect 317578 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 359518 309978
rect 359574 309922 359642 309978
rect 359698 309922 390238 309978
rect 390294 309922 390362 309978
rect 390418 309922 420958 309978
rect 421014 309922 421082 309978
rect 421138 309922 451678 309978
rect 451734 309922 451802 309978
rect 451858 309922 482398 309978
rect 482454 309922 482522 309978
rect 482578 309922 513118 309978
rect 513174 309922 513242 309978
rect 513298 309922 543838 309978
rect 543894 309922 543962 309978
rect 544018 309922 574558 309978
rect 574614 309922 574682 309978
rect 574738 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect 338252 301978 339460 301994
rect 338252 301922 338268 301978
rect 338324 301922 339388 301978
rect 339444 301922 339460 301978
rect 338252 301906 339460 301922
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 209878 298350
rect 209934 298294 210002 298350
rect 210058 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 240598 298350
rect 240654 298294 240722 298350
rect 240778 298294 271318 298350
rect 271374 298294 271442 298350
rect 271498 298294 302038 298350
rect 302094 298294 302162 298350
rect 302218 298294 332758 298350
rect 332814 298294 332882 298350
rect 332938 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 374878 298350
rect 374934 298294 375002 298350
rect 375058 298294 405598 298350
rect 405654 298294 405722 298350
rect 405778 298294 436318 298350
rect 436374 298294 436442 298350
rect 436498 298294 467038 298350
rect 467094 298294 467162 298350
rect 467218 298294 497758 298350
rect 497814 298294 497882 298350
rect 497938 298294 528478 298350
rect 528534 298294 528602 298350
rect 528658 298294 559198 298350
rect 559254 298294 559322 298350
rect 559378 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 209878 298226
rect 209934 298170 210002 298226
rect 210058 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 240598 298226
rect 240654 298170 240722 298226
rect 240778 298170 271318 298226
rect 271374 298170 271442 298226
rect 271498 298170 302038 298226
rect 302094 298170 302162 298226
rect 302218 298170 332758 298226
rect 332814 298170 332882 298226
rect 332938 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 374878 298226
rect 374934 298170 375002 298226
rect 375058 298170 405598 298226
rect 405654 298170 405722 298226
rect 405778 298170 436318 298226
rect 436374 298170 436442 298226
rect 436498 298170 467038 298226
rect 467094 298170 467162 298226
rect 467218 298170 497758 298226
rect 497814 298170 497882 298226
rect 497938 298170 528478 298226
rect 528534 298170 528602 298226
rect 528658 298170 559198 298226
rect 559254 298170 559322 298226
rect 559378 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 209878 298102
rect 209934 298046 210002 298102
rect 210058 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 240598 298102
rect 240654 298046 240722 298102
rect 240778 298046 271318 298102
rect 271374 298046 271442 298102
rect 271498 298046 302038 298102
rect 302094 298046 302162 298102
rect 302218 298046 332758 298102
rect 332814 298046 332882 298102
rect 332938 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 374878 298102
rect 374934 298046 375002 298102
rect 375058 298046 405598 298102
rect 405654 298046 405722 298102
rect 405778 298046 436318 298102
rect 436374 298046 436442 298102
rect 436498 298046 467038 298102
rect 467094 298046 467162 298102
rect 467218 298046 497758 298102
rect 497814 298046 497882 298102
rect 497938 298046 528478 298102
rect 528534 298046 528602 298102
rect 528658 298046 559198 298102
rect 559254 298046 559322 298102
rect 559378 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 209878 297978
rect 209934 297922 210002 297978
rect 210058 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 240598 297978
rect 240654 297922 240722 297978
rect 240778 297922 271318 297978
rect 271374 297922 271442 297978
rect 271498 297922 302038 297978
rect 302094 297922 302162 297978
rect 302218 297922 332758 297978
rect 332814 297922 332882 297978
rect 332938 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 374878 297978
rect 374934 297922 375002 297978
rect 375058 297922 405598 297978
rect 405654 297922 405722 297978
rect 405778 297922 436318 297978
rect 436374 297922 436442 297978
rect 436498 297922 467038 297978
rect 467094 297922 467162 297978
rect 467218 297922 497758 297978
rect 497814 297922 497882 297978
rect 497938 297922 528478 297978
rect 528534 297922 528602 297978
rect 528658 297922 559198 297978
rect 559254 297922 559322 297978
rect 559378 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect 4268 294778 239780 294794
rect 4268 294722 4284 294778
rect 4340 294722 238364 294778
rect 238420 294722 239708 294778
rect 239764 294722 239780 294778
rect 4268 294706 239780 294722
rect 71804 294058 236868 294074
rect 71804 294002 71820 294058
rect 71876 294002 236796 294058
rect 236852 294002 236868 294058
rect 71804 293986 236868 294002
rect 84572 293878 239892 293894
rect 84572 293822 84588 293878
rect 84644 293822 235116 293878
rect 235172 293822 239820 293878
rect 239876 293822 239892 293878
rect 84572 293806 239892 293822
rect 190636 292618 239668 292634
rect 190636 292562 190652 292618
rect 190708 292562 239596 292618
rect 239652 292562 239668 292618
rect 190636 292546 239668 292562
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 194518 292350
rect 194574 292294 194642 292350
rect 194698 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 225238 292350
rect 225294 292294 225362 292350
rect 225418 292294 255958 292350
rect 256014 292294 256082 292350
rect 256138 292294 286678 292350
rect 286734 292294 286802 292350
rect 286858 292294 317398 292350
rect 317454 292294 317522 292350
rect 317578 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 359518 292350
rect 359574 292294 359642 292350
rect 359698 292294 390238 292350
rect 390294 292294 390362 292350
rect 390418 292294 420958 292350
rect 421014 292294 421082 292350
rect 421138 292294 451678 292350
rect 451734 292294 451802 292350
rect 451858 292294 482398 292350
rect 482454 292294 482522 292350
rect 482578 292294 513118 292350
rect 513174 292294 513242 292350
rect 513298 292294 543838 292350
rect 543894 292294 543962 292350
rect 544018 292294 574558 292350
rect 574614 292294 574682 292350
rect 574738 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 194518 292226
rect 194574 292170 194642 292226
rect 194698 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 225238 292226
rect 225294 292170 225362 292226
rect 225418 292170 255958 292226
rect 256014 292170 256082 292226
rect 256138 292170 286678 292226
rect 286734 292170 286802 292226
rect 286858 292170 317398 292226
rect 317454 292170 317522 292226
rect 317578 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 359518 292226
rect 359574 292170 359642 292226
rect 359698 292170 390238 292226
rect 390294 292170 390362 292226
rect 390418 292170 420958 292226
rect 421014 292170 421082 292226
rect 421138 292170 451678 292226
rect 451734 292170 451802 292226
rect 451858 292170 482398 292226
rect 482454 292170 482522 292226
rect 482578 292170 513118 292226
rect 513174 292170 513242 292226
rect 513298 292170 543838 292226
rect 543894 292170 543962 292226
rect 544018 292170 574558 292226
rect 574614 292170 574682 292226
rect 574738 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 194518 292102
rect 194574 292046 194642 292102
rect 194698 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 225238 292102
rect 225294 292046 225362 292102
rect 225418 292046 255958 292102
rect 256014 292046 256082 292102
rect 256138 292046 286678 292102
rect 286734 292046 286802 292102
rect 286858 292046 317398 292102
rect 317454 292046 317522 292102
rect 317578 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 359518 292102
rect 359574 292046 359642 292102
rect 359698 292046 390238 292102
rect 390294 292046 390362 292102
rect 390418 292046 420958 292102
rect 421014 292046 421082 292102
rect 421138 292046 451678 292102
rect 451734 292046 451802 292102
rect 451858 292046 482398 292102
rect 482454 292046 482522 292102
rect 482578 292046 513118 292102
rect 513174 292046 513242 292102
rect 513298 292046 543838 292102
rect 543894 292046 543962 292102
rect 544018 292046 574558 292102
rect 574614 292046 574682 292102
rect 574738 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 194518 291978
rect 194574 291922 194642 291978
rect 194698 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 225238 291978
rect 225294 291922 225362 291978
rect 225418 291922 255958 291978
rect 256014 291922 256082 291978
rect 256138 291922 286678 291978
rect 286734 291922 286802 291978
rect 286858 291922 317398 291978
rect 317454 291922 317522 291978
rect 317578 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 359518 291978
rect 359574 291922 359642 291978
rect 359698 291922 390238 291978
rect 390294 291922 390362 291978
rect 390418 291922 420958 291978
rect 421014 291922 421082 291978
rect 421138 291922 451678 291978
rect 451734 291922 451802 291978
rect 451858 291922 482398 291978
rect 482454 291922 482522 291978
rect 482578 291922 513118 291978
rect 513174 291922 513242 291978
rect 513298 291922 543838 291978
rect 543894 291922 543962 291978
rect 544018 291922 574558 291978
rect 574614 291922 574682 291978
rect 574738 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect 188060 289018 240004 289034
rect 188060 288962 188076 289018
rect 188132 288962 239932 289018
rect 239988 288962 240004 289018
rect 188060 288946 240004 288962
rect 187052 288838 239556 288854
rect 187052 288782 187068 288838
rect 187124 288782 239484 288838
rect 239540 288782 239556 288838
rect 187052 288766 239556 288782
rect 188060 287398 236084 287414
rect 188060 287342 188076 287398
rect 188132 287342 236012 287398
rect 236068 287342 236084 287398
rect 188060 287326 236084 287342
rect 188060 285958 236308 285974
rect 188060 285902 188076 285958
rect 188132 285902 236236 285958
rect 236292 285902 236308 285958
rect 188060 285886 236308 285902
rect 187052 285778 239556 285794
rect 187052 285722 187068 285778
rect 187124 285722 239484 285778
rect 239540 285722 239556 285778
rect 187052 285706 239556 285722
rect 188060 283978 236196 283994
rect 188060 283922 188076 283978
rect 188132 283922 236124 283978
rect 236180 283922 236196 283978
rect 188060 283906 236196 283922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 59878 280350
rect 59934 280294 60002 280350
rect 60058 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 147078 280350
rect 147134 280294 147202 280350
rect 147258 280294 152902 280350
rect 152958 280294 153026 280350
rect 153082 280294 158726 280350
rect 158782 280294 158850 280350
rect 158906 280294 164550 280350
rect 164606 280294 164674 280350
rect 164730 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 209878 280350
rect 209934 280294 210002 280350
rect 210058 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 240598 280350
rect 240654 280294 240722 280350
rect 240778 280294 271318 280350
rect 271374 280294 271442 280350
rect 271498 280294 302038 280350
rect 302094 280294 302162 280350
rect 302218 280294 332758 280350
rect 332814 280294 332882 280350
rect 332938 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 374878 280350
rect 374934 280294 375002 280350
rect 375058 280294 405598 280350
rect 405654 280294 405722 280350
rect 405778 280294 436318 280350
rect 436374 280294 436442 280350
rect 436498 280294 467038 280350
rect 467094 280294 467162 280350
rect 467218 280294 497758 280350
rect 497814 280294 497882 280350
rect 497938 280294 528478 280350
rect 528534 280294 528602 280350
rect 528658 280294 559198 280350
rect 559254 280294 559322 280350
rect 559378 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 59878 280226
rect 59934 280170 60002 280226
rect 60058 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 147078 280226
rect 147134 280170 147202 280226
rect 147258 280170 152902 280226
rect 152958 280170 153026 280226
rect 153082 280170 158726 280226
rect 158782 280170 158850 280226
rect 158906 280170 164550 280226
rect 164606 280170 164674 280226
rect 164730 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 209878 280226
rect 209934 280170 210002 280226
rect 210058 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 240598 280226
rect 240654 280170 240722 280226
rect 240778 280170 271318 280226
rect 271374 280170 271442 280226
rect 271498 280170 302038 280226
rect 302094 280170 302162 280226
rect 302218 280170 332758 280226
rect 332814 280170 332882 280226
rect 332938 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 374878 280226
rect 374934 280170 375002 280226
rect 375058 280170 405598 280226
rect 405654 280170 405722 280226
rect 405778 280170 436318 280226
rect 436374 280170 436442 280226
rect 436498 280170 467038 280226
rect 467094 280170 467162 280226
rect 467218 280170 497758 280226
rect 497814 280170 497882 280226
rect 497938 280170 528478 280226
rect 528534 280170 528602 280226
rect 528658 280170 559198 280226
rect 559254 280170 559322 280226
rect 559378 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 59878 280102
rect 59934 280046 60002 280102
rect 60058 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 147078 280102
rect 147134 280046 147202 280102
rect 147258 280046 152902 280102
rect 152958 280046 153026 280102
rect 153082 280046 158726 280102
rect 158782 280046 158850 280102
rect 158906 280046 164550 280102
rect 164606 280046 164674 280102
rect 164730 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 209878 280102
rect 209934 280046 210002 280102
rect 210058 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 240598 280102
rect 240654 280046 240722 280102
rect 240778 280046 271318 280102
rect 271374 280046 271442 280102
rect 271498 280046 302038 280102
rect 302094 280046 302162 280102
rect 302218 280046 332758 280102
rect 332814 280046 332882 280102
rect 332938 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 374878 280102
rect 374934 280046 375002 280102
rect 375058 280046 405598 280102
rect 405654 280046 405722 280102
rect 405778 280046 436318 280102
rect 436374 280046 436442 280102
rect 436498 280046 467038 280102
rect 467094 280046 467162 280102
rect 467218 280046 497758 280102
rect 497814 280046 497882 280102
rect 497938 280046 528478 280102
rect 528534 280046 528602 280102
rect 528658 280046 559198 280102
rect 559254 280046 559322 280102
rect 559378 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 59878 279978
rect 59934 279922 60002 279978
rect 60058 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 147078 279978
rect 147134 279922 147202 279978
rect 147258 279922 152902 279978
rect 152958 279922 153026 279978
rect 153082 279922 158726 279978
rect 158782 279922 158850 279978
rect 158906 279922 164550 279978
rect 164606 279922 164674 279978
rect 164730 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 209878 279978
rect 209934 279922 210002 279978
rect 210058 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 240598 279978
rect 240654 279922 240722 279978
rect 240778 279922 271318 279978
rect 271374 279922 271442 279978
rect 271498 279922 302038 279978
rect 302094 279922 302162 279978
rect 302218 279922 332758 279978
rect 332814 279922 332882 279978
rect 332938 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 374878 279978
rect 374934 279922 375002 279978
rect 375058 279922 405598 279978
rect 405654 279922 405722 279978
rect 405778 279922 436318 279978
rect 436374 279922 436442 279978
rect 436498 279922 467038 279978
rect 467094 279922 467162 279978
rect 467218 279922 497758 279978
rect 497814 279922 497882 279978
rect 497938 279922 528478 279978
rect 528534 279922 528602 279978
rect 528658 279922 559198 279978
rect 559254 279922 559322 279978
rect 559378 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect 93980 275698 153764 275714
rect 93980 275642 93996 275698
rect 94052 275642 153692 275698
rect 153748 275642 153764 275698
rect 93980 275626 153764 275642
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 44518 274350
rect 44574 274294 44642 274350
rect 44698 274294 75238 274350
rect 75294 274294 75362 274350
rect 75418 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 144166 274350
rect 144222 274294 144290 274350
rect 144346 274294 149990 274350
rect 150046 274294 150114 274350
rect 150170 274294 155814 274350
rect 155870 274294 155938 274350
rect 155994 274294 161638 274350
rect 161694 274294 161762 274350
rect 161818 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 194518 274350
rect 194574 274294 194642 274350
rect 194698 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 225238 274350
rect 225294 274294 225362 274350
rect 225418 274294 255958 274350
rect 256014 274294 256082 274350
rect 256138 274294 286678 274350
rect 286734 274294 286802 274350
rect 286858 274294 317398 274350
rect 317454 274294 317522 274350
rect 317578 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 359518 274350
rect 359574 274294 359642 274350
rect 359698 274294 390238 274350
rect 390294 274294 390362 274350
rect 390418 274294 420958 274350
rect 421014 274294 421082 274350
rect 421138 274294 451678 274350
rect 451734 274294 451802 274350
rect 451858 274294 482398 274350
rect 482454 274294 482522 274350
rect 482578 274294 513118 274350
rect 513174 274294 513242 274350
rect 513298 274294 543838 274350
rect 543894 274294 543962 274350
rect 544018 274294 574558 274350
rect 574614 274294 574682 274350
rect 574738 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 44518 274226
rect 44574 274170 44642 274226
rect 44698 274170 75238 274226
rect 75294 274170 75362 274226
rect 75418 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 144166 274226
rect 144222 274170 144290 274226
rect 144346 274170 149990 274226
rect 150046 274170 150114 274226
rect 150170 274170 155814 274226
rect 155870 274170 155938 274226
rect 155994 274170 161638 274226
rect 161694 274170 161762 274226
rect 161818 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 194518 274226
rect 194574 274170 194642 274226
rect 194698 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 225238 274226
rect 225294 274170 225362 274226
rect 225418 274170 255958 274226
rect 256014 274170 256082 274226
rect 256138 274170 286678 274226
rect 286734 274170 286802 274226
rect 286858 274170 317398 274226
rect 317454 274170 317522 274226
rect 317578 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 359518 274226
rect 359574 274170 359642 274226
rect 359698 274170 390238 274226
rect 390294 274170 390362 274226
rect 390418 274170 420958 274226
rect 421014 274170 421082 274226
rect 421138 274170 451678 274226
rect 451734 274170 451802 274226
rect 451858 274170 482398 274226
rect 482454 274170 482522 274226
rect 482578 274170 513118 274226
rect 513174 274170 513242 274226
rect 513298 274170 543838 274226
rect 543894 274170 543962 274226
rect 544018 274170 574558 274226
rect 574614 274170 574682 274226
rect 574738 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 44518 274102
rect 44574 274046 44642 274102
rect 44698 274046 75238 274102
rect 75294 274046 75362 274102
rect 75418 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 144166 274102
rect 144222 274046 144290 274102
rect 144346 274046 149990 274102
rect 150046 274046 150114 274102
rect 150170 274046 155814 274102
rect 155870 274046 155938 274102
rect 155994 274046 161638 274102
rect 161694 274046 161762 274102
rect 161818 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 194518 274102
rect 194574 274046 194642 274102
rect 194698 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 225238 274102
rect 225294 274046 225362 274102
rect 225418 274046 255958 274102
rect 256014 274046 256082 274102
rect 256138 274046 286678 274102
rect 286734 274046 286802 274102
rect 286858 274046 317398 274102
rect 317454 274046 317522 274102
rect 317578 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 359518 274102
rect 359574 274046 359642 274102
rect 359698 274046 390238 274102
rect 390294 274046 390362 274102
rect 390418 274046 420958 274102
rect 421014 274046 421082 274102
rect 421138 274046 451678 274102
rect 451734 274046 451802 274102
rect 451858 274046 482398 274102
rect 482454 274046 482522 274102
rect 482578 274046 513118 274102
rect 513174 274046 513242 274102
rect 513298 274046 543838 274102
rect 543894 274046 543962 274102
rect 544018 274046 574558 274102
rect 574614 274046 574682 274102
rect 574738 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 44518 273978
rect 44574 273922 44642 273978
rect 44698 273922 75238 273978
rect 75294 273922 75362 273978
rect 75418 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 144166 273978
rect 144222 273922 144290 273978
rect 144346 273922 149990 273978
rect 150046 273922 150114 273978
rect 150170 273922 155814 273978
rect 155870 273922 155938 273978
rect 155994 273922 161638 273978
rect 161694 273922 161762 273978
rect 161818 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 194518 273978
rect 194574 273922 194642 273978
rect 194698 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 225238 273978
rect 225294 273922 225362 273978
rect 225418 273922 255958 273978
rect 256014 273922 256082 273978
rect 256138 273922 286678 273978
rect 286734 273922 286802 273978
rect 286858 273922 317398 273978
rect 317454 273922 317522 273978
rect 317578 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 359518 273978
rect 359574 273922 359642 273978
rect 359698 273922 390238 273978
rect 390294 273922 390362 273978
rect 390418 273922 420958 273978
rect 421014 273922 421082 273978
rect 421138 273922 451678 273978
rect 451734 273922 451802 273978
rect 451858 273922 482398 273978
rect 482454 273922 482522 273978
rect 482578 273922 513118 273978
rect 513174 273922 513242 273978
rect 513298 273922 543838 273978
rect 543894 273922 543962 273978
rect 544018 273922 574558 273978
rect 574614 273922 574682 273978
rect 574738 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect 229948 272098 231044 272114
rect 229948 272042 229964 272098
rect 230020 272042 230972 272098
rect 231028 272042 231044 272098
rect 229948 272026 231044 272042
rect 93980 270658 153876 270674
rect 93980 270602 93996 270658
rect 94052 270602 153804 270658
rect 153860 270602 153876 270658
rect 93980 270586 153876 270602
rect 177980 270658 236420 270674
rect 177980 270602 177996 270658
rect 178052 270602 188076 270658
rect 188132 270602 236348 270658
rect 236404 270602 236420 270658
rect 177980 270586 236420 270602
rect 153676 267058 168884 267074
rect 153676 267002 153692 267058
rect 153748 267002 168812 267058
rect 168868 267002 168884 267058
rect 153676 266986 168884 267002
rect 153788 265438 231044 265454
rect 153788 265382 153804 265438
rect 153860 265382 230972 265438
rect 231028 265382 231044 265438
rect 153788 265366 231044 265382
rect 344300 262918 353012 262934
rect 344300 262862 344316 262918
rect 344372 262862 352940 262918
rect 352996 262862 353012 262918
rect 344300 262846 353012 262862
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 59878 262350
rect 59934 262294 60002 262350
rect 60058 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 209878 262350
rect 209934 262294 210002 262350
rect 210058 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 240598 262350
rect 240654 262294 240722 262350
rect 240778 262294 271318 262350
rect 271374 262294 271442 262350
rect 271498 262294 302038 262350
rect 302094 262294 302162 262350
rect 302218 262294 332758 262350
rect 332814 262294 332882 262350
rect 332938 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 374878 262350
rect 374934 262294 375002 262350
rect 375058 262294 405598 262350
rect 405654 262294 405722 262350
rect 405778 262294 436318 262350
rect 436374 262294 436442 262350
rect 436498 262294 467038 262350
rect 467094 262294 467162 262350
rect 467218 262294 497758 262350
rect 497814 262294 497882 262350
rect 497938 262294 528478 262350
rect 528534 262294 528602 262350
rect 528658 262294 559198 262350
rect 559254 262294 559322 262350
rect 559378 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 59878 262226
rect 59934 262170 60002 262226
rect 60058 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 209878 262226
rect 209934 262170 210002 262226
rect 210058 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 240598 262226
rect 240654 262170 240722 262226
rect 240778 262170 271318 262226
rect 271374 262170 271442 262226
rect 271498 262170 302038 262226
rect 302094 262170 302162 262226
rect 302218 262170 332758 262226
rect 332814 262170 332882 262226
rect 332938 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 374878 262226
rect 374934 262170 375002 262226
rect 375058 262170 405598 262226
rect 405654 262170 405722 262226
rect 405778 262170 436318 262226
rect 436374 262170 436442 262226
rect 436498 262170 467038 262226
rect 467094 262170 467162 262226
rect 467218 262170 497758 262226
rect 497814 262170 497882 262226
rect 497938 262170 528478 262226
rect 528534 262170 528602 262226
rect 528658 262170 559198 262226
rect 559254 262170 559322 262226
rect 559378 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 59878 262102
rect 59934 262046 60002 262102
rect 60058 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 209878 262102
rect 209934 262046 210002 262102
rect 210058 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 240598 262102
rect 240654 262046 240722 262102
rect 240778 262046 271318 262102
rect 271374 262046 271442 262102
rect 271498 262046 302038 262102
rect 302094 262046 302162 262102
rect 302218 262046 332758 262102
rect 332814 262046 332882 262102
rect 332938 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 374878 262102
rect 374934 262046 375002 262102
rect 375058 262046 405598 262102
rect 405654 262046 405722 262102
rect 405778 262046 436318 262102
rect 436374 262046 436442 262102
rect 436498 262046 467038 262102
rect 467094 262046 467162 262102
rect 467218 262046 497758 262102
rect 497814 262046 497882 262102
rect 497938 262046 528478 262102
rect 528534 262046 528602 262102
rect 528658 262046 559198 262102
rect 559254 262046 559322 262102
rect 559378 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 59878 261978
rect 59934 261922 60002 261978
rect 60058 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 209878 261978
rect 209934 261922 210002 261978
rect 210058 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 240598 261978
rect 240654 261922 240722 261978
rect 240778 261922 271318 261978
rect 271374 261922 271442 261978
rect 271498 261922 302038 261978
rect 302094 261922 302162 261978
rect 302218 261922 332758 261978
rect 332814 261922 332882 261978
rect 332938 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 374878 261978
rect 374934 261922 375002 261978
rect 375058 261922 405598 261978
rect 405654 261922 405722 261978
rect 405778 261922 436318 261978
rect 436374 261922 436442 261978
rect 436498 261922 467038 261978
rect 467094 261922 467162 261978
rect 467218 261922 497758 261978
rect 497814 261922 497882 261978
rect 497938 261922 528478 261978
rect 528534 261922 528602 261978
rect 528658 261922 559198 261978
rect 559254 261922 559322 261978
rect 559378 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect 190636 260398 239444 260414
rect 190636 260342 190652 260398
rect 190708 260342 239372 260398
rect 239428 260342 239444 260398
rect 190636 260326 239444 260342
rect 338588 258418 339348 258434
rect 338588 258362 338604 258418
rect 338660 258362 339276 258418
rect 339332 258362 339348 258418
rect 338588 258346 339348 258362
rect 338700 256618 339460 256634
rect 338700 256562 338716 256618
rect 338772 256562 339388 256618
rect 339444 256562 339460 256618
rect 338700 256546 339460 256562
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 44518 256350
rect 44574 256294 44642 256350
rect 44698 256294 75238 256350
rect 75294 256294 75362 256350
rect 75418 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 194518 256350
rect 194574 256294 194642 256350
rect 194698 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 225238 256350
rect 225294 256294 225362 256350
rect 225418 256294 255958 256350
rect 256014 256294 256082 256350
rect 256138 256294 286678 256350
rect 286734 256294 286802 256350
rect 286858 256294 317398 256350
rect 317454 256294 317522 256350
rect 317578 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 359518 256350
rect 359574 256294 359642 256350
rect 359698 256294 390238 256350
rect 390294 256294 390362 256350
rect 390418 256294 420958 256350
rect 421014 256294 421082 256350
rect 421138 256294 451678 256350
rect 451734 256294 451802 256350
rect 451858 256294 482398 256350
rect 482454 256294 482522 256350
rect 482578 256294 513118 256350
rect 513174 256294 513242 256350
rect 513298 256294 543838 256350
rect 543894 256294 543962 256350
rect 544018 256294 574558 256350
rect 574614 256294 574682 256350
rect 574738 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 44518 256226
rect 44574 256170 44642 256226
rect 44698 256170 75238 256226
rect 75294 256170 75362 256226
rect 75418 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 194518 256226
rect 194574 256170 194642 256226
rect 194698 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 225238 256226
rect 225294 256170 225362 256226
rect 225418 256170 255958 256226
rect 256014 256170 256082 256226
rect 256138 256170 286678 256226
rect 286734 256170 286802 256226
rect 286858 256170 317398 256226
rect 317454 256170 317522 256226
rect 317578 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 359518 256226
rect 359574 256170 359642 256226
rect 359698 256170 390238 256226
rect 390294 256170 390362 256226
rect 390418 256170 420958 256226
rect 421014 256170 421082 256226
rect 421138 256170 451678 256226
rect 451734 256170 451802 256226
rect 451858 256170 482398 256226
rect 482454 256170 482522 256226
rect 482578 256170 513118 256226
rect 513174 256170 513242 256226
rect 513298 256170 543838 256226
rect 543894 256170 543962 256226
rect 544018 256170 574558 256226
rect 574614 256170 574682 256226
rect 574738 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 44518 256102
rect 44574 256046 44642 256102
rect 44698 256046 75238 256102
rect 75294 256046 75362 256102
rect 75418 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 194518 256102
rect 194574 256046 194642 256102
rect 194698 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 225238 256102
rect 225294 256046 225362 256102
rect 225418 256046 255958 256102
rect 256014 256046 256082 256102
rect 256138 256046 286678 256102
rect 286734 256046 286802 256102
rect 286858 256046 317398 256102
rect 317454 256046 317522 256102
rect 317578 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 359518 256102
rect 359574 256046 359642 256102
rect 359698 256046 390238 256102
rect 390294 256046 390362 256102
rect 390418 256046 420958 256102
rect 421014 256046 421082 256102
rect 421138 256046 451678 256102
rect 451734 256046 451802 256102
rect 451858 256046 482398 256102
rect 482454 256046 482522 256102
rect 482578 256046 513118 256102
rect 513174 256046 513242 256102
rect 513298 256046 543838 256102
rect 543894 256046 543962 256102
rect 544018 256046 574558 256102
rect 574614 256046 574682 256102
rect 574738 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 44518 255978
rect 44574 255922 44642 255978
rect 44698 255922 75238 255978
rect 75294 255922 75362 255978
rect 75418 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 194518 255978
rect 194574 255922 194642 255978
rect 194698 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 225238 255978
rect 225294 255922 225362 255978
rect 225418 255922 255958 255978
rect 256014 255922 256082 255978
rect 256138 255922 286678 255978
rect 286734 255922 286802 255978
rect 286858 255922 317398 255978
rect 317454 255922 317522 255978
rect 317578 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 359518 255978
rect 359574 255922 359642 255978
rect 359698 255922 390238 255978
rect 390294 255922 390362 255978
rect 390418 255922 420958 255978
rect 421014 255922 421082 255978
rect 421138 255922 451678 255978
rect 451734 255922 451802 255978
rect 451858 255922 482398 255978
rect 482454 255922 482522 255978
rect 482578 255922 513118 255978
rect 513174 255922 513242 255978
rect 513298 255922 543838 255978
rect 543894 255922 543962 255978
rect 544018 255922 574558 255978
rect 574614 255922 574682 255978
rect 574738 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect 190636 255538 241124 255554
rect 190636 255482 190652 255538
rect 190708 255482 241052 255538
rect 241108 255482 241124 255538
rect 190636 255466 241124 255482
rect 338364 253738 339348 253754
rect 338364 253682 338380 253738
rect 338436 253682 339276 253738
rect 339332 253682 339348 253738
rect 338364 253666 339348 253682
rect 190636 252118 239444 252134
rect 190636 252062 190652 252118
rect 190708 252062 239372 252118
rect 239428 252062 239444 252118
rect 190636 252046 239444 252062
rect 174620 251218 241236 251234
rect 174620 251162 174636 251218
rect 174692 251162 241164 251218
rect 241220 251162 241236 251218
rect 174620 251146 241236 251162
rect 338364 249958 340132 249974
rect 338364 249902 338380 249958
rect 338436 249902 340060 249958
rect 340116 249902 340132 249958
rect 338364 249886 340132 249902
rect 338476 247078 339348 247094
rect 338476 247022 338492 247078
rect 338548 247022 339276 247078
rect 339332 247022 339348 247078
rect 338476 247006 339348 247022
rect 338252 245458 339460 245474
rect 338252 245402 338268 245458
rect 338324 245402 339388 245458
rect 339444 245402 339460 245458
rect 338252 245386 339460 245402
rect 338476 245098 339460 245114
rect 338476 245042 338492 245098
rect 338548 245042 339388 245098
rect 339444 245042 339460 245098
rect 338476 245026 339460 245042
rect 337916 244918 339460 244934
rect 337916 244862 337932 244918
rect 337988 244862 339388 244918
rect 339444 244862 339460 244918
rect 337916 244846 339460 244862
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 59878 244350
rect 59934 244294 60002 244350
rect 60058 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 209878 244350
rect 209934 244294 210002 244350
rect 210058 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 240598 244350
rect 240654 244294 240722 244350
rect 240778 244294 271318 244350
rect 271374 244294 271442 244350
rect 271498 244294 302038 244350
rect 302094 244294 302162 244350
rect 302218 244294 332758 244350
rect 332814 244294 332882 244350
rect 332938 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 374878 244350
rect 374934 244294 375002 244350
rect 375058 244294 405598 244350
rect 405654 244294 405722 244350
rect 405778 244294 436318 244350
rect 436374 244294 436442 244350
rect 436498 244294 467038 244350
rect 467094 244294 467162 244350
rect 467218 244294 497758 244350
rect 497814 244294 497882 244350
rect 497938 244294 528478 244350
rect 528534 244294 528602 244350
rect 528658 244294 559198 244350
rect 559254 244294 559322 244350
rect 559378 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 59878 244226
rect 59934 244170 60002 244226
rect 60058 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 209878 244226
rect 209934 244170 210002 244226
rect 210058 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 240598 244226
rect 240654 244170 240722 244226
rect 240778 244170 271318 244226
rect 271374 244170 271442 244226
rect 271498 244170 302038 244226
rect 302094 244170 302162 244226
rect 302218 244170 332758 244226
rect 332814 244170 332882 244226
rect 332938 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 374878 244226
rect 374934 244170 375002 244226
rect 375058 244170 405598 244226
rect 405654 244170 405722 244226
rect 405778 244170 436318 244226
rect 436374 244170 436442 244226
rect 436498 244170 467038 244226
rect 467094 244170 467162 244226
rect 467218 244170 497758 244226
rect 497814 244170 497882 244226
rect 497938 244170 528478 244226
rect 528534 244170 528602 244226
rect 528658 244170 559198 244226
rect 559254 244170 559322 244226
rect 559378 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 59878 244102
rect 59934 244046 60002 244102
rect 60058 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 209878 244102
rect 209934 244046 210002 244102
rect 210058 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 240598 244102
rect 240654 244046 240722 244102
rect 240778 244046 271318 244102
rect 271374 244046 271442 244102
rect 271498 244046 302038 244102
rect 302094 244046 302162 244102
rect 302218 244046 332758 244102
rect 332814 244046 332882 244102
rect 332938 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 374878 244102
rect 374934 244046 375002 244102
rect 375058 244046 405598 244102
rect 405654 244046 405722 244102
rect 405778 244046 436318 244102
rect 436374 244046 436442 244102
rect 436498 244046 467038 244102
rect 467094 244046 467162 244102
rect 467218 244046 497758 244102
rect 497814 244046 497882 244102
rect 497938 244046 528478 244102
rect 528534 244046 528602 244102
rect 528658 244046 559198 244102
rect 559254 244046 559322 244102
rect 559378 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 59878 243978
rect 59934 243922 60002 243978
rect 60058 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 209878 243978
rect 209934 243922 210002 243978
rect 210058 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 240598 243978
rect 240654 243922 240722 243978
rect 240778 243922 271318 243978
rect 271374 243922 271442 243978
rect 271498 243922 302038 243978
rect 302094 243922 302162 243978
rect 302218 243922 332758 243978
rect 332814 243922 332882 243978
rect 332938 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 374878 243978
rect 374934 243922 375002 243978
rect 375058 243922 405598 243978
rect 405654 243922 405722 243978
rect 405778 243922 436318 243978
rect 436374 243922 436442 243978
rect 436498 243922 467038 243978
rect 467094 243922 467162 243978
rect 467218 243922 497758 243978
rect 497814 243922 497882 243978
rect 497938 243922 528478 243978
rect 528534 243922 528602 243978
rect 528658 243922 559198 243978
rect 559254 243922 559322 243978
rect 559378 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect 241148 241858 344836 241874
rect 241148 241802 241164 241858
rect 241220 241802 344764 241858
rect 344820 241802 344836 241858
rect 241148 241786 344836 241802
rect 236332 241678 339796 241694
rect 236332 241622 236348 241678
rect 236404 241622 339724 241678
rect 339780 241622 339796 241678
rect 236332 241606 339796 241622
rect 336908 241498 341364 241514
rect 336908 241442 336924 241498
rect 336980 241442 341292 241498
rect 341348 241442 341364 241498
rect 336908 241426 341364 241442
rect 337244 241318 342484 241334
rect 337244 241262 337260 241318
rect 337316 241262 342412 241318
rect 342468 241262 342484 241318
rect 337244 241246 342484 241262
rect 289756 241138 342932 241154
rect 289756 241082 289772 241138
rect 289828 241082 342860 241138
rect 342916 241082 342932 241138
rect 289756 241066 342932 241082
rect 344748 240418 345620 240434
rect 344748 240362 344764 240418
rect 344820 240362 345548 240418
rect 345604 240362 345620 240418
rect 344748 240346 345620 240362
rect 337132 240238 339684 240254
rect 337132 240182 337148 240238
rect 337204 240182 339612 240238
rect 339668 240182 339684 240238
rect 337132 240166 339684 240182
rect 18380 238978 342708 238994
rect 18380 238922 18396 238978
rect 18452 238922 342636 238978
rect 342692 238922 342708 238978
rect 18380 238906 342708 238922
rect 16700 238798 340020 238814
rect 16700 238742 16716 238798
rect 16772 238742 339948 238798
rect 340004 238742 340020 238798
rect 16700 238726 340020 238742
rect 336796 238618 340916 238634
rect 336796 238562 336812 238618
rect 336868 238562 340844 238618
rect 340900 238562 340916 238618
rect 336796 238546 340916 238562
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 359518 238350
rect 359574 238294 359642 238350
rect 359698 238294 390238 238350
rect 390294 238294 390362 238350
rect 390418 238294 420958 238350
rect 421014 238294 421082 238350
rect 421138 238294 451678 238350
rect 451734 238294 451802 238350
rect 451858 238294 482398 238350
rect 482454 238294 482522 238350
rect 482578 238294 513118 238350
rect 513174 238294 513242 238350
rect 513298 238294 543838 238350
rect 543894 238294 543962 238350
rect 544018 238294 574558 238350
rect 574614 238294 574682 238350
rect 574738 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 359518 238226
rect 359574 238170 359642 238226
rect 359698 238170 390238 238226
rect 390294 238170 390362 238226
rect 390418 238170 420958 238226
rect 421014 238170 421082 238226
rect 421138 238170 451678 238226
rect 451734 238170 451802 238226
rect 451858 238170 482398 238226
rect 482454 238170 482522 238226
rect 482578 238170 513118 238226
rect 513174 238170 513242 238226
rect 513298 238170 543838 238226
rect 543894 238170 543962 238226
rect 544018 238170 574558 238226
rect 574614 238170 574682 238226
rect 574738 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 359518 238102
rect 359574 238046 359642 238102
rect 359698 238046 390238 238102
rect 390294 238046 390362 238102
rect 390418 238046 420958 238102
rect 421014 238046 421082 238102
rect 421138 238046 451678 238102
rect 451734 238046 451802 238102
rect 451858 238046 482398 238102
rect 482454 238046 482522 238102
rect 482578 238046 513118 238102
rect 513174 238046 513242 238102
rect 513298 238046 543838 238102
rect 543894 238046 543962 238102
rect 544018 238046 574558 238102
rect 574614 238046 574682 238102
rect 574738 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 359518 237978
rect 359574 237922 359642 237978
rect 359698 237922 390238 237978
rect 390294 237922 390362 237978
rect 390418 237922 420958 237978
rect 421014 237922 421082 237978
rect 421138 237922 451678 237978
rect 451734 237922 451802 237978
rect 451858 237922 482398 237978
rect 482454 237922 482522 237978
rect 482578 237922 513118 237978
rect 513174 237922 513242 237978
rect 513298 237922 543838 237978
rect 543894 237922 543962 237978
rect 544018 237922 574558 237978
rect 574614 237922 574682 237978
rect 574738 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect 62620 237718 170564 237734
rect 62620 237662 62636 237718
rect 62692 237662 170492 237718
rect 170548 237662 170564 237718
rect 62620 237646 170564 237662
rect 64412 237538 100228 237554
rect 64412 237482 64428 237538
rect 64484 237482 100156 237538
rect 100212 237482 100228 237538
rect 64412 237466 100228 237482
rect 245068 237178 269908 237194
rect 245068 237122 245084 237178
rect 245140 237122 269836 237178
rect 269892 237122 269908 237178
rect 245068 237106 269908 237122
rect 244172 236998 277300 237014
rect 244172 236942 244188 236998
rect 244244 236942 277228 236998
rect 277284 236942 277300 236998
rect 244172 236926 277300 236942
rect 355388 236638 356708 236654
rect 355388 236582 355404 236638
rect 355460 236582 356636 236638
rect 356692 236582 356708 236638
rect 355388 236566 356708 236582
rect 239804 234658 353572 234674
rect 239804 234602 239820 234658
rect 239876 234602 353500 234658
rect 353556 234602 353572 234658
rect 239804 234586 353572 234602
rect 21740 234478 340132 234494
rect 21740 234422 21756 234478
rect 21812 234422 340060 234478
rect 340116 234422 340132 234478
rect 21740 234406 340132 234422
rect 26780 234298 346180 234314
rect 26780 234242 26796 234298
rect 26852 234242 346108 234298
rect 346164 234242 346180 234298
rect 26780 234226 346180 234242
rect 236668 231418 270020 231434
rect 236668 231362 236684 231418
rect 236740 231362 269948 231418
rect 270004 231362 270020 231418
rect 236668 231346 270020 231362
rect 236780 231238 269796 231254
rect 236780 231182 236796 231238
rect 236852 231182 269724 231238
rect 269780 231182 269796 231238
rect 236780 231166 269796 231182
rect 209900 231058 267220 231074
rect 209900 231002 209916 231058
rect 209972 231002 267148 231058
rect 267204 231002 267220 231058
rect 209900 230986 267220 231002
rect 241820 227998 270804 228014
rect 241820 227942 241836 227998
rect 241892 227942 270732 227998
rect 270788 227942 270804 227998
rect 241820 227926 270804 227942
rect 240028 227818 270916 227834
rect 240028 227762 240044 227818
rect 240100 227762 270844 227818
rect 270900 227762 270916 227818
rect 240028 227746 270916 227762
rect 238460 227638 271028 227654
rect 238460 227582 238476 227638
rect 238532 227582 270956 227638
rect 271012 227582 271028 227638
rect 238460 227566 271028 227582
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 374878 226350
rect 374934 226294 375002 226350
rect 375058 226294 405598 226350
rect 405654 226294 405722 226350
rect 405778 226294 436318 226350
rect 436374 226294 436442 226350
rect 436498 226294 467038 226350
rect 467094 226294 467162 226350
rect 467218 226294 497758 226350
rect 497814 226294 497882 226350
rect 497938 226294 528478 226350
rect 528534 226294 528602 226350
rect 528658 226294 559198 226350
rect 559254 226294 559322 226350
rect 559378 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 374878 226226
rect 374934 226170 375002 226226
rect 375058 226170 405598 226226
rect 405654 226170 405722 226226
rect 405778 226170 436318 226226
rect 436374 226170 436442 226226
rect 436498 226170 467038 226226
rect 467094 226170 467162 226226
rect 467218 226170 497758 226226
rect 497814 226170 497882 226226
rect 497938 226170 528478 226226
rect 528534 226170 528602 226226
rect 528658 226170 559198 226226
rect 559254 226170 559322 226226
rect 559378 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 374878 226102
rect 374934 226046 375002 226102
rect 375058 226046 405598 226102
rect 405654 226046 405722 226102
rect 405778 226046 436318 226102
rect 436374 226046 436442 226102
rect 436498 226046 467038 226102
rect 467094 226046 467162 226102
rect 467218 226046 497758 226102
rect 497814 226046 497882 226102
rect 497938 226046 528478 226102
rect 528534 226046 528602 226102
rect 528658 226046 559198 226102
rect 559254 226046 559322 226102
rect 559378 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 374878 225978
rect 374934 225922 375002 225978
rect 375058 225922 405598 225978
rect 405654 225922 405722 225978
rect 405778 225922 436318 225978
rect 436374 225922 436442 225978
rect 436498 225922 467038 225978
rect 467094 225922 467162 225978
rect 467218 225922 497758 225978
rect 497814 225922 497882 225978
rect 497938 225922 528478 225978
rect 528534 225922 528602 225978
rect 528658 225922 559198 225978
rect 559254 225922 559322 225978
rect 559378 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect 243388 224578 267444 224594
rect 243388 224522 243404 224578
rect 243460 224522 267372 224578
rect 267428 224522 267444 224578
rect 243388 224506 267444 224522
rect 243500 224398 275620 224414
rect 243500 224342 243516 224398
rect 243572 224342 275548 224398
rect 275604 224342 275620 224398
rect 243500 224326 275620 224342
rect 33388 224218 225220 224234
rect 33388 224162 33404 224218
rect 33460 224162 225148 224218
rect 225204 224162 225220 224218
rect 33388 224146 225220 224162
rect 233420 224218 273940 224234
rect 233420 224162 233436 224218
rect 233492 224162 273868 224218
rect 273924 224162 273940 224218
rect 233420 224146 273940 224162
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 359518 220350
rect 359574 220294 359642 220350
rect 359698 220294 390238 220350
rect 390294 220294 390362 220350
rect 390418 220294 420958 220350
rect 421014 220294 421082 220350
rect 421138 220294 451678 220350
rect 451734 220294 451802 220350
rect 451858 220294 482398 220350
rect 482454 220294 482522 220350
rect 482578 220294 513118 220350
rect 513174 220294 513242 220350
rect 513298 220294 543838 220350
rect 543894 220294 543962 220350
rect 544018 220294 574558 220350
rect 574614 220294 574682 220350
rect 574738 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 359518 220226
rect 359574 220170 359642 220226
rect 359698 220170 390238 220226
rect 390294 220170 390362 220226
rect 390418 220170 420958 220226
rect 421014 220170 421082 220226
rect 421138 220170 451678 220226
rect 451734 220170 451802 220226
rect 451858 220170 482398 220226
rect 482454 220170 482522 220226
rect 482578 220170 513118 220226
rect 513174 220170 513242 220226
rect 513298 220170 543838 220226
rect 543894 220170 543962 220226
rect 544018 220170 574558 220226
rect 574614 220170 574682 220226
rect 574738 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 359518 220102
rect 359574 220046 359642 220102
rect 359698 220046 390238 220102
rect 390294 220046 390362 220102
rect 390418 220046 420958 220102
rect 421014 220046 421082 220102
rect 421138 220046 451678 220102
rect 451734 220046 451802 220102
rect 451858 220046 482398 220102
rect 482454 220046 482522 220102
rect 482578 220046 513118 220102
rect 513174 220046 513242 220102
rect 513298 220046 543838 220102
rect 543894 220046 543962 220102
rect 544018 220046 574558 220102
rect 574614 220046 574682 220102
rect 574738 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 359518 219978
rect 359574 219922 359642 219978
rect 359698 219922 390238 219978
rect 390294 219922 390362 219978
rect 390418 219922 420958 219978
rect 421014 219922 421082 219978
rect 421138 219922 451678 219978
rect 451734 219922 451802 219978
rect 451858 219922 482398 219978
rect 482454 219922 482522 219978
rect 482578 219922 513118 219978
rect 513174 219922 513242 219978
rect 513298 219922 543838 219978
rect 543894 219922 543962 219978
rect 544018 219922 574558 219978
rect 574614 219922 574682 219978
rect 574738 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect 355388 213598 356820 213614
rect 355388 213542 355404 213598
rect 355460 213542 356748 213598
rect 356804 213542 356820 213598
rect 355388 213526 356820 213542
rect 239580 211438 267668 211454
rect 239580 211382 239596 211438
rect 239652 211382 267596 211438
rect 267652 211382 267668 211438
rect 239580 211366 267668 211382
rect 240140 211258 269236 211274
rect 240140 211202 240156 211258
rect 240212 211202 269164 211258
rect 269220 211202 269236 211258
rect 240140 211186 269236 211202
rect 241036 211078 345844 211094
rect 241036 211022 241052 211078
rect 241108 211022 345772 211078
rect 345828 211022 345844 211078
rect 241036 211006 345844 211022
rect 184476 210898 339796 210914
rect 184476 210842 184492 210898
rect 184548 210842 339724 210898
rect 339780 210842 339796 210898
rect 184476 210826 339796 210842
rect 41116 210178 274164 210194
rect 41116 210122 41132 210178
rect 41188 210122 274092 210178
rect 274148 210122 274164 210178
rect 41116 210106 274164 210122
rect 267020 209098 298244 209114
rect 267020 209042 267036 209098
rect 267092 209042 298172 209098
rect 298228 209042 298244 209098
rect 267020 209026 298244 209042
rect 41452 208738 274276 208754
rect 41452 208682 41468 208738
rect 41524 208682 274204 208738
rect 274260 208682 274276 208738
rect 41452 208666 274276 208682
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 374878 208350
rect 374934 208294 375002 208350
rect 375058 208294 405598 208350
rect 405654 208294 405722 208350
rect 405778 208294 436318 208350
rect 436374 208294 436442 208350
rect 436498 208294 467038 208350
rect 467094 208294 467162 208350
rect 467218 208294 497758 208350
rect 497814 208294 497882 208350
rect 497938 208294 528478 208350
rect 528534 208294 528602 208350
rect 528658 208294 559198 208350
rect 559254 208294 559322 208350
rect 559378 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 374878 208226
rect 374934 208170 375002 208226
rect 375058 208170 405598 208226
rect 405654 208170 405722 208226
rect 405778 208170 436318 208226
rect 436374 208170 436442 208226
rect 436498 208170 467038 208226
rect 467094 208170 467162 208226
rect 467218 208170 497758 208226
rect 497814 208170 497882 208226
rect 497938 208170 528478 208226
rect 528534 208170 528602 208226
rect 528658 208170 559198 208226
rect 559254 208170 559322 208226
rect 559378 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 374878 208102
rect 374934 208046 375002 208102
rect 375058 208046 405598 208102
rect 405654 208046 405722 208102
rect 405778 208046 436318 208102
rect 436374 208046 436442 208102
rect 436498 208046 467038 208102
rect 467094 208046 467162 208102
rect 467218 208046 497758 208102
rect 497814 208046 497882 208102
rect 497938 208046 528478 208102
rect 528534 208046 528602 208102
rect 528658 208046 559198 208102
rect 559254 208046 559322 208102
rect 559378 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 374878 207978
rect 374934 207922 375002 207978
rect 375058 207922 405598 207978
rect 405654 207922 405722 207978
rect 405778 207922 436318 207978
rect 436374 207922 436442 207978
rect 436498 207922 467038 207978
rect 467094 207922 467162 207978
rect 467218 207922 497758 207978
rect 497814 207922 497882 207978
rect 497938 207922 528478 207978
rect 528534 207922 528602 207978
rect 528658 207922 559198 207978
rect 559254 207922 559322 207978
rect 559378 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 44518 202350
rect 44574 202294 44642 202350
rect 44698 202294 75238 202350
rect 75294 202294 75362 202350
rect 75418 202294 105958 202350
rect 106014 202294 106082 202350
rect 106138 202294 136678 202350
rect 136734 202294 136802 202350
rect 136858 202294 167398 202350
rect 167454 202294 167522 202350
rect 167578 202294 198118 202350
rect 198174 202294 198242 202350
rect 198298 202294 228838 202350
rect 228894 202294 228962 202350
rect 229018 202294 259558 202350
rect 259614 202294 259682 202350
rect 259738 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 359518 202350
rect 359574 202294 359642 202350
rect 359698 202294 390238 202350
rect 390294 202294 390362 202350
rect 390418 202294 420958 202350
rect 421014 202294 421082 202350
rect 421138 202294 451678 202350
rect 451734 202294 451802 202350
rect 451858 202294 482398 202350
rect 482454 202294 482522 202350
rect 482578 202294 513118 202350
rect 513174 202294 513242 202350
rect 513298 202294 543838 202350
rect 543894 202294 543962 202350
rect 544018 202294 574558 202350
rect 574614 202294 574682 202350
rect 574738 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 44518 202226
rect 44574 202170 44642 202226
rect 44698 202170 75238 202226
rect 75294 202170 75362 202226
rect 75418 202170 105958 202226
rect 106014 202170 106082 202226
rect 106138 202170 136678 202226
rect 136734 202170 136802 202226
rect 136858 202170 167398 202226
rect 167454 202170 167522 202226
rect 167578 202170 198118 202226
rect 198174 202170 198242 202226
rect 198298 202170 228838 202226
rect 228894 202170 228962 202226
rect 229018 202170 259558 202226
rect 259614 202170 259682 202226
rect 259738 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 359518 202226
rect 359574 202170 359642 202226
rect 359698 202170 390238 202226
rect 390294 202170 390362 202226
rect 390418 202170 420958 202226
rect 421014 202170 421082 202226
rect 421138 202170 451678 202226
rect 451734 202170 451802 202226
rect 451858 202170 482398 202226
rect 482454 202170 482522 202226
rect 482578 202170 513118 202226
rect 513174 202170 513242 202226
rect 513298 202170 543838 202226
rect 543894 202170 543962 202226
rect 544018 202170 574558 202226
rect 574614 202170 574682 202226
rect 574738 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 44518 202102
rect 44574 202046 44642 202102
rect 44698 202046 75238 202102
rect 75294 202046 75362 202102
rect 75418 202046 105958 202102
rect 106014 202046 106082 202102
rect 106138 202046 136678 202102
rect 136734 202046 136802 202102
rect 136858 202046 167398 202102
rect 167454 202046 167522 202102
rect 167578 202046 198118 202102
rect 198174 202046 198242 202102
rect 198298 202046 228838 202102
rect 228894 202046 228962 202102
rect 229018 202046 259558 202102
rect 259614 202046 259682 202102
rect 259738 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 359518 202102
rect 359574 202046 359642 202102
rect 359698 202046 390238 202102
rect 390294 202046 390362 202102
rect 390418 202046 420958 202102
rect 421014 202046 421082 202102
rect 421138 202046 451678 202102
rect 451734 202046 451802 202102
rect 451858 202046 482398 202102
rect 482454 202046 482522 202102
rect 482578 202046 513118 202102
rect 513174 202046 513242 202102
rect 513298 202046 543838 202102
rect 543894 202046 543962 202102
rect 544018 202046 574558 202102
rect 574614 202046 574682 202102
rect 574738 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 44518 201978
rect 44574 201922 44642 201978
rect 44698 201922 75238 201978
rect 75294 201922 75362 201978
rect 75418 201922 105958 201978
rect 106014 201922 106082 201978
rect 106138 201922 136678 201978
rect 136734 201922 136802 201978
rect 136858 201922 167398 201978
rect 167454 201922 167522 201978
rect 167578 201922 198118 201978
rect 198174 201922 198242 201978
rect 198298 201922 228838 201978
rect 228894 201922 228962 201978
rect 229018 201922 259558 201978
rect 259614 201922 259682 201978
rect 259738 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 359518 201978
rect 359574 201922 359642 201978
rect 359698 201922 390238 201978
rect 390294 201922 390362 201978
rect 390418 201922 420958 201978
rect 421014 201922 421082 201978
rect 421138 201922 451678 201978
rect 451734 201922 451802 201978
rect 451858 201922 482398 201978
rect 482454 201922 482522 201978
rect 482578 201922 513118 201978
rect 513174 201922 513242 201978
rect 513298 201922 543838 201978
rect 543894 201922 543962 201978
rect 544018 201922 574558 201978
rect 574614 201922 574682 201978
rect 574738 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect 309020 197578 338452 197594
rect 309020 197522 309036 197578
rect 309092 197522 338380 197578
rect 338436 197522 338452 197578
rect 309020 197506 338452 197522
rect 310700 197398 344164 197414
rect 310700 197342 310716 197398
rect 310772 197342 344092 197398
rect 344148 197342 344164 197398
rect 310700 197326 344164 197342
rect 319100 193978 340356 193994
rect 319100 193922 319116 193978
rect 319172 193922 340284 193978
rect 340340 193922 340356 193978
rect 319100 193906 340356 193922
rect 334220 192358 341140 192374
rect 334220 192302 334236 192358
rect 334292 192302 341068 192358
rect 341124 192302 341140 192358
rect 334220 192286 341140 192302
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 59878 190350
rect 59934 190294 60002 190350
rect 60058 190294 90598 190350
rect 90654 190294 90722 190350
rect 90778 190294 121318 190350
rect 121374 190294 121442 190350
rect 121498 190294 152038 190350
rect 152094 190294 152162 190350
rect 152218 190294 182758 190350
rect 182814 190294 182882 190350
rect 182938 190294 213478 190350
rect 213534 190294 213602 190350
rect 213658 190294 244198 190350
rect 244254 190294 244322 190350
rect 244378 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 309822 190350
rect 309878 190294 309946 190350
rect 310002 190294 318390 190350
rect 318446 190294 318514 190350
rect 318570 190294 326958 190350
rect 327014 190294 327082 190350
rect 327138 190294 335526 190350
rect 335582 190294 335650 190350
rect 335706 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 374878 190350
rect 374934 190294 375002 190350
rect 375058 190294 405598 190350
rect 405654 190294 405722 190350
rect 405778 190294 436318 190350
rect 436374 190294 436442 190350
rect 436498 190294 467038 190350
rect 467094 190294 467162 190350
rect 467218 190294 497758 190350
rect 497814 190294 497882 190350
rect 497938 190294 528478 190350
rect 528534 190294 528602 190350
rect 528658 190294 559198 190350
rect 559254 190294 559322 190350
rect 559378 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 59878 190226
rect 59934 190170 60002 190226
rect 60058 190170 90598 190226
rect 90654 190170 90722 190226
rect 90778 190170 121318 190226
rect 121374 190170 121442 190226
rect 121498 190170 152038 190226
rect 152094 190170 152162 190226
rect 152218 190170 182758 190226
rect 182814 190170 182882 190226
rect 182938 190170 213478 190226
rect 213534 190170 213602 190226
rect 213658 190170 244198 190226
rect 244254 190170 244322 190226
rect 244378 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 309822 190226
rect 309878 190170 309946 190226
rect 310002 190170 318390 190226
rect 318446 190170 318514 190226
rect 318570 190170 326958 190226
rect 327014 190170 327082 190226
rect 327138 190170 335526 190226
rect 335582 190170 335650 190226
rect 335706 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 374878 190226
rect 374934 190170 375002 190226
rect 375058 190170 405598 190226
rect 405654 190170 405722 190226
rect 405778 190170 436318 190226
rect 436374 190170 436442 190226
rect 436498 190170 467038 190226
rect 467094 190170 467162 190226
rect 467218 190170 497758 190226
rect 497814 190170 497882 190226
rect 497938 190170 528478 190226
rect 528534 190170 528602 190226
rect 528658 190170 559198 190226
rect 559254 190170 559322 190226
rect 559378 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 59878 190102
rect 59934 190046 60002 190102
rect 60058 190046 90598 190102
rect 90654 190046 90722 190102
rect 90778 190046 121318 190102
rect 121374 190046 121442 190102
rect 121498 190046 152038 190102
rect 152094 190046 152162 190102
rect 152218 190046 182758 190102
rect 182814 190046 182882 190102
rect 182938 190046 213478 190102
rect 213534 190046 213602 190102
rect 213658 190046 244198 190102
rect 244254 190046 244322 190102
rect 244378 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 309822 190102
rect 309878 190046 309946 190102
rect 310002 190046 318390 190102
rect 318446 190046 318514 190102
rect 318570 190046 326958 190102
rect 327014 190046 327082 190102
rect 327138 190046 335526 190102
rect 335582 190046 335650 190102
rect 335706 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 374878 190102
rect 374934 190046 375002 190102
rect 375058 190046 405598 190102
rect 405654 190046 405722 190102
rect 405778 190046 436318 190102
rect 436374 190046 436442 190102
rect 436498 190046 467038 190102
rect 467094 190046 467162 190102
rect 467218 190046 497758 190102
rect 497814 190046 497882 190102
rect 497938 190046 528478 190102
rect 528534 190046 528602 190102
rect 528658 190046 559198 190102
rect 559254 190046 559322 190102
rect 559378 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 59878 189978
rect 59934 189922 60002 189978
rect 60058 189922 90598 189978
rect 90654 189922 90722 189978
rect 90778 189922 121318 189978
rect 121374 189922 121442 189978
rect 121498 189922 152038 189978
rect 152094 189922 152162 189978
rect 152218 189922 182758 189978
rect 182814 189922 182882 189978
rect 182938 189922 213478 189978
rect 213534 189922 213602 189978
rect 213658 189922 244198 189978
rect 244254 189922 244322 189978
rect 244378 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 309822 189978
rect 309878 189922 309946 189978
rect 310002 189922 318390 189978
rect 318446 189922 318514 189978
rect 318570 189922 326958 189978
rect 327014 189922 327082 189978
rect 327138 189922 335526 189978
rect 335582 189922 335650 189978
rect 335706 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 374878 189978
rect 374934 189922 375002 189978
rect 375058 189922 405598 189978
rect 405654 189922 405722 189978
rect 405778 189922 436318 189978
rect 436374 189922 436442 189978
rect 436498 189922 467038 189978
rect 467094 189922 467162 189978
rect 467218 189922 497758 189978
rect 497814 189922 497882 189978
rect 497938 189922 528478 189978
rect 528534 189922 528602 189978
rect 528658 189922 559198 189978
rect 559254 189922 559322 189978
rect 559378 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 44518 184350
rect 44574 184294 44642 184350
rect 44698 184294 75238 184350
rect 75294 184294 75362 184350
rect 75418 184294 105958 184350
rect 106014 184294 106082 184350
rect 106138 184294 136678 184350
rect 136734 184294 136802 184350
rect 136858 184294 167398 184350
rect 167454 184294 167522 184350
rect 167578 184294 198118 184350
rect 198174 184294 198242 184350
rect 198298 184294 228838 184350
rect 228894 184294 228962 184350
rect 229018 184294 259558 184350
rect 259614 184294 259682 184350
rect 259738 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 305538 184350
rect 305594 184294 305662 184350
rect 305718 184294 314106 184350
rect 314162 184294 314230 184350
rect 314286 184294 322674 184350
rect 322730 184294 322798 184350
rect 322854 184294 331242 184350
rect 331298 184294 331366 184350
rect 331422 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 359518 184350
rect 359574 184294 359642 184350
rect 359698 184294 390238 184350
rect 390294 184294 390362 184350
rect 390418 184294 420958 184350
rect 421014 184294 421082 184350
rect 421138 184294 451678 184350
rect 451734 184294 451802 184350
rect 451858 184294 482398 184350
rect 482454 184294 482522 184350
rect 482578 184294 513118 184350
rect 513174 184294 513242 184350
rect 513298 184294 543838 184350
rect 543894 184294 543962 184350
rect 544018 184294 574558 184350
rect 574614 184294 574682 184350
rect 574738 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 44518 184226
rect 44574 184170 44642 184226
rect 44698 184170 75238 184226
rect 75294 184170 75362 184226
rect 75418 184170 105958 184226
rect 106014 184170 106082 184226
rect 106138 184170 136678 184226
rect 136734 184170 136802 184226
rect 136858 184170 167398 184226
rect 167454 184170 167522 184226
rect 167578 184170 198118 184226
rect 198174 184170 198242 184226
rect 198298 184170 228838 184226
rect 228894 184170 228962 184226
rect 229018 184170 259558 184226
rect 259614 184170 259682 184226
rect 259738 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 305538 184226
rect 305594 184170 305662 184226
rect 305718 184170 314106 184226
rect 314162 184170 314230 184226
rect 314286 184170 322674 184226
rect 322730 184170 322798 184226
rect 322854 184170 331242 184226
rect 331298 184170 331366 184226
rect 331422 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 359518 184226
rect 359574 184170 359642 184226
rect 359698 184170 390238 184226
rect 390294 184170 390362 184226
rect 390418 184170 420958 184226
rect 421014 184170 421082 184226
rect 421138 184170 451678 184226
rect 451734 184170 451802 184226
rect 451858 184170 482398 184226
rect 482454 184170 482522 184226
rect 482578 184170 513118 184226
rect 513174 184170 513242 184226
rect 513298 184170 543838 184226
rect 543894 184170 543962 184226
rect 544018 184170 574558 184226
rect 574614 184170 574682 184226
rect 574738 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 44518 184102
rect 44574 184046 44642 184102
rect 44698 184046 75238 184102
rect 75294 184046 75362 184102
rect 75418 184046 105958 184102
rect 106014 184046 106082 184102
rect 106138 184046 136678 184102
rect 136734 184046 136802 184102
rect 136858 184046 167398 184102
rect 167454 184046 167522 184102
rect 167578 184046 198118 184102
rect 198174 184046 198242 184102
rect 198298 184046 228838 184102
rect 228894 184046 228962 184102
rect 229018 184046 259558 184102
rect 259614 184046 259682 184102
rect 259738 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 305538 184102
rect 305594 184046 305662 184102
rect 305718 184046 314106 184102
rect 314162 184046 314230 184102
rect 314286 184046 322674 184102
rect 322730 184046 322798 184102
rect 322854 184046 331242 184102
rect 331298 184046 331366 184102
rect 331422 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 359518 184102
rect 359574 184046 359642 184102
rect 359698 184046 390238 184102
rect 390294 184046 390362 184102
rect 390418 184046 420958 184102
rect 421014 184046 421082 184102
rect 421138 184046 451678 184102
rect 451734 184046 451802 184102
rect 451858 184046 482398 184102
rect 482454 184046 482522 184102
rect 482578 184046 513118 184102
rect 513174 184046 513242 184102
rect 513298 184046 543838 184102
rect 543894 184046 543962 184102
rect 544018 184046 574558 184102
rect 574614 184046 574682 184102
rect 574738 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 44518 183978
rect 44574 183922 44642 183978
rect 44698 183922 75238 183978
rect 75294 183922 75362 183978
rect 75418 183922 105958 183978
rect 106014 183922 106082 183978
rect 106138 183922 136678 183978
rect 136734 183922 136802 183978
rect 136858 183922 167398 183978
rect 167454 183922 167522 183978
rect 167578 183922 198118 183978
rect 198174 183922 198242 183978
rect 198298 183922 228838 183978
rect 228894 183922 228962 183978
rect 229018 183922 259558 183978
rect 259614 183922 259682 183978
rect 259738 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 305538 183978
rect 305594 183922 305662 183978
rect 305718 183922 314106 183978
rect 314162 183922 314230 183978
rect 314286 183922 322674 183978
rect 322730 183922 322798 183978
rect 322854 183922 331242 183978
rect 331298 183922 331366 183978
rect 331422 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 359518 183978
rect 359574 183922 359642 183978
rect 359698 183922 390238 183978
rect 390294 183922 390362 183978
rect 390418 183922 420958 183978
rect 421014 183922 421082 183978
rect 421138 183922 451678 183978
rect 451734 183922 451802 183978
rect 451858 183922 482398 183978
rect 482454 183922 482522 183978
rect 482578 183922 513118 183978
rect 513174 183922 513242 183978
rect 513298 183922 543838 183978
rect 543894 183922 543962 183978
rect 544018 183922 574558 183978
rect 574614 183922 574682 183978
rect 574738 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 59878 172350
rect 59934 172294 60002 172350
rect 60058 172294 90598 172350
rect 90654 172294 90722 172350
rect 90778 172294 121318 172350
rect 121374 172294 121442 172350
rect 121498 172294 152038 172350
rect 152094 172294 152162 172350
rect 152218 172294 182758 172350
rect 182814 172294 182882 172350
rect 182938 172294 213478 172350
rect 213534 172294 213602 172350
rect 213658 172294 244198 172350
rect 244254 172294 244322 172350
rect 244378 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 309822 172350
rect 309878 172294 309946 172350
rect 310002 172294 318390 172350
rect 318446 172294 318514 172350
rect 318570 172294 326958 172350
rect 327014 172294 327082 172350
rect 327138 172294 335526 172350
rect 335582 172294 335650 172350
rect 335706 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 374878 172350
rect 374934 172294 375002 172350
rect 375058 172294 405598 172350
rect 405654 172294 405722 172350
rect 405778 172294 436318 172350
rect 436374 172294 436442 172350
rect 436498 172294 467038 172350
rect 467094 172294 467162 172350
rect 467218 172294 497758 172350
rect 497814 172294 497882 172350
rect 497938 172294 528478 172350
rect 528534 172294 528602 172350
rect 528658 172294 559198 172350
rect 559254 172294 559322 172350
rect 559378 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 59878 172226
rect 59934 172170 60002 172226
rect 60058 172170 90598 172226
rect 90654 172170 90722 172226
rect 90778 172170 121318 172226
rect 121374 172170 121442 172226
rect 121498 172170 152038 172226
rect 152094 172170 152162 172226
rect 152218 172170 182758 172226
rect 182814 172170 182882 172226
rect 182938 172170 213478 172226
rect 213534 172170 213602 172226
rect 213658 172170 244198 172226
rect 244254 172170 244322 172226
rect 244378 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 309822 172226
rect 309878 172170 309946 172226
rect 310002 172170 318390 172226
rect 318446 172170 318514 172226
rect 318570 172170 326958 172226
rect 327014 172170 327082 172226
rect 327138 172170 335526 172226
rect 335582 172170 335650 172226
rect 335706 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 374878 172226
rect 374934 172170 375002 172226
rect 375058 172170 405598 172226
rect 405654 172170 405722 172226
rect 405778 172170 436318 172226
rect 436374 172170 436442 172226
rect 436498 172170 467038 172226
rect 467094 172170 467162 172226
rect 467218 172170 497758 172226
rect 497814 172170 497882 172226
rect 497938 172170 528478 172226
rect 528534 172170 528602 172226
rect 528658 172170 559198 172226
rect 559254 172170 559322 172226
rect 559378 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 59878 172102
rect 59934 172046 60002 172102
rect 60058 172046 90598 172102
rect 90654 172046 90722 172102
rect 90778 172046 121318 172102
rect 121374 172046 121442 172102
rect 121498 172046 152038 172102
rect 152094 172046 152162 172102
rect 152218 172046 182758 172102
rect 182814 172046 182882 172102
rect 182938 172046 213478 172102
rect 213534 172046 213602 172102
rect 213658 172046 244198 172102
rect 244254 172046 244322 172102
rect 244378 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 309822 172102
rect 309878 172046 309946 172102
rect 310002 172046 318390 172102
rect 318446 172046 318514 172102
rect 318570 172046 326958 172102
rect 327014 172046 327082 172102
rect 327138 172046 335526 172102
rect 335582 172046 335650 172102
rect 335706 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 374878 172102
rect 374934 172046 375002 172102
rect 375058 172046 405598 172102
rect 405654 172046 405722 172102
rect 405778 172046 436318 172102
rect 436374 172046 436442 172102
rect 436498 172046 467038 172102
rect 467094 172046 467162 172102
rect 467218 172046 497758 172102
rect 497814 172046 497882 172102
rect 497938 172046 528478 172102
rect 528534 172046 528602 172102
rect 528658 172046 559198 172102
rect 559254 172046 559322 172102
rect 559378 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 59878 171978
rect 59934 171922 60002 171978
rect 60058 171922 90598 171978
rect 90654 171922 90722 171978
rect 90778 171922 121318 171978
rect 121374 171922 121442 171978
rect 121498 171922 152038 171978
rect 152094 171922 152162 171978
rect 152218 171922 182758 171978
rect 182814 171922 182882 171978
rect 182938 171922 213478 171978
rect 213534 171922 213602 171978
rect 213658 171922 244198 171978
rect 244254 171922 244322 171978
rect 244378 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 309822 171978
rect 309878 171922 309946 171978
rect 310002 171922 318390 171978
rect 318446 171922 318514 171978
rect 318570 171922 326958 171978
rect 327014 171922 327082 171978
rect 327138 171922 335526 171978
rect 335582 171922 335650 171978
rect 335706 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 374878 171978
rect 374934 171922 375002 171978
rect 375058 171922 405598 171978
rect 405654 171922 405722 171978
rect 405778 171922 436318 171978
rect 436374 171922 436442 171978
rect 436498 171922 467038 171978
rect 467094 171922 467162 171978
rect 467218 171922 497758 171978
rect 497814 171922 497882 171978
rect 497938 171922 528478 171978
rect 528534 171922 528602 171978
rect 528658 171922 559198 171978
rect 559254 171922 559322 171978
rect 559378 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect 351804 167338 356596 167354
rect 351804 167282 351820 167338
rect 351876 167282 356524 167338
rect 356580 167282 356596 167338
rect 351804 167266 356596 167282
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 44518 166350
rect 44574 166294 44642 166350
rect 44698 166294 75238 166350
rect 75294 166294 75362 166350
rect 75418 166294 105958 166350
rect 106014 166294 106082 166350
rect 106138 166294 136678 166350
rect 136734 166294 136802 166350
rect 136858 166294 167398 166350
rect 167454 166294 167522 166350
rect 167578 166294 198118 166350
rect 198174 166294 198242 166350
rect 198298 166294 228838 166350
rect 228894 166294 228962 166350
rect 229018 166294 259558 166350
rect 259614 166294 259682 166350
rect 259738 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 305538 166350
rect 305594 166294 305662 166350
rect 305718 166294 314106 166350
rect 314162 166294 314230 166350
rect 314286 166294 322674 166350
rect 322730 166294 322798 166350
rect 322854 166294 331242 166350
rect 331298 166294 331366 166350
rect 331422 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 44518 166226
rect 44574 166170 44642 166226
rect 44698 166170 75238 166226
rect 75294 166170 75362 166226
rect 75418 166170 105958 166226
rect 106014 166170 106082 166226
rect 106138 166170 136678 166226
rect 136734 166170 136802 166226
rect 136858 166170 167398 166226
rect 167454 166170 167522 166226
rect 167578 166170 198118 166226
rect 198174 166170 198242 166226
rect 198298 166170 228838 166226
rect 228894 166170 228962 166226
rect 229018 166170 259558 166226
rect 259614 166170 259682 166226
rect 259738 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 305538 166226
rect 305594 166170 305662 166226
rect 305718 166170 314106 166226
rect 314162 166170 314230 166226
rect 314286 166170 322674 166226
rect 322730 166170 322798 166226
rect 322854 166170 331242 166226
rect 331298 166170 331366 166226
rect 331422 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 44518 166102
rect 44574 166046 44642 166102
rect 44698 166046 75238 166102
rect 75294 166046 75362 166102
rect 75418 166046 105958 166102
rect 106014 166046 106082 166102
rect 106138 166046 136678 166102
rect 136734 166046 136802 166102
rect 136858 166046 167398 166102
rect 167454 166046 167522 166102
rect 167578 166046 198118 166102
rect 198174 166046 198242 166102
rect 198298 166046 228838 166102
rect 228894 166046 228962 166102
rect 229018 166046 259558 166102
rect 259614 166046 259682 166102
rect 259738 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 305538 166102
rect 305594 166046 305662 166102
rect 305718 166046 314106 166102
rect 314162 166046 314230 166102
rect 314286 166046 322674 166102
rect 322730 166046 322798 166102
rect 322854 166046 331242 166102
rect 331298 166046 331366 166102
rect 331422 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 44518 165978
rect 44574 165922 44642 165978
rect 44698 165922 75238 165978
rect 75294 165922 75362 165978
rect 75418 165922 105958 165978
rect 106014 165922 106082 165978
rect 106138 165922 136678 165978
rect 136734 165922 136802 165978
rect 136858 165922 167398 165978
rect 167454 165922 167522 165978
rect 167578 165922 198118 165978
rect 198174 165922 198242 165978
rect 198298 165922 228838 165978
rect 228894 165922 228962 165978
rect 229018 165922 259558 165978
rect 259614 165922 259682 165978
rect 259738 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 305538 165978
rect 305594 165922 305662 165978
rect 305718 165922 314106 165978
rect 314162 165922 314230 165978
rect 314286 165922 322674 165978
rect 322730 165922 322798 165978
rect 322854 165922 331242 165978
rect 331298 165922 331366 165978
rect 331422 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect 354268 165538 488980 165554
rect 354268 165482 354284 165538
rect 354340 165482 488908 165538
rect 488964 165482 488980 165538
rect 354268 165466 488980 165482
rect 356060 164818 489316 164834
rect 356060 164762 356076 164818
rect 356132 164762 489244 164818
rect 489300 164762 489316 164818
rect 356060 164746 489316 164762
rect 337020 164638 590564 164654
rect 337020 164582 337036 164638
rect 337092 164582 590492 164638
rect 590548 164582 590564 164638
rect 337020 164566 590564 164582
rect 354940 164098 487860 164114
rect 354940 164042 354956 164098
rect 355012 164042 487788 164098
rect 487844 164042 487860 164098
rect 354940 164026 487860 164042
rect 355052 163918 493236 163934
rect 355052 163862 355068 163918
rect 355124 163862 493164 163918
rect 493220 163862 493236 163918
rect 355052 163846 493236 163862
rect 350796 163738 554388 163754
rect 350796 163682 350812 163738
rect 350868 163682 554316 163738
rect 554372 163682 554388 163738
rect 350796 163666 554388 163682
rect 346876 162838 539380 162854
rect 346876 162782 346892 162838
rect 346948 162782 539308 162838
rect 539364 162782 539380 162838
rect 346876 162766 539380 162782
rect 353484 162478 483828 162494
rect 353484 162422 353500 162478
rect 353556 162422 483756 162478
rect 483812 162422 483828 162478
rect 353484 162406 483828 162422
rect 354380 162298 491892 162314
rect 354380 162242 354396 162298
rect 354452 162242 491820 162298
rect 491876 162242 491892 162298
rect 354380 162226 491892 162242
rect 348444 162118 559204 162134
rect 348444 162062 348460 162118
rect 348516 162062 559132 162118
rect 559188 162062 559204 162118
rect 348444 162046 559204 162062
rect 340604 161218 546548 161234
rect 340604 161162 340620 161218
rect 340676 161162 546476 161218
rect 546532 161162 546548 161218
rect 340604 161146 546548 161162
rect 346316 160858 480468 160874
rect 346316 160802 346332 160858
rect 346388 160802 480396 160858
rect 480452 160802 480468 160858
rect 346316 160786 480468 160802
rect 342060 160678 554836 160694
rect 342060 160622 342076 160678
rect 342132 160622 554764 160678
rect 554820 160622 554836 160678
rect 342060 160606 554836 160622
rect 340268 160498 555284 160514
rect 340268 160442 340284 160498
rect 340340 160442 555212 160498
rect 555268 160442 555284 160498
rect 340268 160426 555284 160442
rect 355276 159598 532436 159614
rect 355276 159542 355292 159598
rect 355348 159542 532364 159598
rect 532420 159542 532436 159598
rect 355276 159526 532436 159542
rect 354156 158878 554612 158894
rect 354156 158822 354172 158878
rect 354228 158822 554540 158878
rect 554596 158822 554612 158878
rect 354156 158806 554612 158822
rect 344188 158698 556404 158714
rect 344188 158642 344204 158698
rect 344260 158642 556332 158698
rect 556388 158642 556404 158698
rect 344188 158626 556404 158642
rect 346876 157978 553940 157994
rect 346876 157922 346892 157978
rect 346948 157922 553868 157978
rect 553924 157922 553940 157978
rect 346876 157906 553940 157922
rect 339484 157798 497940 157814
rect 339484 157742 339500 157798
rect 339556 157742 497868 157798
rect 497924 157742 497940 157798
rect 339484 157726 497940 157742
rect 353596 157618 477108 157634
rect 353596 157562 353612 157618
rect 353668 157562 477036 157618
rect 477092 157562 477108 157618
rect 353596 157546 477108 157562
rect 298940 157438 306644 157454
rect 298940 157382 298956 157438
rect 299012 157382 306572 157438
rect 306628 157382 306644 157438
rect 298940 157366 306644 157382
rect 346092 157438 460308 157454
rect 346092 157382 346108 157438
rect 346164 157382 460236 157438
rect 460292 157382 460308 157438
rect 346092 157366 460308 157382
rect 461228 156538 494580 156554
rect 461228 156482 461244 156538
rect 461300 156482 494508 156538
rect 494564 156482 494580 156538
rect 461228 156466 494580 156482
rect 421580 156358 554500 156374
rect 421580 156302 421596 156358
rect 421652 156302 554428 156358
rect 554484 156302 554500 156358
rect 421580 156286 554500 156302
rect 341948 156178 460196 156194
rect 341948 156122 341964 156178
rect 342020 156122 460124 156178
rect 460180 156122 460196 156178
rect 341948 156106 460196 156122
rect 355164 155638 485172 155654
rect 355164 155582 355180 155638
rect 355236 155582 485100 155638
rect 485156 155582 485172 155638
rect 355164 155566 485172 155582
rect 345308 155458 557860 155474
rect 345308 155402 345324 155458
rect 345380 155402 557788 155458
rect 557844 155402 557860 155458
rect 345308 155386 557860 155402
rect 460332 154918 475764 154934
rect 460332 154862 460348 154918
rect 460404 154862 475692 154918
rect 475748 154862 475764 154918
rect 460332 154846 475764 154862
rect 458428 154738 555172 154754
rect 458428 154682 458444 154738
rect 458500 154682 555100 154738
rect 555156 154682 555172 154738
rect 458428 154666 555172 154682
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 59878 154350
rect 59934 154294 60002 154350
rect 60058 154294 90598 154350
rect 90654 154294 90722 154350
rect 90778 154294 121318 154350
rect 121374 154294 121442 154350
rect 121498 154294 152038 154350
rect 152094 154294 152162 154350
rect 152218 154294 182758 154350
rect 182814 154294 182882 154350
rect 182938 154294 213478 154350
rect 213534 154294 213602 154350
rect 213658 154294 244198 154350
rect 244254 154294 244322 154350
rect 244378 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 59878 154226
rect 59934 154170 60002 154226
rect 60058 154170 90598 154226
rect 90654 154170 90722 154226
rect 90778 154170 121318 154226
rect 121374 154170 121442 154226
rect 121498 154170 152038 154226
rect 152094 154170 152162 154226
rect 152218 154170 182758 154226
rect 182814 154170 182882 154226
rect 182938 154170 213478 154226
rect 213534 154170 213602 154226
rect 213658 154170 244198 154226
rect 244254 154170 244322 154226
rect 244378 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 59878 154102
rect 59934 154046 60002 154102
rect 60058 154046 90598 154102
rect 90654 154046 90722 154102
rect 90778 154046 121318 154102
rect 121374 154046 121442 154102
rect 121498 154046 152038 154102
rect 152094 154046 152162 154102
rect 152218 154046 182758 154102
rect 182814 154046 182882 154102
rect 182938 154046 213478 154102
rect 213534 154046 213602 154102
rect 213658 154046 244198 154102
rect 244254 154046 244322 154102
rect 244378 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 59878 153978
rect 59934 153922 60002 153978
rect 60058 153922 90598 153978
rect 90654 153922 90722 153978
rect 90778 153922 121318 153978
rect 121374 153922 121442 153978
rect 121498 153922 152038 153978
rect 152094 153922 152162 153978
rect 152218 153922 182758 153978
rect 182814 153922 182882 153978
rect 182938 153922 213478 153978
rect 213534 153922 213602 153978
rect 213658 153922 244198 153978
rect 244254 153922 244322 153978
rect 244378 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect 272284 153658 499956 153674
rect 272284 153602 272300 153658
rect 272356 153602 499884 153658
rect 499940 153602 499956 153658
rect 272284 153586 499956 153602
rect 274636 153478 498612 153494
rect 274636 153422 274652 153478
rect 274708 153422 498540 153478
rect 498596 153422 498612 153478
rect 274636 153406 498612 153422
rect 497292 152938 556180 152954
rect 497292 152882 497308 152938
rect 497364 152882 556108 152938
rect 556164 152882 556180 152938
rect 497292 152866 556180 152882
rect 296588 152758 590228 152774
rect 296588 152702 296604 152758
rect 296660 152702 590156 152758
rect 590212 152702 590228 152758
rect 296588 152686 590228 152702
rect 348668 152578 463780 152594
rect 348668 152522 348684 152578
rect 348740 152522 463708 152578
rect 463764 152522 463780 152578
rect 348668 152506 463780 152522
rect 350572 152218 558308 152234
rect 350572 152162 350588 152218
rect 350644 152162 558236 152218
rect 558292 152162 558308 152218
rect 350572 152146 558308 152162
rect 350124 152038 558196 152054
rect 350124 151982 350140 152038
rect 350196 151982 558124 152038
rect 558180 151982 558196 152038
rect 350124 151966 558196 151982
rect 457196 151318 590564 151334
rect 457196 151262 457212 151318
rect 457268 151262 590492 151318
rect 590548 151262 590564 151318
rect 457196 151246 590564 151262
rect 350348 150598 555060 150614
rect 350348 150542 350364 150598
rect 350420 150542 554988 150598
rect 555044 150542 555060 150598
rect 350348 150526 555060 150542
rect 346540 150418 557972 150434
rect 346540 150362 346556 150418
rect 346612 150362 557900 150418
rect 557956 150362 557972 150418
rect 346540 150346 557972 150362
rect 456972 150058 553828 150074
rect 456972 150002 456988 150058
rect 457044 150002 553756 150058
rect 553812 150002 553828 150058
rect 456972 149986 553828 150002
rect 461116 149878 477108 149894
rect 461116 149822 461132 149878
rect 461188 149822 477036 149878
rect 477092 149822 477108 149878
rect 461116 149806 477108 149822
rect 342060 149698 554948 149714
rect 342060 149642 342076 149698
rect 342132 149642 554876 149698
rect 554932 149642 554948 149698
rect 342060 149626 554948 149642
rect 346764 148618 557860 148634
rect 346764 148562 346780 148618
rect 346836 148562 557788 148618
rect 557844 148562 557860 148618
rect 346764 148546 557860 148562
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 44518 148350
rect 44574 148294 44642 148350
rect 44698 148294 75238 148350
rect 75294 148294 75362 148350
rect 75418 148294 105958 148350
rect 106014 148294 106082 148350
rect 106138 148294 136678 148350
rect 136734 148294 136802 148350
rect 136858 148294 167398 148350
rect 167454 148294 167522 148350
rect 167578 148294 198118 148350
rect 198174 148294 198242 148350
rect 198298 148294 228838 148350
rect 228894 148294 228962 148350
rect 229018 148294 259558 148350
rect 259614 148294 259682 148350
rect 259738 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 44518 148226
rect 44574 148170 44642 148226
rect 44698 148170 75238 148226
rect 75294 148170 75362 148226
rect 75418 148170 105958 148226
rect 106014 148170 106082 148226
rect 106138 148170 136678 148226
rect 136734 148170 136802 148226
rect 136858 148170 167398 148226
rect 167454 148170 167522 148226
rect 167578 148170 198118 148226
rect 198174 148170 198242 148226
rect 198298 148170 228838 148226
rect 228894 148170 228962 148226
rect 229018 148170 259558 148226
rect 259614 148170 259682 148226
rect 259738 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 44518 148102
rect 44574 148046 44642 148102
rect 44698 148046 75238 148102
rect 75294 148046 75362 148102
rect 75418 148046 105958 148102
rect 106014 148046 106082 148102
rect 106138 148046 136678 148102
rect 136734 148046 136802 148102
rect 136858 148046 167398 148102
rect 167454 148046 167522 148102
rect 167578 148046 198118 148102
rect 198174 148046 198242 148102
rect 198298 148046 228838 148102
rect 228894 148046 228962 148102
rect 229018 148046 259558 148102
rect 259614 148046 259682 148102
rect 259738 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 44518 147978
rect 44574 147922 44642 147978
rect 44698 147922 75238 147978
rect 75294 147922 75362 147978
rect 75418 147922 105958 147978
rect 106014 147922 106082 147978
rect 106138 147922 136678 147978
rect 136734 147922 136802 147978
rect 136858 147922 167398 147978
rect 167454 147922 167522 147978
rect 167578 147922 198118 147978
rect 198174 147922 198242 147978
rect 198298 147922 228838 147978
rect 228894 147922 228962 147978
rect 229018 147922 259558 147978
rect 259614 147922 259682 147978
rect 259738 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect 337636 147718 461316 147734
rect 337636 147662 350028 147718
rect 350084 147662 461244 147718
rect 461300 147662 461316 147718
rect 337636 147646 461316 147662
rect 337636 147014 337724 147646
rect 311596 146998 337724 147014
rect 311596 146942 311612 146998
rect 311668 146942 337724 146998
rect 311596 146926 337724 146942
rect 350796 146098 463668 146114
rect 350796 146042 350812 146098
rect 350868 146042 463596 146098
rect 463652 146042 463668 146098
rect 350796 146026 463668 146042
rect 366252 145918 460532 145934
rect 366252 145862 366268 145918
rect 366324 145862 460460 145918
rect 460516 145862 460532 145918
rect 366252 145846 460532 145862
rect 349340 145738 461764 145754
rect 349340 145682 349356 145738
rect 349412 145682 421708 145738
rect 421764 145682 461692 145738
rect 461748 145682 461764 145738
rect 349340 145666 461764 145682
rect 422476 145558 461652 145574
rect 422476 145502 422492 145558
rect 422548 145502 461580 145558
rect 461636 145502 461652 145558
rect 422476 145486 461652 145502
rect 352588 144478 460420 144494
rect 352588 144422 352604 144478
rect 352660 144422 460348 144478
rect 460404 144422 460420 144478
rect 352588 144406 460420 144422
rect 352476 144298 460644 144314
rect 352476 144242 352492 144298
rect 352548 144242 460572 144298
rect 460628 144242 460644 144298
rect 352476 144226 460644 144242
rect 351916 143938 352676 143954
rect 351916 143882 351932 143938
rect 351988 143882 352604 143938
rect 352660 143882 352676 143938
rect 351916 143866 352676 143882
rect 337636 142678 462996 142694
rect 337636 142622 352716 142678
rect 352772 142622 462924 142678
rect 462980 142622 462996 142678
rect 337636 142606 462996 142622
rect 337636 141974 337724 142606
rect 293228 141958 337724 141974
rect 293228 141902 293244 141958
rect 293300 141902 337724 141958
rect 293228 141886 337724 141902
rect 351020 141058 462884 141074
rect 351020 141002 351036 141058
rect 351092 141002 462812 141058
rect 462868 141002 462884 141058
rect 351020 140986 462884 141002
rect 352028 140878 461204 140894
rect 352028 140822 352044 140878
rect 352100 140822 461132 140878
rect 461188 140822 461204 140878
rect 352028 140806 461204 140822
rect 339148 139438 463108 139454
rect 339148 139382 339164 139438
rect 339220 139382 463036 139438
rect 463092 139382 463108 139438
rect 339148 139366 463108 139382
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 59878 136350
rect 59934 136294 60002 136350
rect 60058 136294 90598 136350
rect 90654 136294 90722 136350
rect 90778 136294 121318 136350
rect 121374 136294 121442 136350
rect 121498 136294 152038 136350
rect 152094 136294 152162 136350
rect 152218 136294 182758 136350
rect 182814 136294 182882 136350
rect 182938 136294 213478 136350
rect 213534 136294 213602 136350
rect 213658 136294 244198 136350
rect 244254 136294 244322 136350
rect 244378 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 479878 136350
rect 479934 136294 480002 136350
rect 480058 136294 510598 136350
rect 510654 136294 510722 136350
rect 510778 136294 541318 136350
rect 541374 136294 541442 136350
rect 541498 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 59878 136226
rect 59934 136170 60002 136226
rect 60058 136170 90598 136226
rect 90654 136170 90722 136226
rect 90778 136170 121318 136226
rect 121374 136170 121442 136226
rect 121498 136170 152038 136226
rect 152094 136170 152162 136226
rect 152218 136170 182758 136226
rect 182814 136170 182882 136226
rect 182938 136170 213478 136226
rect 213534 136170 213602 136226
rect 213658 136170 244198 136226
rect 244254 136170 244322 136226
rect 244378 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 479878 136226
rect 479934 136170 480002 136226
rect 480058 136170 510598 136226
rect 510654 136170 510722 136226
rect 510778 136170 541318 136226
rect 541374 136170 541442 136226
rect 541498 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 59878 136102
rect 59934 136046 60002 136102
rect 60058 136046 90598 136102
rect 90654 136046 90722 136102
rect 90778 136046 121318 136102
rect 121374 136046 121442 136102
rect 121498 136046 152038 136102
rect 152094 136046 152162 136102
rect 152218 136046 182758 136102
rect 182814 136046 182882 136102
rect 182938 136046 213478 136102
rect 213534 136046 213602 136102
rect 213658 136046 244198 136102
rect 244254 136046 244322 136102
rect 244378 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 479878 136102
rect 479934 136046 480002 136102
rect 480058 136046 510598 136102
rect 510654 136046 510722 136102
rect 510778 136046 541318 136102
rect 541374 136046 541442 136102
rect 541498 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 59878 135978
rect 59934 135922 60002 135978
rect 60058 135922 90598 135978
rect 90654 135922 90722 135978
rect 90778 135922 121318 135978
rect 121374 135922 121442 135978
rect 121498 135922 152038 135978
rect 152094 135922 152162 135978
rect 152218 135922 182758 135978
rect 182814 135922 182882 135978
rect 182938 135922 213478 135978
rect 213534 135922 213602 135978
rect 213658 135922 244198 135978
rect 244254 135922 244322 135978
rect 244378 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 479878 135978
rect 479934 135922 480002 135978
rect 480058 135922 510598 135978
rect 510654 135922 510722 135978
rect 510778 135922 541318 135978
rect 541374 135922 541442 135978
rect 541498 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 44518 130350
rect 44574 130294 44642 130350
rect 44698 130294 75238 130350
rect 75294 130294 75362 130350
rect 75418 130294 105958 130350
rect 106014 130294 106082 130350
rect 106138 130294 136678 130350
rect 136734 130294 136802 130350
rect 136858 130294 167398 130350
rect 167454 130294 167522 130350
rect 167578 130294 198118 130350
rect 198174 130294 198242 130350
rect 198298 130294 228838 130350
rect 228894 130294 228962 130350
rect 229018 130294 259558 130350
rect 259614 130294 259682 130350
rect 259738 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 464518 130350
rect 464574 130294 464642 130350
rect 464698 130294 495238 130350
rect 495294 130294 495362 130350
rect 495418 130294 525958 130350
rect 526014 130294 526082 130350
rect 526138 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 44518 130226
rect 44574 130170 44642 130226
rect 44698 130170 75238 130226
rect 75294 130170 75362 130226
rect 75418 130170 105958 130226
rect 106014 130170 106082 130226
rect 106138 130170 136678 130226
rect 136734 130170 136802 130226
rect 136858 130170 167398 130226
rect 167454 130170 167522 130226
rect 167578 130170 198118 130226
rect 198174 130170 198242 130226
rect 198298 130170 228838 130226
rect 228894 130170 228962 130226
rect 229018 130170 259558 130226
rect 259614 130170 259682 130226
rect 259738 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 464518 130226
rect 464574 130170 464642 130226
rect 464698 130170 495238 130226
rect 495294 130170 495362 130226
rect 495418 130170 525958 130226
rect 526014 130170 526082 130226
rect 526138 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 44518 130102
rect 44574 130046 44642 130102
rect 44698 130046 75238 130102
rect 75294 130046 75362 130102
rect 75418 130046 105958 130102
rect 106014 130046 106082 130102
rect 106138 130046 136678 130102
rect 136734 130046 136802 130102
rect 136858 130046 167398 130102
rect 167454 130046 167522 130102
rect 167578 130046 198118 130102
rect 198174 130046 198242 130102
rect 198298 130046 228838 130102
rect 228894 130046 228962 130102
rect 229018 130046 259558 130102
rect 259614 130046 259682 130102
rect 259738 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 464518 130102
rect 464574 130046 464642 130102
rect 464698 130046 495238 130102
rect 495294 130046 495362 130102
rect 495418 130046 525958 130102
rect 526014 130046 526082 130102
rect 526138 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 44518 129978
rect 44574 129922 44642 129978
rect 44698 129922 75238 129978
rect 75294 129922 75362 129978
rect 75418 129922 105958 129978
rect 106014 129922 106082 129978
rect 106138 129922 136678 129978
rect 136734 129922 136802 129978
rect 136858 129922 167398 129978
rect 167454 129922 167522 129978
rect 167578 129922 198118 129978
rect 198174 129922 198242 129978
rect 198298 129922 228838 129978
rect 228894 129922 228962 129978
rect 229018 129922 259558 129978
rect 259614 129922 259682 129978
rect 259738 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 464518 129978
rect 464574 129922 464642 129978
rect 464698 129922 495238 129978
rect 495294 129922 495362 129978
rect 495418 129922 525958 129978
rect 526014 129922 526082 129978
rect 526138 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect 423260 122518 460756 122534
rect 423260 122462 423276 122518
rect 423332 122462 460684 122518
rect 460740 122462 460756 122518
rect 423260 122446 460756 122462
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 59878 118350
rect 59934 118294 60002 118350
rect 60058 118294 90598 118350
rect 90654 118294 90722 118350
rect 90778 118294 121318 118350
rect 121374 118294 121442 118350
rect 121498 118294 152038 118350
rect 152094 118294 152162 118350
rect 152218 118294 182758 118350
rect 182814 118294 182882 118350
rect 182938 118294 213478 118350
rect 213534 118294 213602 118350
rect 213658 118294 244198 118350
rect 244254 118294 244322 118350
rect 244378 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 479878 118350
rect 479934 118294 480002 118350
rect 480058 118294 510598 118350
rect 510654 118294 510722 118350
rect 510778 118294 541318 118350
rect 541374 118294 541442 118350
rect 541498 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 59878 118226
rect 59934 118170 60002 118226
rect 60058 118170 90598 118226
rect 90654 118170 90722 118226
rect 90778 118170 121318 118226
rect 121374 118170 121442 118226
rect 121498 118170 152038 118226
rect 152094 118170 152162 118226
rect 152218 118170 182758 118226
rect 182814 118170 182882 118226
rect 182938 118170 213478 118226
rect 213534 118170 213602 118226
rect 213658 118170 244198 118226
rect 244254 118170 244322 118226
rect 244378 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 479878 118226
rect 479934 118170 480002 118226
rect 480058 118170 510598 118226
rect 510654 118170 510722 118226
rect 510778 118170 541318 118226
rect 541374 118170 541442 118226
rect 541498 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 59878 118102
rect 59934 118046 60002 118102
rect 60058 118046 90598 118102
rect 90654 118046 90722 118102
rect 90778 118046 121318 118102
rect 121374 118046 121442 118102
rect 121498 118046 152038 118102
rect 152094 118046 152162 118102
rect 152218 118046 182758 118102
rect 182814 118046 182882 118102
rect 182938 118046 213478 118102
rect 213534 118046 213602 118102
rect 213658 118046 244198 118102
rect 244254 118046 244322 118102
rect 244378 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 479878 118102
rect 479934 118046 480002 118102
rect 480058 118046 510598 118102
rect 510654 118046 510722 118102
rect 510778 118046 541318 118102
rect 541374 118046 541442 118102
rect 541498 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 59878 117978
rect 59934 117922 60002 117978
rect 60058 117922 90598 117978
rect 90654 117922 90722 117978
rect 90778 117922 121318 117978
rect 121374 117922 121442 117978
rect 121498 117922 152038 117978
rect 152094 117922 152162 117978
rect 152218 117922 182758 117978
rect 182814 117922 182882 117978
rect 182938 117922 213478 117978
rect 213534 117922 213602 117978
rect 213658 117922 244198 117978
rect 244254 117922 244322 117978
rect 244378 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 479878 117978
rect 479934 117922 480002 117978
rect 480058 117922 510598 117978
rect 510654 117922 510722 117978
rect 510778 117922 541318 117978
rect 541374 117922 541442 117978
rect 541498 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect 553628 116938 555284 116954
rect 553628 116882 553644 116938
rect 553700 116882 555212 116938
rect 555268 116882 555284 116938
rect 553628 116866 555284 116882
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 44518 112350
rect 44574 112294 44642 112350
rect 44698 112294 75238 112350
rect 75294 112294 75362 112350
rect 75418 112294 105958 112350
rect 106014 112294 106082 112350
rect 106138 112294 136678 112350
rect 136734 112294 136802 112350
rect 136858 112294 167398 112350
rect 167454 112294 167522 112350
rect 167578 112294 198118 112350
rect 198174 112294 198242 112350
rect 198298 112294 228838 112350
rect 228894 112294 228962 112350
rect 229018 112294 259558 112350
rect 259614 112294 259682 112350
rect 259738 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 464518 112350
rect 464574 112294 464642 112350
rect 464698 112294 495238 112350
rect 495294 112294 495362 112350
rect 495418 112294 525958 112350
rect 526014 112294 526082 112350
rect 526138 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 44518 112226
rect 44574 112170 44642 112226
rect 44698 112170 75238 112226
rect 75294 112170 75362 112226
rect 75418 112170 105958 112226
rect 106014 112170 106082 112226
rect 106138 112170 136678 112226
rect 136734 112170 136802 112226
rect 136858 112170 167398 112226
rect 167454 112170 167522 112226
rect 167578 112170 198118 112226
rect 198174 112170 198242 112226
rect 198298 112170 228838 112226
rect 228894 112170 228962 112226
rect 229018 112170 259558 112226
rect 259614 112170 259682 112226
rect 259738 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 464518 112226
rect 464574 112170 464642 112226
rect 464698 112170 495238 112226
rect 495294 112170 495362 112226
rect 495418 112170 525958 112226
rect 526014 112170 526082 112226
rect 526138 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 44518 112102
rect 44574 112046 44642 112102
rect 44698 112046 75238 112102
rect 75294 112046 75362 112102
rect 75418 112046 105958 112102
rect 106014 112046 106082 112102
rect 106138 112046 136678 112102
rect 136734 112046 136802 112102
rect 136858 112046 167398 112102
rect 167454 112046 167522 112102
rect 167578 112046 198118 112102
rect 198174 112046 198242 112102
rect 198298 112046 228838 112102
rect 228894 112046 228962 112102
rect 229018 112046 259558 112102
rect 259614 112046 259682 112102
rect 259738 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 464518 112102
rect 464574 112046 464642 112102
rect 464698 112046 495238 112102
rect 495294 112046 495362 112102
rect 495418 112046 525958 112102
rect 526014 112046 526082 112102
rect 526138 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 44518 111978
rect 44574 111922 44642 111978
rect 44698 111922 75238 111978
rect 75294 111922 75362 111978
rect 75418 111922 105958 111978
rect 106014 111922 106082 111978
rect 106138 111922 136678 111978
rect 136734 111922 136802 111978
rect 136858 111922 167398 111978
rect 167454 111922 167522 111978
rect 167578 111922 198118 111978
rect 198174 111922 198242 111978
rect 198298 111922 228838 111978
rect 228894 111922 228962 111978
rect 229018 111922 259558 111978
rect 259614 111922 259682 111978
rect 259738 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 464518 111978
rect 464574 111922 464642 111978
rect 464698 111922 495238 111978
rect 495294 111922 495362 111978
rect 495418 111922 525958 111978
rect 526014 111922 526082 111978
rect 526138 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect 268588 110098 398260 110114
rect 268588 110042 268604 110098
rect 268660 110042 398188 110098
rect 398244 110042 398260 110098
rect 268588 110026 398260 110042
rect 268700 106678 396580 106694
rect 268700 106622 268716 106678
rect 268772 106622 396508 106678
rect 396564 106622 396580 106678
rect 268700 106606 396580 106622
rect 553292 105418 554164 105434
rect 553292 105362 553308 105418
rect 553364 105362 554092 105418
rect 554148 105362 554164 105418
rect 553292 105346 554164 105362
rect 293116 104158 392436 104174
rect 293116 104102 293132 104158
rect 293188 104102 392364 104158
rect 392420 104102 392436 104158
rect 293116 104086 392436 104102
rect 296476 103978 389300 103994
rect 296476 103922 296492 103978
rect 296548 103922 389228 103978
rect 389284 103922 389300 103978
rect 296476 103906 389300 103922
rect 553740 103978 554388 103994
rect 553740 103922 553756 103978
rect 553812 103922 554316 103978
rect 554372 103922 554388 103978
rect 553740 103906 554388 103922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 59878 100350
rect 59934 100294 60002 100350
rect 60058 100294 90598 100350
rect 90654 100294 90722 100350
rect 90778 100294 121318 100350
rect 121374 100294 121442 100350
rect 121498 100294 152038 100350
rect 152094 100294 152162 100350
rect 152218 100294 182758 100350
rect 182814 100294 182882 100350
rect 182938 100294 213478 100350
rect 213534 100294 213602 100350
rect 213658 100294 244198 100350
rect 244254 100294 244322 100350
rect 244378 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 479878 100350
rect 479934 100294 480002 100350
rect 480058 100294 510598 100350
rect 510654 100294 510722 100350
rect 510778 100294 541318 100350
rect 541374 100294 541442 100350
rect 541498 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 59878 100226
rect 59934 100170 60002 100226
rect 60058 100170 90598 100226
rect 90654 100170 90722 100226
rect 90778 100170 121318 100226
rect 121374 100170 121442 100226
rect 121498 100170 152038 100226
rect 152094 100170 152162 100226
rect 152218 100170 182758 100226
rect 182814 100170 182882 100226
rect 182938 100170 213478 100226
rect 213534 100170 213602 100226
rect 213658 100170 244198 100226
rect 244254 100170 244322 100226
rect 244378 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 479878 100226
rect 479934 100170 480002 100226
rect 480058 100170 510598 100226
rect 510654 100170 510722 100226
rect 510778 100170 541318 100226
rect 541374 100170 541442 100226
rect 541498 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 59878 100102
rect 59934 100046 60002 100102
rect 60058 100046 90598 100102
rect 90654 100046 90722 100102
rect 90778 100046 121318 100102
rect 121374 100046 121442 100102
rect 121498 100046 152038 100102
rect 152094 100046 152162 100102
rect 152218 100046 182758 100102
rect 182814 100046 182882 100102
rect 182938 100046 213478 100102
rect 213534 100046 213602 100102
rect 213658 100046 244198 100102
rect 244254 100046 244322 100102
rect 244378 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 479878 100102
rect 479934 100046 480002 100102
rect 480058 100046 510598 100102
rect 510654 100046 510722 100102
rect 510778 100046 541318 100102
rect 541374 100046 541442 100102
rect 541498 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 59878 99978
rect 59934 99922 60002 99978
rect 60058 99922 90598 99978
rect 90654 99922 90722 99978
rect 90778 99922 121318 99978
rect 121374 99922 121442 99978
rect 121498 99922 152038 99978
rect 152094 99922 152162 99978
rect 152218 99922 182758 99978
rect 182814 99922 182882 99978
rect 182938 99922 213478 99978
rect 213534 99922 213602 99978
rect 213658 99922 244198 99978
rect 244254 99922 244322 99978
rect 244378 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 479878 99978
rect 479934 99922 480002 99978
rect 480058 99922 510598 99978
rect 510654 99922 510722 99978
rect 510778 99922 541318 99978
rect 541374 99922 541442 99978
rect 541498 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect 553180 99658 554388 99674
rect 553180 99602 553196 99658
rect 553252 99602 554316 99658
rect 554372 99602 554388 99658
rect 553180 99586 554388 99602
rect 353932 98218 457732 98234
rect 353932 98162 353948 98218
rect 354004 98162 457660 98218
rect 457716 98162 457732 98218
rect 353932 98146 457732 98162
rect 342508 94978 457732 94994
rect 342508 94922 342524 94978
rect 342580 94922 457660 94978
rect 457716 94922 457732 94978
rect 342508 94906 457732 94922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 44518 94350
rect 44574 94294 44642 94350
rect 44698 94294 75238 94350
rect 75294 94294 75362 94350
rect 75418 94294 105958 94350
rect 106014 94294 106082 94350
rect 106138 94294 136678 94350
rect 136734 94294 136802 94350
rect 136858 94294 167398 94350
rect 167454 94294 167522 94350
rect 167578 94294 198118 94350
rect 198174 94294 198242 94350
rect 198298 94294 228838 94350
rect 228894 94294 228962 94350
rect 229018 94294 259558 94350
rect 259614 94294 259682 94350
rect 259738 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 374518 94350
rect 374574 94294 374642 94350
rect 374698 94294 405238 94350
rect 405294 94294 405362 94350
rect 405418 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 464518 94350
rect 464574 94294 464642 94350
rect 464698 94294 495238 94350
rect 495294 94294 495362 94350
rect 495418 94294 525958 94350
rect 526014 94294 526082 94350
rect 526138 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 44518 94226
rect 44574 94170 44642 94226
rect 44698 94170 75238 94226
rect 75294 94170 75362 94226
rect 75418 94170 105958 94226
rect 106014 94170 106082 94226
rect 106138 94170 136678 94226
rect 136734 94170 136802 94226
rect 136858 94170 167398 94226
rect 167454 94170 167522 94226
rect 167578 94170 198118 94226
rect 198174 94170 198242 94226
rect 198298 94170 228838 94226
rect 228894 94170 228962 94226
rect 229018 94170 259558 94226
rect 259614 94170 259682 94226
rect 259738 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 374518 94226
rect 374574 94170 374642 94226
rect 374698 94170 405238 94226
rect 405294 94170 405362 94226
rect 405418 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 464518 94226
rect 464574 94170 464642 94226
rect 464698 94170 495238 94226
rect 495294 94170 495362 94226
rect 495418 94170 525958 94226
rect 526014 94170 526082 94226
rect 526138 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 44518 94102
rect 44574 94046 44642 94102
rect 44698 94046 75238 94102
rect 75294 94046 75362 94102
rect 75418 94046 105958 94102
rect 106014 94046 106082 94102
rect 106138 94046 136678 94102
rect 136734 94046 136802 94102
rect 136858 94046 167398 94102
rect 167454 94046 167522 94102
rect 167578 94046 198118 94102
rect 198174 94046 198242 94102
rect 198298 94046 228838 94102
rect 228894 94046 228962 94102
rect 229018 94046 259558 94102
rect 259614 94046 259682 94102
rect 259738 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 374518 94102
rect 374574 94046 374642 94102
rect 374698 94046 405238 94102
rect 405294 94046 405362 94102
rect 405418 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 464518 94102
rect 464574 94046 464642 94102
rect 464698 94046 495238 94102
rect 495294 94046 495362 94102
rect 495418 94046 525958 94102
rect 526014 94046 526082 94102
rect 526138 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 44518 93978
rect 44574 93922 44642 93978
rect 44698 93922 75238 93978
rect 75294 93922 75362 93978
rect 75418 93922 105958 93978
rect 106014 93922 106082 93978
rect 106138 93922 136678 93978
rect 136734 93922 136802 93978
rect 136858 93922 167398 93978
rect 167454 93922 167522 93978
rect 167578 93922 198118 93978
rect 198174 93922 198242 93978
rect 198298 93922 228838 93978
rect 228894 93922 228962 93978
rect 229018 93922 259558 93978
rect 259614 93922 259682 93978
rect 259738 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 374518 93978
rect 374574 93922 374642 93978
rect 374698 93922 405238 93978
rect 405294 93922 405362 93978
rect 405418 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 464518 93978
rect 464574 93922 464642 93978
rect 464698 93922 495238 93978
rect 495294 93922 495362 93978
rect 495418 93922 525958 93978
rect 526014 93922 526082 93978
rect 526138 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 59878 82350
rect 59934 82294 60002 82350
rect 60058 82294 90598 82350
rect 90654 82294 90722 82350
rect 90778 82294 121318 82350
rect 121374 82294 121442 82350
rect 121498 82294 152038 82350
rect 152094 82294 152162 82350
rect 152218 82294 182758 82350
rect 182814 82294 182882 82350
rect 182938 82294 213478 82350
rect 213534 82294 213602 82350
rect 213658 82294 244198 82350
rect 244254 82294 244322 82350
rect 244378 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 389878 82350
rect 389934 82294 390002 82350
rect 390058 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 510598 82350
rect 510654 82294 510722 82350
rect 510778 82294 541318 82350
rect 541374 82294 541442 82350
rect 541498 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 59878 82226
rect 59934 82170 60002 82226
rect 60058 82170 90598 82226
rect 90654 82170 90722 82226
rect 90778 82170 121318 82226
rect 121374 82170 121442 82226
rect 121498 82170 152038 82226
rect 152094 82170 152162 82226
rect 152218 82170 182758 82226
rect 182814 82170 182882 82226
rect 182938 82170 213478 82226
rect 213534 82170 213602 82226
rect 213658 82170 244198 82226
rect 244254 82170 244322 82226
rect 244378 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 389878 82226
rect 389934 82170 390002 82226
rect 390058 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 510598 82226
rect 510654 82170 510722 82226
rect 510778 82170 541318 82226
rect 541374 82170 541442 82226
rect 541498 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82147 597980 82170
rect -1916 82102 299528 82147
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 59878 82102
rect 59934 82046 60002 82102
rect 60058 82046 90598 82102
rect 90654 82046 90722 82102
rect 90778 82046 121318 82102
rect 121374 82046 121442 82102
rect 121498 82046 152038 82102
rect 152094 82046 152162 82102
rect 152218 82046 182758 82102
rect 182814 82046 182882 82102
rect 182938 82046 213478 82102
rect 213534 82046 213602 82102
rect 213658 82046 244198 82102
rect 244254 82046 244322 82102
rect 244378 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82091 299528 82102
rect 299584 82091 299632 82147
rect 299688 82091 299736 82147
rect 299792 82091 307844 82147
rect 307900 82091 307948 82147
rect 308004 82091 308052 82147
rect 308108 82091 316160 82147
rect 316216 82091 316264 82147
rect 316320 82091 316368 82147
rect 316424 82091 324476 82147
rect 324532 82091 324580 82147
rect 324636 82091 324684 82147
rect 324740 82102 597980 82147
rect 324740 82091 347154 82102
rect 286142 82046 347154 82091
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 389878 82102
rect 389934 82046 390002 82102
rect 390058 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 510598 82102
rect 510654 82046 510722 82102
rect 510778 82046 541318 82102
rect 541374 82046 541442 82102
rect 541498 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 82043 597980 82046
rect -1916 81987 299528 82043
rect 299584 81987 299632 82043
rect 299688 81987 299736 82043
rect 299792 81987 307844 82043
rect 307900 81987 307948 82043
rect 308004 81987 308052 82043
rect 308108 81987 316160 82043
rect 316216 81987 316264 82043
rect 316320 81987 316368 82043
rect 316424 81987 324476 82043
rect 324532 81987 324580 82043
rect 324636 81987 324684 82043
rect 324740 81987 597980 82043
rect -1916 81978 597980 81987
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 59878 81978
rect 59934 81922 60002 81978
rect 60058 81922 90598 81978
rect 90654 81922 90722 81978
rect 90778 81922 121318 81978
rect 121374 81922 121442 81978
rect 121498 81922 152038 81978
rect 152094 81922 152162 81978
rect 152218 81922 182758 81978
rect 182814 81922 182882 81978
rect 182938 81922 213478 81978
rect 213534 81922 213602 81978
rect 213658 81922 244198 81978
rect 244254 81922 244322 81978
rect 244378 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81939 347154 81978
rect 286142 81922 299528 81939
rect -1916 81883 299528 81922
rect 299584 81883 299632 81939
rect 299688 81883 299736 81939
rect 299792 81883 307844 81939
rect 307900 81883 307948 81939
rect 308004 81883 308052 81939
rect 308108 81883 316160 81939
rect 316216 81883 316264 81939
rect 316320 81883 316368 81939
rect 316424 81883 324476 81939
rect 324532 81883 324580 81939
rect 324636 81883 324684 81939
rect 324740 81922 347154 81939
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 389878 81978
rect 389934 81922 390002 81978
rect 390058 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 510598 81978
rect 510654 81922 510722 81978
rect 510778 81922 541318 81978
rect 541374 81922 541442 81978
rect 541498 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 324740 81883 597980 81922
rect -1916 81826 597980 81883
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 44518 76350
rect 44574 76294 44642 76350
rect 44698 76294 75238 76350
rect 75294 76294 75362 76350
rect 75418 76294 105958 76350
rect 106014 76294 106082 76350
rect 106138 76294 136678 76350
rect 136734 76294 136802 76350
rect 136858 76294 167398 76350
rect 167454 76294 167522 76350
rect 167578 76294 198118 76350
rect 198174 76294 198242 76350
rect 198298 76294 228838 76350
rect 228894 76294 228962 76350
rect 229018 76294 259558 76350
rect 259614 76294 259682 76350
rect 259738 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 295412 76350
rect 295468 76294 295536 76350
rect 295592 76294 303728 76350
rect 303784 76294 303852 76350
rect 303908 76294 312044 76350
rect 312100 76294 312168 76350
rect 312224 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 320360 76350
rect 320416 76294 320484 76350
rect 320540 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 374518 76350
rect 374574 76294 374642 76350
rect 374698 76294 405238 76350
rect 405294 76294 405362 76350
rect 405418 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 525958 76350
rect 526014 76294 526082 76350
rect 526138 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 44518 76226
rect 44574 76170 44642 76226
rect 44698 76170 75238 76226
rect 75294 76170 75362 76226
rect 75418 76170 105958 76226
rect 106014 76170 106082 76226
rect 106138 76170 136678 76226
rect 136734 76170 136802 76226
rect 136858 76170 167398 76226
rect 167454 76170 167522 76226
rect 167578 76170 198118 76226
rect 198174 76170 198242 76226
rect 198298 76170 228838 76226
rect 228894 76170 228962 76226
rect 229018 76170 259558 76226
rect 259614 76170 259682 76226
rect 259738 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 295412 76226
rect 295468 76170 295536 76226
rect 295592 76170 303728 76226
rect 303784 76170 303852 76226
rect 303908 76170 312044 76226
rect 312100 76170 312168 76226
rect 312224 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 320360 76226
rect 320416 76170 320484 76226
rect 320540 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 374518 76226
rect 374574 76170 374642 76226
rect 374698 76170 405238 76226
rect 405294 76170 405362 76226
rect 405418 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 525958 76226
rect 526014 76170 526082 76226
rect 526138 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 44518 76102
rect 44574 76046 44642 76102
rect 44698 76046 75238 76102
rect 75294 76046 75362 76102
rect 75418 76046 105958 76102
rect 106014 76046 106082 76102
rect 106138 76046 136678 76102
rect 136734 76046 136802 76102
rect 136858 76046 167398 76102
rect 167454 76046 167522 76102
rect 167578 76046 198118 76102
rect 198174 76046 198242 76102
rect 198298 76046 228838 76102
rect 228894 76046 228962 76102
rect 229018 76046 259558 76102
rect 259614 76046 259682 76102
rect 259738 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 295412 76102
rect 295468 76046 295536 76102
rect 295592 76046 303728 76102
rect 303784 76046 303852 76102
rect 303908 76046 312044 76102
rect 312100 76046 312168 76102
rect 312224 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 320360 76102
rect 320416 76046 320484 76102
rect 320540 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 374518 76102
rect 374574 76046 374642 76102
rect 374698 76046 405238 76102
rect 405294 76046 405362 76102
rect 405418 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 525958 76102
rect 526014 76046 526082 76102
rect 526138 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 44518 75978
rect 44574 75922 44642 75978
rect 44698 75922 75238 75978
rect 75294 75922 75362 75978
rect 75418 75922 105958 75978
rect 106014 75922 106082 75978
rect 106138 75922 136678 75978
rect 136734 75922 136802 75978
rect 136858 75922 167398 75978
rect 167454 75922 167522 75978
rect 167578 75922 198118 75978
rect 198174 75922 198242 75978
rect 198298 75922 228838 75978
rect 228894 75922 228962 75978
rect 229018 75922 259558 75978
rect 259614 75922 259682 75978
rect 259738 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 295412 75978
rect 295468 75922 295536 75978
rect 295592 75922 303728 75978
rect 303784 75922 303852 75978
rect 303908 75922 312044 75978
rect 312100 75922 312168 75978
rect 312224 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 320360 75978
rect 320416 75922 320484 75978
rect 320540 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 374518 75978
rect 374574 75922 374642 75978
rect 374698 75922 405238 75978
rect 405294 75922 405362 75978
rect 405418 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 525958 75978
rect 526014 75922 526082 75978
rect 526138 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 59878 64350
rect 59934 64294 60002 64350
rect 60058 64294 90598 64350
rect 90654 64294 90722 64350
rect 90778 64294 121318 64350
rect 121374 64294 121442 64350
rect 121498 64294 152038 64350
rect 152094 64294 152162 64350
rect 152218 64294 182758 64350
rect 182814 64294 182882 64350
rect 182938 64294 213478 64350
rect 213534 64294 213602 64350
rect 213658 64294 244198 64350
rect 244254 64294 244322 64350
rect 244378 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 299570 64350
rect 299626 64294 299694 64350
rect 299750 64294 307886 64350
rect 307942 64294 308010 64350
rect 308066 64294 316202 64350
rect 316258 64294 316326 64350
rect 316382 64294 324518 64350
rect 324574 64294 324642 64350
rect 324698 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 389878 64350
rect 389934 64294 390002 64350
rect 390058 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 510598 64350
rect 510654 64294 510722 64350
rect 510778 64294 541318 64350
rect 541374 64294 541442 64350
rect 541498 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 59878 64226
rect 59934 64170 60002 64226
rect 60058 64170 90598 64226
rect 90654 64170 90722 64226
rect 90778 64170 121318 64226
rect 121374 64170 121442 64226
rect 121498 64170 152038 64226
rect 152094 64170 152162 64226
rect 152218 64170 182758 64226
rect 182814 64170 182882 64226
rect 182938 64170 213478 64226
rect 213534 64170 213602 64226
rect 213658 64170 244198 64226
rect 244254 64170 244322 64226
rect 244378 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 299570 64226
rect 299626 64170 299694 64226
rect 299750 64170 307886 64226
rect 307942 64170 308010 64226
rect 308066 64170 316202 64226
rect 316258 64170 316326 64226
rect 316382 64170 324518 64226
rect 324574 64170 324642 64226
rect 324698 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 389878 64226
rect 389934 64170 390002 64226
rect 390058 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 510598 64226
rect 510654 64170 510722 64226
rect 510778 64170 541318 64226
rect 541374 64170 541442 64226
rect 541498 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 59878 64102
rect 59934 64046 60002 64102
rect 60058 64046 90598 64102
rect 90654 64046 90722 64102
rect 90778 64046 121318 64102
rect 121374 64046 121442 64102
rect 121498 64046 152038 64102
rect 152094 64046 152162 64102
rect 152218 64046 182758 64102
rect 182814 64046 182882 64102
rect 182938 64046 213478 64102
rect 213534 64046 213602 64102
rect 213658 64046 244198 64102
rect 244254 64046 244322 64102
rect 244378 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 299570 64102
rect 299626 64046 299694 64102
rect 299750 64046 307886 64102
rect 307942 64046 308010 64102
rect 308066 64046 316202 64102
rect 316258 64046 316326 64102
rect 316382 64046 324518 64102
rect 324574 64046 324642 64102
rect 324698 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 389878 64102
rect 389934 64046 390002 64102
rect 390058 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 510598 64102
rect 510654 64046 510722 64102
rect 510778 64046 541318 64102
rect 541374 64046 541442 64102
rect 541498 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 59878 63978
rect 59934 63922 60002 63978
rect 60058 63922 90598 63978
rect 90654 63922 90722 63978
rect 90778 63922 121318 63978
rect 121374 63922 121442 63978
rect 121498 63922 152038 63978
rect 152094 63922 152162 63978
rect 152218 63922 182758 63978
rect 182814 63922 182882 63978
rect 182938 63922 213478 63978
rect 213534 63922 213602 63978
rect 213658 63922 244198 63978
rect 244254 63922 244322 63978
rect 244378 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 299570 63978
rect 299626 63922 299694 63978
rect 299750 63922 307886 63978
rect 307942 63922 308010 63978
rect 308066 63922 316202 63978
rect 316258 63922 316326 63978
rect 316382 63922 324518 63978
rect 324574 63922 324642 63978
rect 324698 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 389878 63978
rect 389934 63922 390002 63978
rect 390058 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 510598 63978
rect 510654 63922 510722 63978
rect 510778 63922 541318 63978
rect 541374 63922 541442 63978
rect 541498 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 44518 58350
rect 44574 58294 44642 58350
rect 44698 58294 75238 58350
rect 75294 58294 75362 58350
rect 75418 58294 105958 58350
rect 106014 58294 106082 58350
rect 106138 58294 136678 58350
rect 136734 58294 136802 58350
rect 136858 58294 167398 58350
rect 167454 58294 167522 58350
rect 167578 58294 198118 58350
rect 198174 58294 198242 58350
rect 198298 58294 228838 58350
rect 228894 58294 228962 58350
rect 229018 58294 259558 58350
rect 259614 58294 259682 58350
rect 259738 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 295412 58350
rect 295468 58294 295536 58350
rect 295592 58294 303728 58350
rect 303784 58294 303852 58350
rect 303908 58294 312044 58350
rect 312100 58294 312168 58350
rect 312224 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 320360 58350
rect 320416 58294 320484 58350
rect 320540 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 374518 58350
rect 374574 58294 374642 58350
rect 374698 58294 405238 58350
rect 405294 58294 405362 58350
rect 405418 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 525958 58350
rect 526014 58294 526082 58350
rect 526138 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 44518 58226
rect 44574 58170 44642 58226
rect 44698 58170 75238 58226
rect 75294 58170 75362 58226
rect 75418 58170 105958 58226
rect 106014 58170 106082 58226
rect 106138 58170 136678 58226
rect 136734 58170 136802 58226
rect 136858 58170 167398 58226
rect 167454 58170 167522 58226
rect 167578 58170 198118 58226
rect 198174 58170 198242 58226
rect 198298 58170 228838 58226
rect 228894 58170 228962 58226
rect 229018 58170 259558 58226
rect 259614 58170 259682 58226
rect 259738 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 295412 58226
rect 295468 58170 295536 58226
rect 295592 58170 303728 58226
rect 303784 58170 303852 58226
rect 303908 58170 312044 58226
rect 312100 58170 312168 58226
rect 312224 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 320360 58226
rect 320416 58170 320484 58226
rect 320540 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 374518 58226
rect 374574 58170 374642 58226
rect 374698 58170 405238 58226
rect 405294 58170 405362 58226
rect 405418 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 525958 58226
rect 526014 58170 526082 58226
rect 526138 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 44518 58102
rect 44574 58046 44642 58102
rect 44698 58046 75238 58102
rect 75294 58046 75362 58102
rect 75418 58046 105958 58102
rect 106014 58046 106082 58102
rect 106138 58046 136678 58102
rect 136734 58046 136802 58102
rect 136858 58046 167398 58102
rect 167454 58046 167522 58102
rect 167578 58046 198118 58102
rect 198174 58046 198242 58102
rect 198298 58046 228838 58102
rect 228894 58046 228962 58102
rect 229018 58046 259558 58102
rect 259614 58046 259682 58102
rect 259738 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 295412 58102
rect 295468 58046 295536 58102
rect 295592 58046 303728 58102
rect 303784 58046 303852 58102
rect 303908 58046 312044 58102
rect 312100 58046 312168 58102
rect 312224 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 320360 58102
rect 320416 58046 320484 58102
rect 320540 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 374518 58102
rect 374574 58046 374642 58102
rect 374698 58046 405238 58102
rect 405294 58046 405362 58102
rect 405418 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 525958 58102
rect 526014 58046 526082 58102
rect 526138 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 44518 57978
rect 44574 57922 44642 57978
rect 44698 57922 75238 57978
rect 75294 57922 75362 57978
rect 75418 57922 105958 57978
rect 106014 57922 106082 57978
rect 106138 57922 136678 57978
rect 136734 57922 136802 57978
rect 136858 57922 167398 57978
rect 167454 57922 167522 57978
rect 167578 57922 198118 57978
rect 198174 57922 198242 57978
rect 198298 57922 228838 57978
rect 228894 57922 228962 57978
rect 229018 57922 259558 57978
rect 259614 57922 259682 57978
rect 259738 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 295412 57978
rect 295468 57922 295536 57978
rect 295592 57922 303728 57978
rect 303784 57922 303852 57978
rect 303908 57922 312044 57978
rect 312100 57922 312168 57978
rect 312224 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 320360 57978
rect 320416 57922 320484 57978
rect 320540 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 374518 57978
rect 374574 57922 374642 57978
rect 374698 57922 405238 57978
rect 405294 57922 405362 57978
rect 405418 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 525958 57978
rect 526014 57922 526082 57978
rect 526138 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect 110780 47998 267556 48014
rect 110780 47942 110796 47998
rect 110852 47942 267484 47998
rect 267540 47942 267556 47998
rect 110780 47926 267556 47942
rect 90620 47818 270132 47834
rect 90620 47762 90636 47818
rect 90692 47762 270060 47818
rect 270116 47762 270132 47818
rect 90620 47746 270132 47762
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect 154460 44758 283124 44774
rect 154460 44702 154476 44758
rect 154532 44702 283052 44758
rect 283108 44702 283124 44758
rect 154460 44686 283124 44702
rect 104060 44578 338788 44594
rect 104060 44522 104076 44578
rect 104132 44522 338716 44578
rect 338772 44522 338788 44578
rect 104060 44506 338788 44522
rect 75500 41158 340244 41174
rect 75500 41102 75516 41158
rect 75572 41102 340172 41158
rect 340228 41102 340244 41158
rect 75500 41086 340244 41102
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect 33500 4978 57220 4994
rect 33500 4922 33516 4978
rect 33572 4922 57148 4978
rect 57204 4922 57220 4978
rect 33500 4906 57220 4922
rect 137212 4978 288388 4994
rect 137212 4922 137228 4978
rect 137284 4922 288316 4978
rect 288372 4922 288388 4978
rect 137212 4906 288388 4922
rect 35180 4798 55204 4814
rect 35180 4742 35196 4798
rect 35252 4742 55132 4798
rect 55188 4742 55204 4798
rect 35180 4726 55204 4742
rect 148636 4798 281444 4814
rect 148636 4742 148652 4798
rect 148708 4742 281372 4798
rect 281428 4742 281444 4798
rect 148636 4726 281444 4742
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use avali_logo  avali_logo
timestamp 0
transform 1 0 60000 0 1 475000
box 0 0 90000 105660
use wrapped_ay8913  ay8913
timestamp 0
transform 1 0 40000 0 1 240000
box 1120 0 51000 51000
use blinker  blinker
timestamp 0
transform 1 0 290000 0 1 50000
box 1258 0 34768 32230
use diceroll  diceroll
timestamp 0
transform 1 0 50000 0 1 315000
box 1258 3050 44662 46000
use hellorld  hellorld
timestamp 0
transform 1 0 140000 0 1 260000
box 1258 1792 26000 26000
use wrapped_mc14500  mc14500
timestamp 0
transform 1 0 300000 0 1 160000
box 1258 0 37000 37000
use multiplexer  multiplexer
timestamp 0
transform 1 0 190000 0 1 240000
box 0 0 150000 140000
use wrapped_sid  sid
timestamp 0
transform 1 0 40000 0 1 50000
box 1258 0 230000 160000
use tholin_avalonsemi_tbb1143  tbb1143
timestamp 0
transform 1 0 120000 0 1 320000
box 1258 2688 46000 43120
use ue1  ue1
timestamp 0
transform 1 0 60000 0 1 390000
box 1258 1568 24000 24000
use wrapped_pdp11  wrapped_pdp11
timestamp 0
transform 1 0 190000 0 1 410000
box 0 0 340000 156860
use wrapped_qcpu  wrapped_qcpu
timestamp 0
transform 1 0 460000 0 1 50000
box 0 1026 95000 100000
use wrapped_sn76489  wrapped_sn76489
timestamp 0
transform 1 0 370000 0 1 50000
box 0 1138 50000 50000
use wrapped_tholin_riscv  wrapped_tholin_riscv
timestamp 0
transform 1 0 355000 0 1 165000
box 0 0 228592 230000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 210574 67478 241266 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 289134 67478 337658 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 355174 67478 390964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 412556 67478 486928 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 535792 67478 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 210574 98198 472888 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 549832 98198 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 210574 128918 488368 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 210574 159638 260964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 284908 159638 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 210574 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 210574 221078 408466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 567550 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 210574 251798 240034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 380638 251798 408466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 567550 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 240034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 380638 282518 408466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 567550 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 163170 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 193230 313238 240034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 380638 313238 408466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 567550 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 408466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 567550 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 49026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 98428 374678 164250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 567550 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 49026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 98428 405398 164250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 567550 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 164250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 567550 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 394566 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 394566 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 48914 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 394566 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 164250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 394566 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 289134 71198 337658 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 355174 71198 399778 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 410574 71198 482968 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 539752 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 210574 101918 473068 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 549472 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 210574 132638 490708 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 578452 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 210574 163358 265522 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 282254 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 210574 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 210574 224798 408466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 567550 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 380638 255518 408466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 567550 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 -1644 286238 240034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 380638 286238 408466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 567550 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 -1644 316958 50964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 84316 316958 163170 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 193230 316958 240034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 380638 316958 408466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 567550 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 -1644 347678 408466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 567550 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 -1644 378398 49026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 96334 378398 164250 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 567550 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 -1644 409118 49026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 96334 409118 164250 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 567550 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 164250 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 567550 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 394566 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 394566 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 48914 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 394566 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 164250 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 394566 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 574710 382322 574710 382322 0 vdd
rlabel via4 559350 388322 559350 388322 0 vss
rlabel metal3 39816 240744 39816 240744 0 ay8913_do\[0\]
rlabel metal2 235690 379512 235690 379512 0 ay8913_do\[10\]
rlabel metal3 234472 381416 234472 381416 0 ay8913_do\[11\]
rlabel metal2 237090 379960 237090 379960 0 ay8913_do\[12\]
rlabel metal2 237706 379960 237706 379960 0 ay8913_do\[13\]
rlabel metal2 238686 379960 238686 379960 0 ay8913_do\[14\]
rlabel metal2 68040 238826 68040 238826 0 ay8913_do\[15\]
rlabel metal2 69832 239106 69832 239106 0 ay8913_do\[16\]
rlabel metal2 240450 379960 240450 379960 0 ay8913_do\[17\]
rlabel metal2 73416 238994 73416 238994 0 ay8913_do\[18\]
rlabel metal2 242046 379960 242046 379960 0 ay8913_do\[19\]
rlabel metal2 42952 239274 42952 239274 0 ay8913_do\[1\]
rlabel metal2 242410 379960 242410 379960 0 ay8913_do\[20\]
rlabel metal2 243082 379960 243082 379960 0 ay8913_do\[21\]
rlabel metal2 116760 311360 116760 311360 0 ay8913_do\[22\]
rlabel metal2 120120 310744 120120 310744 0 ay8913_do\[23\]
rlabel metal2 99960 311696 99960 311696 0 ay8913_do\[24\]
rlabel metal2 168840 311080 168840 311080 0 ay8913_do\[25\]
rlabel metal2 95368 311976 95368 311976 0 ay8913_do\[26\]
rlabel metal2 95144 312424 95144 312424 0 ay8913_do\[27\]
rlabel metal2 44744 239162 44744 239162 0 ay8913_do\[2\]
rlabel metal2 167160 311080 167160 311080 0 ay8913_do\[3\]
rlabel metal2 48328 239106 48328 239106 0 ay8913_do\[4\]
rlabel metal2 50120 238994 50120 238994 0 ay8913_do\[5\]
rlabel metal2 51912 239218 51912 239218 0 ay8913_do\[6\]
rlabel metal2 233730 379960 233730 379960 0 ay8913_do\[7\]
rlabel metal2 234346 379960 234346 379960 0 ay8913_do\[8\]
rlabel metal2 235326 379960 235326 379960 0 ay8913_do\[9\]
rlabel metal2 307944 49210 307944 49210 0 blinker_do\[0\]
rlabel metal3 190680 367234 190680 367234 0 blinker_do\[1\]
rlabel metal3 190680 368354 190680 368354 0 blinker_do\[2\]
rlabel metal3 167398 261800 167398 261800 0 custom_settings\[0\]
rlabel via4 355432 236605 355432 236605 0 custom_settings\[10\]
rlabel metal3 167566 283976 167566 283976 0 custom_settings\[11\]
rlabel metal3 188930 514920 188930 514920 0 custom_settings\[12\]
rlabel metal3 189826 522088 189826 522088 0 custom_settings\[13\]
rlabel metal4 353976 98627 353976 98627 0 custom_settings\[14\]
rlabel metal3 188986 536424 188986 536424 0 custom_settings\[15\]
rlabel metal3 188146 543592 188146 543592 0 custom_settings\[16\]
rlabel metal3 353920 284760 353920 284760 0 custom_settings\[17\]
rlabel metal3 189042 557928 189042 557928 0 custom_settings\[18\]
rlabel metal3 189042 565096 189042 565096 0 custom_settings\[19\]
rlabel metal3 92470 280392 92470 280392 0 custom_settings\[1\]
rlabel metal3 459368 115892 459368 115892 0 custom_settings\[20\]
rlabel metal3 459368 118860 459368 118860 0 custom_settings\[21\]
rlabel metal4 351064 196560 351064 196560 0 custom_settings\[22\]
rlabel metal3 459368 124684 459368 124684 0 custom_settings\[23\]
rlabel metal3 459368 127596 459368 127596 0 custom_settings\[24\]
rlabel metal3 459368 130508 459368 130508 0 custom_settings\[25\]
rlabel metal3 459368 133420 459368 133420 0 custom_settings\[26\]
rlabel metal3 459368 136332 459368 136332 0 custom_settings\[27\]
rlabel metal3 459368 139244 459368 139244 0 custom_settings\[28\]
rlabel metal3 352100 304248 352100 304248 0 custom_settings\[29\]
rlabel metal3 90888 284998 90888 284998 0 custom_settings\[2\]
rlabel metal3 459368 145068 459368 145068 0 custom_settings\[30\]
rlabel metal4 457688 147616 457688 147616 0 custom_settings\[31\]
rlabel metal3 92470 288904 92470 288904 0 custom_settings\[3\]
rlabel metal2 187992 280616 187992 280616 0 custom_settings\[4\]
rlabel metal2 449400 98112 449400 98112 0 custom_settings\[5\]
rlabel metal4 188104 284355 188104 284355 0 custom_settings\[6\]
rlabel metal4 187096 286095 187096 286095 0 custom_settings\[7\]
rlabel metal4 188104 286241 188104 286241 0 custom_settings\[8\]
rlabel metal3 167622 279944 167622 279944 0 custom_settings\[9\]
rlabel metal2 185976 372120 185976 372120 0 diceroll_do\[0\]
rlabel metal2 69720 374528 69720 374528 0 diceroll_do\[1\]
rlabel metal2 70840 362390 70840 362390 0 diceroll_do\[2\]
rlabel metal2 74648 370174 74648 370174 0 diceroll_do\[3\]
rlabel metal2 78456 374542 78456 374542 0 diceroll_do\[4\]
rlabel metal3 200760 379848 200760 379848 0 diceroll_do\[5\]
rlabel metal2 121800 372120 121800 372120 0 diceroll_do\[6\]
rlabel metal2 91560 371448 91560 371448 0 diceroll_do\[7\]
rlabel metal2 93688 370510 93688 370510 0 diceroll_do\[8\]
rlabel metal2 161336 290374 161336 290374 0 hellorld_do
rlabel metal4 201376 379890 201376 379890 0 io_in[0]
rlabel metal2 168056 407008 168056 407008 0 io_in[10]
rlabel metal2 355320 400568 355320 400568 0 io_in[11]
rlabel metal4 423304 122593 423304 122593 0 io_in[12]
rlabel metal3 593194 522536 593194 522536 0 io_in[13]
rlabel metal5 352296 143910 352296 143910 0 io_in[14]
rlabel metal3 352464 256984 352464 256984 0 io_in[15]
rlabel metal3 353682 261800 353682 261800 0 io_in[16]
rlabel metal3 351792 406728 351792 406728 0 io_in[17]
rlabel metal3 259952 406616 259952 406616 0 io_in[18]
rlabel metal2 289128 238896 289128 238896 0 io_in[19]
rlabel metal3 354298 285992 354298 285992 0 io_in[20]
rlabel metal3 186928 566104 186928 566104 0 io_in[21]
rlabel metal2 121576 593250 121576 593250 0 io_in[22]
rlabel metal2 55384 593138 55384 593138 0 io_in[23]
rlabel metal3 353920 236824 353920 236824 0 io_in[24]
rlabel metal3 3990 544824 3990 544824 0 io_in[25]
rlabel metal3 2310 502488 2310 502488 0 io_in[26]
rlabel metal2 93240 434896 93240 434896 0 io_in[27]
rlabel metal3 350504 334376 350504 334376 0 io_in[28]
rlabel metal3 2310 375704 2310 375704 0 io_in[29]
rlabel metal3 2478 333368 2478 333368 0 io_in[30]
rlabel metal3 353626 352520 353626 352520 0 io_in[31]
rlabel metal3 331576 381360 331576 381360 0 io_in[32]
rlabel metal2 336728 396970 336728 396970 0 io_in[33]
rlabel metal2 352632 154056 352632 154056 0 io_in[34]
rlabel metal3 2310 121464 2310 121464 0 io_in[35]
rlabel metal3 351512 381416 351512 381416 0 io_in[36]
rlabel metal3 336392 162414 336392 162414 0 io_in[37]
rlabel metal3 92190 242088 92190 242088 0 io_in[5]
rlabel metal5 92568 332730 92568 332730 0 io_in[6]
rlabel metal3 165928 336518 165928 336518 0 io_in[7]
rlabel metal4 355432 213493 355432 213493 0 io_in[8]
rlabel metal3 91686 259112 91686 259112 0 io_in[9]
rlabel metal3 189042 251048 189042 251048 0 io_oeb[0]
rlabel metal3 188202 262248 188202 262248 0 io_oeb[10]
rlabel metal3 593250 469672 593250 469672 0 io_oeb[11]
rlabel metal3 593138 509320 593138 509320 0 io_oeb[12]
rlabel metal3 593138 549192 593138 549192 0 io_oeb[13]
rlabel metal3 593082 588616 593082 588616 0 io_oeb[14]
rlabel metal2 540568 585578 540568 585578 0 io_oeb[15]
rlabel metal3 189826 268968 189826 268968 0 io_oeb[16]
rlabel metal3 189938 270088 189938 270088 0 io_oeb[17]
rlabel metal3 189882 271208 189882 271208 0 io_oeb[18]
rlabel metal3 189770 272328 189770 272328 0 io_oeb[19]
rlabel metal3 593082 73192 593082 73192 0 io_oeb[1]
rlabel metal2 209608 587202 209608 587202 0 io_oeb[20]
rlabel metal2 143416 588882 143416 588882 0 io_oeb[21]
rlabel metal2 77336 589722 77336 589722 0 io_oeb[22]
rlabel metal2 11032 448602 11032 448602 0 io_oeb[23]
rlabel metal4 4144 470970 4144 470970 0 io_oeb[24]
rlabel metal3 2366 516600 2366 516600 0 io_oeb[25]
rlabel metal4 4200 472752 4200 472752 0 io_oeb[26]
rlabel metal4 167160 356608 167160 356608 0 io_oeb[27]
rlabel metal3 2366 389592 2366 389592 0 io_oeb[28]
rlabel metal3 2422 347256 2422 347256 0 io_oeb[29]
rlabel metal3 190680 252826 190680 252826 0 io_oeb[2]
rlabel metal4 165480 294784 165480 294784 0 io_oeb[30]
rlabel metal3 2366 262808 2366 262808 0 io_oeb[31]
rlabel metal3 2366 220472 2366 220472 0 io_oeb[32]
rlabel metal3 2366 178024 2366 178024 0 io_oeb[33]
rlabel metal4 27720 212352 27720 212352 0 io_oeb[34]
rlabel metal3 190120 290430 190120 290430 0 io_oeb[35]
rlabel metal3 5670 51128 5670 51128 0 io_oeb[36]
rlabel metal3 2086 8792 2086 8792 0 io_oeb[37]
rlabel metal3 188706 254408 188706 254408 0 io_oeb[3]
rlabel metal3 188762 255528 188762 255528 0 io_oeb[4]
rlabel metal3 190680 256186 190680 256186 0 io_oeb[5]
rlabel metal3 188874 257768 188874 257768 0 io_oeb[6]
rlabel metal3 190680 259350 190680 259350 0 io_oeb[7]
rlabel metal3 188594 260008 188594 260008 0 io_oeb[8]
rlabel metal3 593418 390600 593418 390600 0 io_oeb[9]
rlabel metal3 593922 20552 593922 20552 0 io_out[0]
rlabel metal4 540120 410499 540120 410499 0 io_out[10]
rlabel metal2 208446 379960 208446 379960 0 io_out[11]
rlabel metal2 209286 379960 209286 379960 0 io_out[12]
rlabel metal2 209790 379960 209790 379960 0 io_out[13]
rlabel metal2 210322 379960 210322 379960 0 io_out[14]
rlabel metal2 210994 379960 210994 379960 0 io_out[15]
rlabel metal2 211806 379960 211806 379960 0 io_out[16]
rlabel metal2 212338 379960 212338 379960 0 io_out[17]
rlabel metal2 213010 379960 213010 379960 0 io_out[18]
rlabel metal2 213682 379960 213682 379960 0 io_out[19]
rlabel metal2 336952 131656 336952 131656 0 io_out[1]
rlabel metal2 214354 379960 214354 379960 0 io_out[20]
rlabel metal2 215166 379960 215166 379960 0 io_out[21]
rlabel metal2 99512 593194 99512 593194 0 io_out[22]
rlabel metal2 216370 379960 216370 379960 0 io_out[23]
rlabel metal2 217042 379960 217042 379960 0 io_out[24]
rlabel metal2 217714 379960 217714 379960 0 io_out[25]
rlabel metal2 218526 379960 218526 379960 0 io_out[26]
rlabel metal2 219058 379960 219058 379960 0 io_out[27]
rlabel metal2 219730 379960 219730 379960 0 io_out[28]
rlabel metal3 214424 379008 214424 379008 0 io_out[29]
rlabel metal3 591402 99848 591402 99848 0 io_out[2]
rlabel metal2 49560 349048 49560 349048 0 io_out[30]
rlabel metal4 214200 379400 214200 379400 0 io_out[31]
rlabel metal3 6510 234360 6510 234360 0 io_out[32]
rlabel metal3 7350 192024 7350 192024 0 io_out[33]
rlabel metal2 24360 266392 24360 266392 0 io_out[34]
rlabel metal4 31080 243081 31080 243081 0 io_out[35]
rlabel metal4 29400 221193 29400 221193 0 io_out[36]
rlabel metal3 2310 22904 2310 22904 0 io_out[37]
rlabel metal3 591514 139384 591514 139384 0 io_out[3]
rlabel metal3 590562 179144 590562 179144 0 io_out[4]
rlabel metal3 593978 218792 593978 218792 0 io_out[5]
rlabel metal3 593082 258440 593082 258440 0 io_out[6]
rlabel metal3 593138 298088 593138 298088 0 io_out[7]
rlabel metal3 593250 337624 593250 337624 0 io_out[8]
rlabel metal2 206962 379960 206962 379960 0 io_out[9]
rlabel metal3 189602 321608 189602 321608 0 mc14500_do\[0\]
rlabel metal3 188258 332808 188258 332808 0 mc14500_do\[10\]
rlabel metal3 189658 333928 189658 333928 0 mc14500_do\[11\]
rlabel metal3 185570 335048 185570 335048 0 mc14500_do\[12\]
rlabel metal3 186522 336168 186522 336168 0 mc14500_do\[13\]
rlabel metal3 187306 337288 187306 337288 0 mc14500_do\[14\]
rlabel metal2 181272 280616 181272 280616 0 mc14500_do\[15\]
rlabel metal2 179592 282128 179592 282128 0 mc14500_do\[16\]
rlabel metal2 179368 285992 179368 285992 0 mc14500_do\[17\]
rlabel metal3 252280 233128 252280 233128 0 mc14500_do\[18\]
rlabel metal2 181160 286328 181160 286328 0 mc14500_do\[19\]
rlabel metal3 188202 322728 188202 322728 0 mc14500_do\[1\]
rlabel metal2 179704 283304 179704 283304 0 mc14500_do\[20\]
rlabel metal2 177800 286608 177800 286608 0 mc14500_do\[21\]
rlabel metal2 326312 209062 326312 209062 0 mc14500_do\[22\]
rlabel metal2 327432 214102 327432 214102 0 mc14500_do\[23\]
rlabel metal2 328552 215838 328552 215838 0 mc14500_do\[24\]
rlabel metal3 187432 349552 187432 349552 0 mc14500_do\[25\]
rlabel metal3 189714 350728 189714 350728 0 mc14500_do\[26\]
rlabel metal2 331912 214998 331912 214998 0 mc14500_do\[27\]
rlabel metal2 333032 213318 333032 213318 0 mc14500_do\[28\]
rlabel metal2 334152 212478 334152 212478 0 mc14500_do\[29\]
rlabel metal2 303912 208278 303912 208278 0 mc14500_do\[2\]
rlabel metal2 335272 214046 335272 214046 0 mc14500_do\[30\]
rlabel metal2 305032 209958 305032 209958 0 mc14500_do\[3\]
rlabel metal2 306152 209118 306152 209118 0 mc14500_do\[4\]
rlabel metal2 307272 215894 307272 215894 0 mc14500_do\[5\]
rlabel metal2 308392 215110 308392 215110 0 mc14500_do\[6\]
rlabel metal2 309512 206486 309512 206486 0 mc14500_do\[7\]
rlabel metal2 310632 213486 310632 213486 0 mc14500_do\[8\]
rlabel metal2 172984 278264 172984 278264 0 mc14500_do\[9\]
rlabel metal2 301602 160664 301602 160664 0 mc14500_sram_addr\[0\]
rlabel metal2 303170 160440 303170 160440 0 mc14500_sram_addr\[1\]
rlabel metal2 304682 160552 304682 160552 0 mc14500_sram_addr\[2\]
rlabel metal4 306600 157637 306600 157637 0 mc14500_sram_addr\[3\]
rlabel metal2 308168 158522 308168 158522 0 mc14500_sram_addr\[4\]
rlabel metal2 309736 158466 309736 158466 0 mc14500_sram_addr\[5\]
rlabel metal4 336000 193230 336000 193230 0 mc14500_sram_gwe
rlabel metal2 311304 158914 311304 158914 0 mc14500_sram_in\[0\]
rlabel metal2 312872 158746 312872 158746 0 mc14500_sram_in\[1\]
rlabel metal2 329336 222082 329336 222082 0 mc14500_sram_in\[2\]
rlabel metal2 330232 218890 330232 218890 0 mc14500_sram_in\[3\]
rlabel metal2 331128 219562 331128 219562 0 mc14500_sram_in\[4\]
rlabel metal2 332024 218722 332024 218722 0 mc14500_sram_in\[5\]
rlabel metal2 332920 220458 332920 220458 0 mc14500_sram_in\[6\]
rlabel metal2 334264 238504 334264 238504 0 mc14500_sram_in\[7\]
rlabel metal2 248318 379960 248318 379960 0 pdp11_do\[0\]
rlabel metal2 261758 379960 261758 379960 0 pdp11_do\[10\]
rlabel metal2 262738 379960 262738 379960 0 pdp11_do\[11\]
rlabel metal2 264082 379960 264082 379960 0 pdp11_do\[12\]
rlabel metal2 265566 379960 265566 379960 0 pdp11_do\[13\]
rlabel metal2 266770 379960 266770 379960 0 pdp11_do\[14\]
rlabel metal2 379624 408408 379624 408408 0 pdp11_do\[15\]
rlabel metal4 444920 407549 444920 407549 0 pdp11_do\[16\]
rlabel metal2 397320 401968 397320 401968 0 pdp11_do\[17\]
rlabel metal2 455224 408898 455224 408898 0 pdp11_do\[18\]
rlabel metal2 273490 379960 273490 379960 0 pdp11_do\[19\]
rlabel metal4 356552 400247 356552 400247 0 pdp11_do\[1\]
rlabel metal2 274834 379960 274834 379960 0 pdp11_do\[20\]
rlabel metal2 470680 402906 470680 402906 0 pdp11_do\[21\]
rlabel metal2 475832 402850 475832 402850 0 pdp11_do\[22\]
rlabel metal2 279174 379960 279174 379960 0 pdp11_do\[23\]
rlabel metal2 280210 379960 280210 379960 0 pdp11_do\[24\]
rlabel metal2 281694 379960 281694 379960 0 pdp11_do\[25\]
rlabel metal2 283206 379960 283206 379960 0 pdp11_do\[26\]
rlabel metal2 284242 379960 284242 379960 0 pdp11_do\[27\]
rlabel metal2 285894 379960 285894 379960 0 pdp11_do\[28\]
rlabel metal2 286930 379960 286930 379960 0 pdp11_do\[29\]
rlabel metal2 355544 399336 355544 399336 0 pdp11_do\[2\]
rlabel metal2 288274 379960 288274 379960 0 pdp11_do\[30\]
rlabel metal2 289982 379960 289982 379960 0 pdp11_do\[31\]
rlabel metal4 353640 397199 353640 397199 0 pdp11_do\[32\]
rlabel metal2 377944 409010 377944 409010 0 pdp11_do\[3\]
rlabel metal2 355096 392336 355096 392336 0 pdp11_do\[4\]
rlabel metal2 257880 393904 257880 393904 0 pdp11_do\[5\]
rlabel metal2 256382 379960 256382 379960 0 pdp11_do\[6\]
rlabel metal2 257726 379960 257726 379960 0 pdp11_do\[7\]
rlabel metal2 259014 379960 259014 379960 0 pdp11_do\[8\]
rlabel metal2 260246 379960 260246 379960 0 pdp11_do\[9\]
rlabel metal2 248766 379960 248766 379960 0 pdp11_oeb\[0\]
rlabel metal2 262206 379960 262206 379960 0 pdp11_oeb\[10\]
rlabel metal2 263410 379960 263410 379960 0 pdp11_oeb\[11\]
rlabel metal2 264754 379960 264754 379960 0 pdp11_oeb\[12\]
rlabel metal2 266406 379960 266406 379960 0 pdp11_oeb\[13\]
rlabel metal2 267442 379960 267442 379960 0 pdp11_oeb\[14\]
rlabel metal2 268926 379960 268926 379960 0 pdp11_oeb\[15\]
rlabel metal2 270130 379960 270130 379960 0 pdp11_oeb\[16\]
rlabel metal2 271474 379960 271474 379960 0 pdp11_oeb\[17\]
rlabel metal2 272818 379960 272818 379960 0 pdp11_oeb\[18\]
rlabel metal2 274162 379960 274162 379960 0 pdp11_oeb\[19\]
rlabel metal2 249970 379960 249970 379960 0 pdp11_oeb\[1\]
rlabel metal2 275646 379960 275646 379960 0 pdp11_oeb\[20\]
rlabel metal2 276850 379960 276850 379960 0 pdp11_oeb\[21\]
rlabel metal2 278194 379960 278194 379960 0 pdp11_oeb\[22\]
rlabel metal2 279538 379960 279538 379960 0 pdp11_oeb\[23\]
rlabel metal2 280882 379960 280882 379960 0 pdp11_oeb\[24\]
rlabel metal2 282366 379960 282366 379960 0 pdp11_oeb\[25\]
rlabel metal2 283570 379960 283570 379960 0 pdp11_oeb\[26\]
rlabel metal2 285278 379960 285278 379960 0 pdp11_oeb\[27\]
rlabel metal2 286258 379960 286258 379960 0 pdp11_oeb\[28\]
rlabel metal2 287910 379960 287910 379960 0 pdp11_oeb\[29\]
rlabel metal2 251314 379960 251314 379960 0 pdp11_oeb\[2\]
rlabel metal2 289310 379960 289310 379960 0 pdp11_oeb\[30\]
rlabel metal2 290486 379960 290486 379960 0 pdp11_oeb\[31\]
rlabel metal2 291998 379960 291998 379960 0 pdp11_oeb\[32\]
rlabel metal4 446040 417441 446040 417441 0 pdp11_oeb\[3\]
rlabel metal2 261240 394072 261240 394072 0 pdp11_oeb\[4\]
rlabel metal2 255710 379960 255710 379960 0 pdp11_oeb\[5\]
rlabel metal2 256886 379960 256886 379960 0 pdp11_oeb\[6\]
rlabel metal2 258398 379960 258398 379960 0 pdp11_oeb\[7\]
rlabel metal2 259378 379960 259378 379960 0 pdp11_oeb\[8\]
rlabel metal2 261086 379960 261086 379960 0 pdp11_oeb\[9\]
rlabel metal2 279160 196154 279160 196154 0 qcpu_do\[0\]
rlabel metal2 288190 240072 288190 240072 0 qcpu_do\[10\]
rlabel metal2 289016 195482 289016 195482 0 qcpu_do\[11\]
rlabel metal4 494536 149240 494536 149240 0 qcpu_do\[12\]
rlabel metal2 525448 152838 525448 152838 0 qcpu_do\[13\]
rlabel metal2 291704 198002 291704 198002 0 qcpu_do\[14\]
rlabel metal2 292600 197834 292600 197834 0 qcpu_do\[15\]
rlabel metal2 293496 197778 293496 197778 0 qcpu_do\[16\]
rlabel metal2 520856 152152 520856 152152 0 qcpu_do\[17\]
rlabel metal2 295288 196434 295288 196434 0 qcpu_do\[18\]
rlabel metal2 524216 151592 524216 151592 0 qcpu_do\[19\]
rlabel metal2 280056 196378 280056 196378 0 qcpu_do\[1\]
rlabel metal2 297080 197722 297080 197722 0 qcpu_do\[20\]
rlabel metal2 297976 195426 297976 195426 0 qcpu_do\[21\]
rlabel metal2 522536 156632 522536 156632 0 qcpu_do\[22\]
rlabel metal2 538888 152222 538888 152222 0 qcpu_do\[23\]
rlabel metal2 540232 152166 540232 152166 0 qcpu_do\[24\]
rlabel metal2 541576 152110 541576 152110 0 qcpu_do\[25\]
rlabel metal2 302456 238714 302456 238714 0 qcpu_do\[26\]
rlabel metal2 303352 238938 303352 238938 0 qcpu_do\[27\]
rlabel metal3 303856 236936 303856 236936 0 qcpu_do\[28\]
rlabel metal2 305144 238770 305144 238770 0 qcpu_do\[29\]
rlabel metal3 284704 236936 284704 236936 0 qcpu_do\[2\]
rlabel metal2 306040 238658 306040 238658 0 qcpu_do\[30\]
rlabel metal2 307384 238504 307384 238504 0 qcpu_do\[31\]
rlabel metal2 307832 238994 307832 238994 0 qcpu_do\[32\]
rlabel metal2 281848 200130 281848 200130 0 qcpu_do\[3\]
rlabel metal2 282744 238770 282744 238770 0 qcpu_do\[4\]
rlabel metal2 283640 200186 283640 200186 0 qcpu_do\[5\]
rlabel metal2 284536 200354 284536 200354 0 qcpu_do\[6\]
rlabel metal2 285432 196098 285432 196098 0 qcpu_do\[7\]
rlabel metal3 494760 149072 494760 149072 0 qcpu_do\[8\]
rlabel metal2 287224 238826 287224 238826 0 qcpu_do\[9\]
rlabel metal3 354872 183400 354872 183400 0 qcpu_oeb\[0\]
rlabel metal4 421624 155417 421624 155417 0 qcpu_oeb\[10\]
rlabel metal3 345240 262360 345240 262360 0 qcpu_oeb\[11\]
rlabel metal2 420840 159488 420840 159488 0 qcpu_oeb\[12\]
rlabel metal4 468664 156184 468664 156184 0 qcpu_oeb\[13\]
rlabel metal4 346360 160915 346360 160915 0 qcpu_oeb\[14\]
rlabel metal3 344624 262136 344624 262136 0 qcpu_oeb\[15\]
rlabel metal4 342104 150407 342104 150407 0 qcpu_oeb\[16\]
rlabel metal3 403480 149352 403480 149352 0 qcpu_oeb\[17\]
rlabel metal5 452704 150570 452704 150570 0 qcpu_oeb\[18\]
rlabel metal3 558208 147896 558208 147896 0 qcpu_oeb\[19\]
rlabel metal3 345800 256984 345800 256984 0 qcpu_oeb\[1\]
rlabel metal3 556486 88088 556486 88088 0 qcpu_oeb\[20\]
rlabel metal3 507416 161560 507416 161560 0 qcpu_oeb\[21\]
rlabel metal3 340998 326536 340998 326536 0 qcpu_oeb\[22\]
rlabel metal3 403704 147448 403704 147448 0 qcpu_oeb\[23\]
rlabel metal4 342664 240390 342664 240390 0 qcpu_oeb\[24\]
rlabel metal3 405776 140952 405776 140952 0 qcpu_oeb\[25\]
rlabel metal3 339864 329770 339864 329770 0 qcpu_oeb\[26\]
rlabel metal3 558040 143528 558040 143528 0 qcpu_oeb\[27\]
rlabel metal3 507024 163128 507024 163128 0 qcpu_oeb\[28\]
rlabel metal3 346696 280504 346696 280504 0 qcpu_oeb\[29\]
rlabel metal3 452424 50232 452424 50232 0 qcpu_oeb\[2\]
rlabel metal3 344302 333704 344302 333704 0 qcpu_oeb\[30\]
rlabel metal3 343238 334600 343238 334600 0 qcpu_oeb\[31\]
rlabel metal3 343350 335496 343350 335496 0 qcpu_oeb\[32\]
rlabel metal3 454328 50120 454328 50120 0 qcpu_oeb\[3\]
rlabel metal3 340662 310408 340662 310408 0 qcpu_oeb\[4\]
rlabel metal3 341768 241976 341768 241976 0 qcpu_oeb\[5\]
rlabel metal3 345408 283864 345408 283864 0 qcpu_oeb\[6\]
rlabel metal3 345366 313096 345366 313096 0 qcpu_oeb\[7\]
rlabel metal3 340606 313992 340606 313992 0 qcpu_oeb\[8\]
rlabel metal3 555926 70840 555926 70840 0 qcpu_oeb\[9\]
rlabel metal2 309064 238504 309064 238504 0 qcpu_sram_addr\[0\]
rlabel metal3 310184 236936 310184 236936 0 qcpu_sram_addr\[1\]
rlabel metal2 310520 219002 310520 219002 0 qcpu_sram_addr\[2\]
rlabel metal2 311416 218946 311416 218946 0 qcpu_sram_addr\[3\]
rlabel metal2 312312 218778 312312 218778 0 qcpu_sram_addr\[4\]
rlabel metal2 313208 220570 313208 220570 0 qcpu_sram_addr\[5\]
rlabel metal2 314104 238938 314104 238938 0 qcpu_sram_gwe
rlabel metal3 555646 117880 555646 117880 0 qcpu_sram_in\[0\]
rlabel metal3 554904 119854 554904 119854 0 qcpu_sram_in\[1\]
rlabel metal5 401128 139410 401128 139410 0 qcpu_sram_in\[2\]
rlabel metal3 318416 236936 318416 236936 0 qcpu_sram_in\[3\]
rlabel metal3 331856 195832 331856 195832 0 qcpu_sram_in\[4\]
rlabel metal3 554680 125846 554680 125846 0 qcpu_sram_in\[5\]
rlabel metal2 337176 193704 337176 193704 0 qcpu_sram_in\[6\]
rlabel metal2 337400 195216 337400 195216 0 qcpu_sram_in\[7\]
rlabel metal3 339864 336210 339864 336210 0 qcpu_sram_out\[0\]
rlabel metal2 341208 243544 341208 243544 0 qcpu_sram_out\[1\]
rlabel metal2 326984 158802 326984 158802 0 qcpu_sram_out\[2\]
rlabel metal2 328552 158746 328552 158746 0 qcpu_sram_out\[3\]
rlabel metal2 330120 158522 330120 158522 0 qcpu_sram_out\[4\]
rlabel metal2 331688 158690 331688 158690 0 qcpu_sram_out\[5\]
rlabel metal2 333256 158914 333256 158914 0 qcpu_sram_out\[6\]
rlabel metal2 334824 158858 334824 158858 0 qcpu_sram_out\[7\]
rlabel metal4 237832 347383 237832 347383 0 rst_ay8913
rlabel metal3 190680 364938 190680 364938 0 rst_blinker
rlabel metal2 315294 379960 315294 379960 0 rst_diceroll
rlabel metal2 167272 339080 167272 339080 0 rst_hellorld
rlabel metal3 338366 165032 338366 165032 0 rst_mc14500
rlabel metal3 189770 421736 189770 421736 0 rst_pdp11
rlabel metal4 190680 319299 190680 319299 0 rst_qcpu
rlabel metal2 212296 48930 212296 48930 0 rst_sid
rlabel metal2 337064 143808 337064 143808 0 rst_sn76489
rlabel metal3 167454 326088 167454 326088 0 rst_tbb1143
rlabel metal2 292670 379960 292670 379960 0 rst_tholin_riscv
rlabel metal2 211624 392784 211624 392784 0 rst_ue1
rlabel metal3 188090 294728 188090 294728 0 sid_do\[0\]
rlabel metal3 186410 305928 186410 305928 0 sid_do\[10\]
rlabel metal3 185626 307048 185626 307048 0 sid_do\[11\]
rlabel metal3 189826 308168 189826 308168 0 sid_do\[12\]
rlabel metal3 185570 309288 185570 309288 0 sid_do\[13\]
rlabel metal4 190456 267680 190456 267680 0 sid_do\[14\]
rlabel metal3 187250 311528 187250 311528 0 sid_do\[15\]
rlabel metal3 184898 312648 184898 312648 0 sid_do\[16\]
rlabel metal3 184058 313768 184058 313768 0 sid_do\[17\]
rlabel metal3 188258 314888 188258 314888 0 sid_do\[18\]
rlabel metal3 227024 211064 227024 211064 0 sid_do\[19\]
rlabel metal3 188986 295848 188986 295848 0 sid_do\[1\]
rlabel metal3 269864 210896 269864 210896 0 sid_do\[20\]
rlabel metal3 188538 296968 188538 296968 0 sid_do\[2\]
rlabel metal3 272776 209832 272776 209832 0 sid_do\[3\]
rlabel metal3 188818 299208 188818 299208 0 sid_do\[4\]
rlabel metal3 188650 300328 188650 300328 0 sid_do\[5\]
rlabel metal3 271278 166264 271278 166264 0 sid_do\[6\]
rlabel metal3 189042 302568 189042 302568 0 sid_do\[7\]
rlabel metal3 188930 303688 188930 303688 0 sid_do\[8\]
rlabel metal3 188146 304808 188146 304808 0 sid_do\[9\]
rlabel metal2 167272 267960 167272 267960 0 sid_oeb
rlabel metal2 373338 99960 373338 99960 0 sn76489_do\[0\]
rlabel metal2 263032 225386 263032 225386 0 sn76489_do\[10\]
rlabel metal2 263928 225778 263928 225778 0 sn76489_do\[11\]
rlabel metal4 264824 209552 264824 209552 0 sn76489_do\[12\]
rlabel metal2 265720 225834 265720 225834 0 sn76489_do\[13\]
rlabel metal2 267064 238504 267064 238504 0 sn76489_do\[14\]
rlabel metal2 396858 99960 396858 99960 0 sn76489_do\[15\]
rlabel metal2 398482 99960 398482 99960 0 sn76489_do\[16\]
rlabel metal2 400274 99960 400274 99960 0 sn76489_do\[17\]
rlabel metal2 401842 99960 401842 99960 0 sn76489_do\[18\]
rlabel metal2 403410 99960 403410 99960 0 sn76489_do\[19\]
rlabel metal2 374962 99960 374962 99960 0 sn76489_do\[1\]
rlabel metal2 404978 99960 404978 99960 0 sn76489_do\[20\]
rlabel metal2 406686 99960 406686 99960 0 sn76489_do\[21\]
rlabel metal2 408114 99960 408114 99960 0 sn76489_do\[22\]
rlabel metal2 406616 103768 406616 103768 0 sn76489_do\[23\]
rlabel metal2 411250 99960 411250 99960 0 sn76489_do\[24\]
rlabel metal2 412818 99960 412818 99960 0 sn76489_do\[25\]
rlabel metal2 414386 99960 414386 99960 0 sn76489_do\[26\]
rlabel metal2 415954 99960 415954 99960 0 sn76489_do\[27\]
rlabel metal2 376698 99960 376698 99960 0 sn76489_do\[2\]
rlabel metal2 378210 99960 378210 99960 0 sn76489_do\[3\]
rlabel metal2 379834 99960 379834 99960 0 sn76489_do\[4\]
rlabel metal2 381458 99960 381458 99960 0 sn76489_do\[5\]
rlabel metal2 383166 99960 383166 99960 0 sn76489_do\[6\]
rlabel metal2 384314 99960 384314 99960 0 sn76489_do\[7\]
rlabel metal2 261240 224994 261240 224994 0 sn76489_do\[8\]
rlabel metal2 262136 228354 262136 228354 0 sn76489_do\[9\]
rlabel metal4 186424 354648 186424 354648 0 tbb1143_do\[0\]
rlabel metal4 179816 356888 179816 356888 0 tbb1143_do\[1\]
rlabel metal3 166502 356328 166502 356328 0 tbb1143_do\[2\]
rlabel metal3 188314 363048 188314 363048 0 tbb1143_do\[3\]
rlabel metal3 165928 363174 165928 363174 0 tbb1143_do\[4\]
rlabel metal2 358232 163968 358232 163968 0 tholin_riscv_do\[0\]
rlabel metal2 427672 164640 427672 164640 0 tholin_riscv_do\[10\]
rlabel metal3 345254 355208 345254 355208 0 tholin_riscv_do\[11\]
rlabel metal3 340886 356104 340886 356104 0 tholin_riscv_do\[12\]
rlabel metal2 448616 163912 448616 163912 0 tholin_riscv_do\[13\]
rlabel metal3 342566 357896 342566 357896 0 tholin_riscv_do\[14\]
rlabel metal3 345198 358792 345198 358792 0 tholin_riscv_do\[15\]
rlabel metal2 469336 163744 469336 163744 0 tholin_riscv_do\[16\]
rlabel metal2 477064 163968 477064 163968 0 tholin_riscv_do\[17\]
rlabel metal2 483966 165032 483966 165032 0 tholin_riscv_do\[18\]
rlabel metal2 490728 163520 490728 163520 0 tholin_riscv_do\[19\]
rlabel metal3 357448 165144 357448 165144 0 tholin_riscv_do\[1\]
rlabel metal2 497896 163968 497896 163968 0 tholin_riscv_do\[20\]
rlabel metal2 504056 164752 504056 164752 0 tholin_riscv_do\[21\]
rlabel metal2 511602 165032 511602 165032 0 tholin_riscv_do\[22\]
rlabel metal2 517944 164360 517944 164360 0 tholin_riscv_do\[23\]
rlabel metal2 525490 165032 525490 165032 0 tholin_riscv_do\[24\]
rlabel metal2 532392 163968 532392 163968 0 tholin_riscv_do\[25\]
rlabel metal4 539336 162857 539336 162857 0 tholin_riscv_do\[26\]
rlabel metal2 546504 163968 546504 163968 0 tholin_riscv_do\[27\]
rlabel metal3 450968 165032 450968 165032 0 tholin_riscv_do\[28\]
rlabel metal4 584808 278969 584808 278969 0 tholin_riscv_do\[29\]
rlabel metal2 372120 163744 372120 163744 0 tholin_riscv_do\[2\]
rlabel metal2 567784 163912 567784 163912 0 tholin_riscv_do\[30\]
rlabel metal4 586376 280645 586376 280645 0 tholin_riscv_do\[31\]
rlabel metal4 586488 279943 586488 279943 0 tholin_riscv_do\[32\]
rlabel metal2 379848 164808 379848 164808 0 tholin_riscv_do\[3\]
rlabel metal2 386610 165032 386610 165032 0 tholin_riscv_do\[4\]
rlabel metal3 346878 349832 346878 349832 0 tholin_riscv_do\[5\]
rlabel metal2 399896 164584 399896 164584 0 tholin_riscv_do\[6\]
rlabel metal2 407442 165032 407442 165032 0 tholin_riscv_do\[7\]
rlabel metal3 340942 352520 340942 352520 0 tholin_riscv_do\[8\]
rlabel metal2 421330 165032 421330 165032 0 tholin_riscv_do\[9\]
rlabel metal4 356664 392975 356664 392975 0 tholin_riscv_oeb\[0\]
rlabel metal2 427994 394968 427994 394968 0 tholin_riscv_oeb\[10\]
rlabel metal2 421624 399504 421624 399504 0 tholin_riscv_oeb\[11\]
rlabel metal2 350504 391384 350504 391384 0 tholin_riscv_oeb\[12\]
rlabel metal2 429240 395752 429240 395752 0 tholin_riscv_oeb\[13\]
rlabel metal2 302526 379960 302526 379960 0 tholin_riscv_oeb\[14\]
rlabel metal2 303366 379960 303366 379960 0 tholin_riscv_oeb\[15\]
rlabel metal2 303730 379960 303730 379960 0 tholin_riscv_oeb\[16\]
rlabel metal2 304402 379960 304402 379960 0 tholin_riscv_oeb\[17\]
rlabel metal2 305074 379960 305074 379960 0 tholin_riscv_oeb\[18\]
rlabel metal2 305886 379960 305886 379960 0 tholin_riscv_oeb\[19\]
rlabel metal2 355208 393176 355208 393176 0 tholin_riscv_oeb\[1\]
rlabel metal2 306726 379960 306726 379960 0 tholin_riscv_oeb\[20\]
rlabel metal2 307090 379960 307090 379960 0 tholin_riscv_oeb\[21\]
rlabel metal2 307762 379960 307762 379960 0 tholin_riscv_oeb\[22\]
rlabel metal2 308434 379960 308434 379960 0 tholin_riscv_oeb\[23\]
rlabel metal2 309246 379960 309246 379960 0 tholin_riscv_oeb\[24\]
rlabel metal2 309778 379960 309778 379960 0 tholin_riscv_oeb\[25\]
rlabel metal2 310450 379960 310450 379960 0 tholin_riscv_oeb\[26\]
rlabel metal2 311122 379960 311122 379960 0 tholin_riscv_oeb\[27\]
rlabel metal2 312158 379960 312158 379960 0 tholin_riscv_oeb\[28\]
rlabel metal2 312830 379960 312830 379960 0 tholin_riscv_oeb\[29\]
rlabel metal2 354872 394184 354872 394184 0 tholin_riscv_oeb\[2\]
rlabel metal2 313446 379960 313446 379960 0 tholin_riscv_oeb\[30\]
rlabel metal2 313810 379960 313810 379960 0 tholin_riscv_oeb\[31\]
rlabel metal4 356104 394020 356104 394020 0 tholin_riscv_oeb\[32\]
rlabel metal4 379848 393960 379848 393960 0 tholin_riscv_oeb\[3\]
rlabel metal2 354984 394240 354984 394240 0 tholin_riscv_oeb\[4\]
rlabel metal2 355432 392504 355432 392504 0 tholin_riscv_oeb\[5\]
rlabel metal2 400386 394968 400386 394968 0 tholin_riscv_oeb\[6\]
rlabel metal2 354760 391048 354760 391048 0 tholin_riscv_oeb\[7\]
rlabel metal2 403144 395640 403144 395640 0 tholin_riscv_oeb\[8\]
rlabel metal2 421050 394968 421050 394968 0 tholin_riscv_oeb\[9\]
rlabel metal2 323106 379960 323106 379960 0 ue1_do\[0\]
rlabel metal3 86016 397544 86016 397544 0 ue1_do\[1\]
rlabel metal2 324562 379960 324562 379960 0 ue1_do\[2\]
rlabel metal2 68600 415702 68600 415702 0 ue1_do\[3\]
rlabel metal2 326046 379960 326046 379960 0 ue1_do\[4\]
rlabel metal2 326466 379960 326466 379960 0 ue1_do\[5\]
rlabel metal2 327250 379960 327250 379960 0 ue1_do\[6\]
rlabel metal2 327810 379960 327810 379960 0 ue1_do\[7\]
rlabel metal2 328594 379960 328594 379960 0 ue1_do\[8\]
rlabel metal2 329406 379960 329406 379960 0 ue1_do\[9\]
rlabel metal2 185640 398776 185640 398776 0 ue1_oeb
rlabel metal4 584696 199907 584696 199907 0 user_irq[0]
rlabel metal2 336840 108472 336840 108472 0 user_irq[1]
rlabel metal2 284984 109200 284984 109200 0 user_irq[2]
rlabel metal3 46984 47040 46984 47040 0 wb_clk_i
rlabel metal2 195832 232162 195832 232162 0 wb_rst_i
rlabel metal2 15400 2310 15400 2310 0 wbs_ack_o
rlabel metal2 22792 116662 22792 116662 0 wbs_adr_i[0]
rlabel metal3 64288 49560 64288 49560 0 wbs_adr_i[10]
rlabel metal2 93240 2366 93240 2366 0 wbs_adr_i[11]
rlabel metal2 98952 2310 98952 2310 0 wbs_adr_i[12]
rlabel metal3 209160 236936 209160 236936 0 wbs_adr_i[13]
rlabel metal2 209272 235802 209272 235802 0 wbs_adr_i[14]
rlabel metal2 116312 2366 116312 2366 0 wbs_adr_i[15]
rlabel metal2 121800 24150 121800 24150 0 wbs_adr_i[16]
rlabel metal2 211960 235858 211960 235858 0 wbs_adr_i[17]
rlabel metal2 212856 235466 212856 235466 0 wbs_adr_i[18]
rlabel metal2 138936 24318 138936 24318 0 wbs_adr_i[19]
rlabel metal2 30408 106526 30408 106526 0 wbs_adr_i[1]
rlabel metal2 144648 25102 144648 25102 0 wbs_adr_i[20]
rlabel metal2 215544 234178 215544 234178 0 wbs_adr_i[21]
rlabel metal2 216440 234234 216440 234234 0 wbs_adr_i[22]
rlabel metal2 161784 25270 161784 25270 0 wbs_adr_i[23]
rlabel metal2 167496 22638 167496 22638 0 wbs_adr_i[24]
rlabel metal2 219128 232554 219128 232554 0 wbs_adr_i[25]
rlabel metal2 220024 232162 220024 232162 0 wbs_adr_i[26]
rlabel metal3 230328 45192 230328 45192 0 wbs_adr_i[27]
rlabel metal2 190344 22862 190344 22862 0 wbs_adr_i[28]
rlabel metal2 196056 24374 196056 24374 0 wbs_adr_i[29]
rlabel metal2 38024 114086 38024 114086 0 wbs_adr_i[2]
rlabel metal4 266952 141512 266952 141512 0 wbs_adr_i[30]
rlabel metal3 241808 44408 241808 44408 0 wbs_adr_i[31]
rlabel metal2 45640 25270 45640 25270 0 wbs_adr_i[3]
rlabel metal2 53256 24318 53256 24318 0 wbs_adr_i[4]
rlabel metal2 58968 2254 58968 2254 0 wbs_adr_i[5]
rlabel metal2 64680 2646 64680 2646 0 wbs_adr_i[6]
rlabel metal2 70392 2422 70392 2422 0 wbs_adr_i[7]
rlabel metal2 76104 2534 76104 2534 0 wbs_adr_i[8]
rlabel metal3 61320 47992 61320 47992 0 wbs_adr_i[9]
rlabel metal3 351568 261240 351568 261240 0 wbs_cyc_i
rlabel metal2 24696 107310 24696 107310 0 wbs_dat_i[0]
rlabel metal2 234360 237146 234360 237146 0 wbs_dat_i[10]
rlabel metal3 236040 237048 236040 237048 0 wbs_dat_i[11]
rlabel metal2 236712 238504 236712 238504 0 wbs_dat_i[12]
rlabel metal3 237776 236936 237776 236936 0 wbs_dat_i[13]
rlabel metal2 237944 236418 237944 236418 0 wbs_dat_i[14]
rlabel metal3 239456 236936 239456 236936 0 wbs_dat_i[15]
rlabel metal2 239736 236474 239736 236474 0 wbs_dat_i[16]
rlabel metal3 241248 236936 241248 236936 0 wbs_dat_i[17]
rlabel metal2 241528 226674 241528 226674 0 wbs_dat_i[18]
rlabel metal3 242928 237048 242928 237048 0 wbs_dat_i[19]
rlabel metal2 32536 2310 32536 2310 0 wbs_dat_i[1]
rlabel metal2 243544 238504 243544 238504 0 wbs_dat_i[20]
rlabel metal4 244216 237737 244216 237737 0 wbs_dat_i[21]
rlabel metal2 158200 3150 158200 3150 0 wbs_dat_i[22]
rlabel metal2 163912 3990 163912 3990 0 wbs_dat_i[23]
rlabel metal2 169400 14910 169400 14910 0 wbs_dat_i[24]
rlabel metal2 280616 140616 280616 140616 0 wbs_dat_i[25]
rlabel metal2 248696 238994 248696 238994 0 wbs_dat_i[26]
rlabel metal2 186536 15750 186536 15750 0 wbs_dat_i[27]
rlabel metal2 192248 6510 192248 6510 0 wbs_dat_i[28]
rlabel metal2 251384 239106 251384 239106 0 wbs_dat_i[29]
rlabel metal2 39928 110726 39928 110726 0 wbs_dat_i[2]
rlabel metal2 252280 239274 252280 239274 0 wbs_dat_i[30]
rlabel metal2 209384 15806 209384 15806 0 wbs_dat_i[31]
rlabel metal2 47544 2366 47544 2366 0 wbs_dat_i[3]
rlabel metal4 55160 4093 55160 4093 0 wbs_dat_i[4]
rlabel metal2 60872 2702 60872 2702 0 wbs_dat_i[5]
rlabel metal2 66584 2590 66584 2590 0 wbs_dat_i[6]
rlabel metal2 72296 2478 72296 2478 0 wbs_dat_i[7]
rlabel metal2 78008 24262 78008 24262 0 wbs_dat_i[8]
rlabel metal2 233464 238490 233464 238490 0 wbs_dat_i[9]
rlabel metal2 26824 2310 26824 2310 0 wbs_dat_o[0]
rlabel metal2 91336 20902 91336 20902 0 wbs_dat_o[10]
rlabel metal2 97272 2646 97272 2646 0 wbs_dat_o[11]
rlabel metal2 102984 2310 102984 2310 0 wbs_dat_o[12]
rlabel metal2 108472 20958 108472 20958 0 wbs_dat_o[13]
rlabel metal2 114296 21686 114296 21686 0 wbs_dat_o[14]
rlabel metal2 119896 21742 119896 21742 0 wbs_dat_o[15]
rlabel metal2 125608 23366 125608 23366 0 wbs_dat_o[16]
rlabel metal4 337176 143317 337176 143317 0 wbs_dat_o[17]
rlabel metal4 288344 122007 288344 122007 0 wbs_dat_o[18]
rlabel metal2 142856 21798 142856 21798 0 wbs_dat_o[19]
rlabel metal3 186760 232680 186760 232680 0 wbs_dat_o[1]
rlabel metal2 148680 1918 148680 1918 0 wbs_dat_o[20]
rlabel metal4 283080 139657 283080 139657 0 wbs_dat_o[21]
rlabel metal4 289800 122823 289800 122823 0 wbs_dat_o[22]
rlabel metal2 165816 2590 165816 2590 0 wbs_dat_o[23]
rlabel metal2 171528 2534 171528 2534 0 wbs_dat_o[24]
rlabel metal2 177016 21854 177016 21854 0 wbs_dat_o[25]
rlabel metal2 182728 19166 182728 19166 0 wbs_dat_o[26]
rlabel metal2 188440 19222 188440 19222 0 wbs_dat_o[27]
rlabel metal2 194376 2646 194376 2646 0 wbs_dat_o[28]
rlabel metal3 269752 46536 269752 46536 0 wbs_dat_o[29]
rlabel metal3 41440 4200 41440 4200 0 wbs_dat_o[2]
rlabel metal2 284760 121352 284760 121352 0 wbs_dat_o[30]
rlabel metal2 211512 2254 211512 2254 0 wbs_dat_o[31]
rlabel metal2 49448 2310 49448 2310 0 wbs_dat_o[3]
rlabel metal4 57176 4183 57176 4183 0 wbs_dat_o[4]
rlabel metal4 336952 143835 336952 143835 0 wbs_dat_o[5]
rlabel metal2 68488 21630 68488 21630 0 wbs_dat_o[6]
rlabel metal2 74424 2254 74424 2254 0 wbs_dat_o[7]
rlabel metal3 344008 238728 344008 238728 0 wbs_dat_o[8]
rlabel metal2 338632 241528 338632 241528 0 wbs_dat_o[9]
rlabel metal2 18984 114870 18984 114870 0 wbs_stb_i
rlabel metal2 21112 2310 21112 2310 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
