magic
tech gf180mcuD
magscale 1 5
timestamp 1702305931
<< obsm1 >>
rect 672 1538 109312 113385
<< metal2 >>
rect 2912 114600 2968 115000
rect 6160 114600 6216 115000
rect 9408 114600 9464 115000
rect 12656 114600 12712 115000
rect 15904 114600 15960 115000
rect 19152 114600 19208 115000
rect 22400 114600 22456 115000
rect 25648 114600 25704 115000
rect 28896 114600 28952 115000
rect 32144 114600 32200 115000
rect 35392 114600 35448 115000
rect 38640 114600 38696 115000
rect 41888 114600 41944 115000
rect 45136 114600 45192 115000
rect 48384 114600 48440 115000
rect 51632 114600 51688 115000
rect 54880 114600 54936 115000
rect 58128 114600 58184 115000
rect 61376 114600 61432 115000
rect 64624 114600 64680 115000
rect 67872 114600 67928 115000
rect 71120 114600 71176 115000
rect 74368 114600 74424 115000
rect 77616 114600 77672 115000
rect 80864 114600 80920 115000
rect 84112 114600 84168 115000
rect 87360 114600 87416 115000
rect 90608 114600 90664 115000
rect 93856 114600 93912 115000
rect 97104 114600 97160 115000
rect 100352 114600 100408 115000
rect 103600 114600 103656 115000
rect 106848 114600 106904 115000
rect 2912 0 2968 400
rect 6160 0 6216 400
rect 9408 0 9464 400
rect 12656 0 12712 400
rect 15904 0 15960 400
rect 19152 0 19208 400
rect 22400 0 22456 400
rect 25648 0 25704 400
rect 28896 0 28952 400
rect 32144 0 32200 400
rect 35392 0 35448 400
rect 38640 0 38696 400
rect 41888 0 41944 400
rect 45136 0 45192 400
rect 48384 0 48440 400
rect 51632 0 51688 400
rect 54880 0 54936 400
rect 58128 0 58184 400
rect 61376 0 61432 400
rect 64624 0 64680 400
rect 67872 0 67928 400
rect 71120 0 71176 400
rect 74368 0 74424 400
rect 77616 0 77672 400
rect 80864 0 80920 400
rect 84112 0 84168 400
rect 87360 0 87416 400
rect 90608 0 90664 400
rect 93856 0 93912 400
rect 97104 0 97160 400
rect 100352 0 100408 400
rect 103600 0 103656 400
rect 106848 0 106904 400
<< obsm2 >>
rect 462 114570 2882 114674
rect 2998 114570 6130 114674
rect 6246 114570 9378 114674
rect 9494 114570 12626 114674
rect 12742 114570 15874 114674
rect 15990 114570 19122 114674
rect 19238 114570 22370 114674
rect 22486 114570 25618 114674
rect 25734 114570 28866 114674
rect 28982 114570 32114 114674
rect 32230 114570 35362 114674
rect 35478 114570 38610 114674
rect 38726 114570 41858 114674
rect 41974 114570 45106 114674
rect 45222 114570 48354 114674
rect 48470 114570 51602 114674
rect 51718 114570 54850 114674
rect 54966 114570 58098 114674
rect 58214 114570 61346 114674
rect 61462 114570 64594 114674
rect 64710 114570 67842 114674
rect 67958 114570 71090 114674
rect 71206 114570 74338 114674
rect 74454 114570 77586 114674
rect 77702 114570 80834 114674
rect 80950 114570 84082 114674
rect 84198 114570 87330 114674
rect 87446 114570 90578 114674
rect 90694 114570 93826 114674
rect 93942 114570 97074 114674
rect 97190 114570 100322 114674
rect 100438 114570 103570 114674
rect 103686 114570 106818 114674
rect 106934 114570 109242 114674
rect 462 430 109242 114570
rect 462 289 2882 430
rect 2998 289 6130 430
rect 6246 289 9378 430
rect 9494 289 12626 430
rect 12742 289 15874 430
rect 15990 289 19122 430
rect 19238 289 22370 430
rect 22486 289 25618 430
rect 25734 289 28866 430
rect 28982 289 32114 430
rect 32230 289 35362 430
rect 35478 289 38610 430
rect 38726 289 41858 430
rect 41974 289 45106 430
rect 45222 289 48354 430
rect 48470 289 51602 430
rect 51718 289 54850 430
rect 54966 289 58098 430
rect 58214 289 61346 430
rect 61462 289 64594 430
rect 64710 289 67842 430
rect 67958 289 71090 430
rect 71206 289 74338 430
rect 74454 289 77586 430
rect 77702 289 80834 430
rect 80950 289 84082 430
rect 84198 289 87330 430
rect 87446 289 90578 430
rect 90694 289 93826 430
rect 93942 289 97074 430
rect 97190 289 100322 430
rect 100438 289 103570 430
rect 103686 289 106818 430
rect 106934 289 109242 430
<< metal3 >>
rect 0 111888 400 111944
rect 0 108864 400 108920
rect 0 105840 400 105896
rect 0 102816 400 102872
rect 0 99792 400 99848
rect 0 96768 400 96824
rect 0 93744 400 93800
rect 0 90720 400 90776
rect 0 87696 400 87752
rect 0 84672 400 84728
rect 0 81648 400 81704
rect 0 78624 400 78680
rect 0 75600 400 75656
rect 0 72576 400 72632
rect 0 69552 400 69608
rect 0 66528 400 66584
rect 0 63504 400 63560
rect 0 60480 400 60536
rect 0 57456 400 57512
rect 0 54432 400 54488
rect 0 51408 400 51464
rect 0 48384 400 48440
rect 0 45360 400 45416
rect 0 42336 400 42392
rect 0 39312 400 39368
rect 0 36288 400 36344
rect 0 33264 400 33320
rect 0 30240 400 30296
rect 0 27216 400 27272
rect 0 24192 400 24248
rect 0 21168 400 21224
rect 0 18144 400 18200
rect 0 15120 400 15176
rect 0 12096 400 12152
rect 0 9072 400 9128
rect 0 6048 400 6104
rect 0 3024 400 3080
<< obsm3 >>
rect 400 111974 109191 113554
rect 430 111858 109191 111974
rect 400 108950 109191 111858
rect 430 108834 109191 108950
rect 400 105926 109191 108834
rect 430 105810 109191 105926
rect 400 102902 109191 105810
rect 430 102786 109191 102902
rect 400 99878 109191 102786
rect 430 99762 109191 99878
rect 400 96854 109191 99762
rect 430 96738 109191 96854
rect 400 93830 109191 96738
rect 430 93714 109191 93830
rect 400 90806 109191 93714
rect 430 90690 109191 90806
rect 400 87782 109191 90690
rect 430 87666 109191 87782
rect 400 84758 109191 87666
rect 430 84642 109191 84758
rect 400 81734 109191 84642
rect 430 81618 109191 81734
rect 400 78710 109191 81618
rect 430 78594 109191 78710
rect 400 75686 109191 78594
rect 430 75570 109191 75686
rect 400 72662 109191 75570
rect 430 72546 109191 72662
rect 400 69638 109191 72546
rect 430 69522 109191 69638
rect 400 66614 109191 69522
rect 430 66498 109191 66614
rect 400 63590 109191 66498
rect 430 63474 109191 63590
rect 400 60566 109191 63474
rect 430 60450 109191 60566
rect 400 57542 109191 60450
rect 430 57426 109191 57542
rect 400 54518 109191 57426
rect 430 54402 109191 54518
rect 400 51494 109191 54402
rect 430 51378 109191 51494
rect 400 48470 109191 51378
rect 430 48354 109191 48470
rect 400 45446 109191 48354
rect 430 45330 109191 45446
rect 400 42422 109191 45330
rect 430 42306 109191 42422
rect 400 39398 109191 42306
rect 430 39282 109191 39398
rect 400 36374 109191 39282
rect 430 36258 109191 36374
rect 400 33350 109191 36258
rect 430 33234 109191 33350
rect 400 30326 109191 33234
rect 430 30210 109191 30326
rect 400 27302 109191 30210
rect 430 27186 109191 27302
rect 400 24278 109191 27186
rect 430 24162 109191 24278
rect 400 21254 109191 24162
rect 430 21138 109191 21254
rect 400 18230 109191 21138
rect 430 18114 109191 18230
rect 400 15206 109191 18114
rect 430 15090 109191 15206
rect 400 12182 109191 15090
rect 430 12066 109191 12182
rect 400 9158 109191 12066
rect 430 9042 109191 9158
rect 400 6134 109191 9042
rect 430 6018 109191 6134
rect 400 3110 109191 6018
rect 430 2994 109191 3110
rect 400 294 109191 2994
<< metal4 >>
rect 2224 1538 2384 113318
rect 9904 1538 10064 113318
rect 17584 1538 17744 113318
rect 25264 1538 25424 113318
rect 32944 1538 33104 113318
rect 40624 1538 40784 113318
rect 48304 1538 48464 113318
rect 55984 1538 56144 113318
rect 63664 1538 63824 113318
rect 71344 1538 71504 113318
rect 79024 1538 79184 113318
rect 86704 1538 86864 113318
rect 94384 1538 94544 113318
rect 102064 1538 102224 113318
<< obsm4 >>
rect 1134 113348 107786 113559
rect 1134 1508 2194 113348
rect 2414 1508 9874 113348
rect 10094 1508 17554 113348
rect 17774 1508 25234 113348
rect 25454 1508 32914 113348
rect 33134 1508 40594 113348
rect 40814 1508 48274 113348
rect 48494 1508 55954 113348
rect 56174 1508 63634 113348
rect 63854 1508 71314 113348
rect 71534 1508 78994 113348
rect 79214 1508 86674 113348
rect 86894 1508 94354 113348
rect 94574 1508 102034 113348
rect 102254 1508 107786 113348
rect 1134 289 107786 1508
<< labels >>
rlabel metal3 s 0 9072 400 9128 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 12096 400 12152 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 0 15120 400 15176 6 io_in[0]
port 3 nsew signal input
rlabel metal3 s 0 45360 400 45416 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 0 48384 400 48440 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 0 51408 400 51464 6 io_in[12]
port 6 nsew signal input
rlabel metal3 s 0 54432 400 54488 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 0 57456 400 57512 6 io_in[14]
port 8 nsew signal input
rlabel metal3 s 0 60480 400 60536 6 io_in[15]
port 9 nsew signal input
rlabel metal3 s 0 63504 400 63560 6 io_in[16]
port 10 nsew signal input
rlabel metal3 s 0 66528 400 66584 6 io_in[17]
port 11 nsew signal input
rlabel metal3 s 0 69552 400 69608 6 io_in[18]
port 12 nsew signal input
rlabel metal3 s 0 72576 400 72632 6 io_in[19]
port 13 nsew signal input
rlabel metal3 s 0 18144 400 18200 6 io_in[1]
port 14 nsew signal input
rlabel metal3 s 0 75600 400 75656 6 io_in[20]
port 15 nsew signal input
rlabel metal3 s 0 78624 400 78680 6 io_in[21]
port 16 nsew signal input
rlabel metal3 s 0 81648 400 81704 6 io_in[22]
port 17 nsew signal input
rlabel metal3 s 0 84672 400 84728 6 io_in[23]
port 18 nsew signal input
rlabel metal3 s 0 87696 400 87752 6 io_in[24]
port 19 nsew signal input
rlabel metal3 s 0 90720 400 90776 6 io_in[25]
port 20 nsew signal input
rlabel metal3 s 0 93744 400 93800 6 io_in[26]
port 21 nsew signal input
rlabel metal3 s 0 96768 400 96824 6 io_in[27]
port 22 nsew signal input
rlabel metal3 s 0 99792 400 99848 6 io_in[28]
port 23 nsew signal input
rlabel metal3 s 0 102816 400 102872 6 io_in[29]
port 24 nsew signal input
rlabel metal3 s 0 21168 400 21224 6 io_in[2]
port 25 nsew signal input
rlabel metal3 s 0 105840 400 105896 6 io_in[30]
port 26 nsew signal input
rlabel metal3 s 0 108864 400 108920 6 io_in[31]
port 27 nsew signal input
rlabel metal3 s 0 111888 400 111944 6 io_in[32]
port 28 nsew signal input
rlabel metal3 s 0 24192 400 24248 6 io_in[3]
port 29 nsew signal input
rlabel metal3 s 0 27216 400 27272 6 io_in[4]
port 30 nsew signal input
rlabel metal3 s 0 30240 400 30296 6 io_in[5]
port 31 nsew signal input
rlabel metal3 s 0 33264 400 33320 6 io_in[6]
port 32 nsew signal input
rlabel metal3 s 0 36288 400 36344 6 io_in[7]
port 33 nsew signal input
rlabel metal3 s 0 39312 400 39368 6 io_in[8]
port 34 nsew signal input
rlabel metal3 s 0 42336 400 42392 6 io_in[9]
port 35 nsew signal input
rlabel metal2 s 2912 114600 2968 115000 6 io_oeb[0]
port 36 nsew signal output
rlabel metal2 s 35392 114600 35448 115000 6 io_oeb[10]
port 37 nsew signal output
rlabel metal2 s 38640 114600 38696 115000 6 io_oeb[11]
port 38 nsew signal output
rlabel metal2 s 41888 114600 41944 115000 6 io_oeb[12]
port 39 nsew signal output
rlabel metal2 s 45136 114600 45192 115000 6 io_oeb[13]
port 40 nsew signal output
rlabel metal2 s 48384 114600 48440 115000 6 io_oeb[14]
port 41 nsew signal output
rlabel metal2 s 51632 114600 51688 115000 6 io_oeb[15]
port 42 nsew signal output
rlabel metal2 s 54880 114600 54936 115000 6 io_oeb[16]
port 43 nsew signal output
rlabel metal2 s 58128 114600 58184 115000 6 io_oeb[17]
port 44 nsew signal output
rlabel metal2 s 61376 114600 61432 115000 6 io_oeb[18]
port 45 nsew signal output
rlabel metal2 s 64624 114600 64680 115000 6 io_oeb[19]
port 46 nsew signal output
rlabel metal2 s 6160 114600 6216 115000 6 io_oeb[1]
port 47 nsew signal output
rlabel metal2 s 67872 114600 67928 115000 6 io_oeb[20]
port 48 nsew signal output
rlabel metal2 s 71120 114600 71176 115000 6 io_oeb[21]
port 49 nsew signal output
rlabel metal2 s 74368 114600 74424 115000 6 io_oeb[22]
port 50 nsew signal output
rlabel metal2 s 77616 114600 77672 115000 6 io_oeb[23]
port 51 nsew signal output
rlabel metal2 s 80864 114600 80920 115000 6 io_oeb[24]
port 52 nsew signal output
rlabel metal2 s 84112 114600 84168 115000 6 io_oeb[25]
port 53 nsew signal output
rlabel metal2 s 87360 114600 87416 115000 6 io_oeb[26]
port 54 nsew signal output
rlabel metal2 s 90608 114600 90664 115000 6 io_oeb[27]
port 55 nsew signal output
rlabel metal2 s 93856 114600 93912 115000 6 io_oeb[28]
port 56 nsew signal output
rlabel metal2 s 97104 114600 97160 115000 6 io_oeb[29]
port 57 nsew signal output
rlabel metal2 s 9408 114600 9464 115000 6 io_oeb[2]
port 58 nsew signal output
rlabel metal2 s 100352 114600 100408 115000 6 io_oeb[30]
port 59 nsew signal output
rlabel metal2 s 103600 114600 103656 115000 6 io_oeb[31]
port 60 nsew signal output
rlabel metal2 s 106848 114600 106904 115000 6 io_oeb[32]
port 61 nsew signal output
rlabel metal2 s 12656 114600 12712 115000 6 io_oeb[3]
port 62 nsew signal output
rlabel metal2 s 15904 114600 15960 115000 6 io_oeb[4]
port 63 nsew signal output
rlabel metal2 s 19152 114600 19208 115000 6 io_oeb[5]
port 64 nsew signal output
rlabel metal2 s 22400 114600 22456 115000 6 io_oeb[6]
port 65 nsew signal output
rlabel metal2 s 25648 114600 25704 115000 6 io_oeb[7]
port 66 nsew signal output
rlabel metal2 s 28896 114600 28952 115000 6 io_oeb[8]
port 67 nsew signal output
rlabel metal2 s 32144 114600 32200 115000 6 io_oeb[9]
port 68 nsew signal output
rlabel metal2 s 2912 0 2968 400 6 io_out[0]
port 69 nsew signal output
rlabel metal2 s 35392 0 35448 400 6 io_out[10]
port 70 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 io_out[11]
port 71 nsew signal output
rlabel metal2 s 41888 0 41944 400 6 io_out[12]
port 72 nsew signal output
rlabel metal2 s 45136 0 45192 400 6 io_out[13]
port 73 nsew signal output
rlabel metal2 s 48384 0 48440 400 6 io_out[14]
port 74 nsew signal output
rlabel metal2 s 51632 0 51688 400 6 io_out[15]
port 75 nsew signal output
rlabel metal2 s 54880 0 54936 400 6 io_out[16]
port 76 nsew signal output
rlabel metal2 s 58128 0 58184 400 6 io_out[17]
port 77 nsew signal output
rlabel metal2 s 61376 0 61432 400 6 io_out[18]
port 78 nsew signal output
rlabel metal2 s 64624 0 64680 400 6 io_out[19]
port 79 nsew signal output
rlabel metal2 s 6160 0 6216 400 6 io_out[1]
port 80 nsew signal output
rlabel metal2 s 67872 0 67928 400 6 io_out[20]
port 81 nsew signal output
rlabel metal2 s 71120 0 71176 400 6 io_out[21]
port 82 nsew signal output
rlabel metal2 s 74368 0 74424 400 6 io_out[22]
port 83 nsew signal output
rlabel metal2 s 77616 0 77672 400 6 io_out[23]
port 84 nsew signal output
rlabel metal2 s 80864 0 80920 400 6 io_out[24]
port 85 nsew signal output
rlabel metal2 s 84112 0 84168 400 6 io_out[25]
port 86 nsew signal output
rlabel metal2 s 87360 0 87416 400 6 io_out[26]
port 87 nsew signal output
rlabel metal2 s 90608 0 90664 400 6 io_out[27]
port 88 nsew signal output
rlabel metal2 s 93856 0 93912 400 6 io_out[28]
port 89 nsew signal output
rlabel metal2 s 97104 0 97160 400 6 io_out[29]
port 90 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 io_out[2]
port 91 nsew signal output
rlabel metal2 s 100352 0 100408 400 6 io_out[30]
port 92 nsew signal output
rlabel metal2 s 103600 0 103656 400 6 io_out[31]
port 93 nsew signal output
rlabel metal2 s 106848 0 106904 400 6 io_out[32]
port 94 nsew signal output
rlabel metal2 s 12656 0 12712 400 6 io_out[3]
port 95 nsew signal output
rlabel metal2 s 15904 0 15960 400 6 io_out[4]
port 96 nsew signal output
rlabel metal2 s 19152 0 19208 400 6 io_out[5]
port 97 nsew signal output
rlabel metal2 s 22400 0 22456 400 6 io_out[6]
port 98 nsew signal output
rlabel metal2 s 25648 0 25704 400 6 io_out[7]
port 99 nsew signal output
rlabel metal2 s 28896 0 28952 400 6 io_out[8]
port 100 nsew signal output
rlabel metal2 s 32144 0 32200 400 6 io_out[9]
port 101 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 rst_n
port 102 nsew signal input
rlabel metal4 s 2224 1538 2384 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal3 s 0 3024 400 3080 6 wb_clk_i
port 105 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 115000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 45147814
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_tholin_riscv/runs/23_12_11_14_09/results/signoff/wrapped_tholin_riscv.magic.gds
string GDS_START 563000
<< end >>

