module wrapped_ay8913 (rst_n,
    vdd,
    vss,
    wb_clk_i,
    custom_settings,
    io_in_1,
    io_in_2,
    io_out);
 input rst_n;
 inout vdd;
 inout vss;
 input wb_clk_i;
 input [3:0] custom_settings;
 input [7:0] io_in_1;
 input [1:0] io_in_2;
 output [27:0] io_out;

 wire net20;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net21;
 wire net38;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire \blink.LED ;
 wire \blink.counter[0] ;
 wire \blink.counter[10] ;
 wire \blink.counter[11] ;
 wire \blink.counter[12] ;
 wire \blink.counter[13] ;
 wire \blink.counter[14] ;
 wire \blink.counter[15] ;
 wire \blink.counter[16] ;
 wire \blink.counter[17] ;
 wire \blink.counter[18] ;
 wire \blink.counter[19] ;
 wire \blink.counter[1] ;
 wire \blink.counter[20] ;
 wire \blink.counter[21] ;
 wire \blink.counter[22] ;
 wire \blink.counter[23] ;
 wire \blink.counter[24] ;
 wire \blink.counter[25] ;
 wire \blink.counter[26] ;
 wire \blink.counter[27] ;
 wire \blink.counter[28] ;
 wire \blink.counter[29] ;
 wire \blink.counter[2] ;
 wire \blink.counter[30] ;
 wire \blink.counter[31] ;
 wire \blink.counter[3] ;
 wire \blink.counter[4] ;
 wire \blink.counter[5] ;
 wire \blink.counter[6] ;
 wire \blink.counter[7] ;
 wire \blink.counter[8] ;
 wire \blink.counter[9] ;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \tt_um_rejunity_ay8913.DAC_clk ;
 wire \tt_um_rejunity_ay8913.DAC_dat ;
 wire \tt_um_rejunity_ay8913.DAC_le ;
 wire \tt_um_rejunity_ay8913.active ;
 wire \tt_um_rejunity_ay8913.amplitude_A[0] ;
 wire \tt_um_rejunity_ay8913.amplitude_B[0] ;
 wire \tt_um_rejunity_ay8913.amplitude_C[0] ;
 wire \tt_um_rejunity_ay8913.clk_counter[0] ;
 wire \tt_um_rejunity_ay8913.clk_counter[1] ;
 wire \tt_um_rejunity_ay8913.clk_counter[2] ;
 wire \tt_um_rejunity_ay8913.clk_counter[3] ;
 wire \tt_um_rejunity_ay8913.clk_counter[4] ;
 wire \tt_um_rejunity_ay8913.clk_counter[5] ;
 wire \tt_um_rejunity_ay8913.clk_counter[6] ;
 wire \tt_um_rejunity_ay8913.envelope_A ;
 wire \tt_um_rejunity_ay8913.envelope_B ;
 wire \tt_um_rejunity_ay8913.envelope_C ;
 wire \tt_um_rejunity_ay8913.envelope_alternate ;
 wire \tt_um_rejunity_ay8913.envelope_attack ;
 wire \tt_um_rejunity_ay8913.envelope_continue ;
 wire \tt_um_rejunity_ay8913.envelope_generator.envelope_counter[0] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.envelope_counter[1] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.envelope_counter[2] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.envelope_counter[3] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.hold ;
 wire \tt_um_rejunity_ay8913.envelope_generator.invert_output ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[0] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[10] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[11] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[12] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[13] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[14] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[15] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[1] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[2] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[3] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[4] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[5] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[6] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[7] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[8] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.period[9] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0 ;
 wire \tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal ;
 wire \tt_um_rejunity_ay8913.envelope_generator.stop ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[0] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[10] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[11] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[12] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[13] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[14] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[15] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[1] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[2] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[3] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[4] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[5] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[6] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[7] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[8] ;
 wire \tt_um_rejunity_ay8913.envelope_generator.tone.counter[9] ;
 wire \tt_um_rejunity_ay8913.latched_register[0] ;
 wire \tt_um_rejunity_ay8913.latched_register[1] ;
 wire \tt_um_rejunity_ay8913.latched_register[2] ;
 wire \tt_um_rejunity_ay8913.latched_register[3] ;
 wire \tt_um_rejunity_ay8913.noise_disable_A ;
 wire \tt_um_rejunity_ay8913.noise_disable_B ;
 wire \tt_um_rejunity_ay8913.noise_disable_C ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[0] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[10] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[11] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[12] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[13] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[14] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[15] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[16] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[1] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[2] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[3] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[4] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[5] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[6] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[7] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[8] ;
 wire \tt_um_rejunity_ay8913.noise_generator.lfsr[9] ;
 wire \tt_um_rejunity_ay8913.noise_generator.period[0] ;
 wire \tt_um_rejunity_ay8913.noise_generator.period[1] ;
 wire \tt_um_rejunity_ay8913.noise_generator.period[2] ;
 wire \tt_um_rejunity_ay8913.noise_generator.period[3] ;
 wire \tt_um_rejunity_ay8913.noise_generator.period[4] ;
 wire \tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0 ;
 wire \tt_um_rejunity_ay8913.noise_generator.signal_edge.signal ;
 wire \tt_um_rejunity_ay8913.noise_generator.tone.counter[0] ;
 wire \tt_um_rejunity_ay8913.noise_generator.tone.counter[1] ;
 wire \tt_um_rejunity_ay8913.noise_generator.tone.counter[2] ;
 wire \tt_um_rejunity_ay8913.noise_generator.tone.counter[3] ;
 wire \tt_um_rejunity_ay8913.noise_generator.tone.counter[4] ;
 wire \tt_um_rejunity_ay8913.pwm_A.accumulator[2] ;
 wire \tt_um_rejunity_ay8913.pwm_A.accumulator[3] ;
 wire \tt_um_rejunity_ay8913.pwm_A.accumulator[4] ;
 wire \tt_um_rejunity_ay8913.pwm_A.accumulator[5] ;
 wire \tt_um_rejunity_ay8913.pwm_A.accumulator[6] ;
 wire \tt_um_rejunity_ay8913.pwm_A.accumulator[7] ;
 wire \tt_um_rejunity_ay8913.pwm_A.accumulator[8] ;
 wire \tt_um_rejunity_ay8913.pwm_A.accumulator[9] ;
 wire \tt_um_rejunity_ay8913.pwm_B.accumulator[2] ;
 wire \tt_um_rejunity_ay8913.pwm_B.accumulator[3] ;
 wire \tt_um_rejunity_ay8913.pwm_B.accumulator[4] ;
 wire \tt_um_rejunity_ay8913.pwm_B.accumulator[5] ;
 wire \tt_um_rejunity_ay8913.pwm_B.accumulator[6] ;
 wire \tt_um_rejunity_ay8913.pwm_B.accumulator[7] ;
 wire \tt_um_rejunity_ay8913.pwm_B.accumulator[8] ;
 wire \tt_um_rejunity_ay8913.pwm_B.accumulator[9] ;
 wire \tt_um_rejunity_ay8913.pwm_C.accumulator[2] ;
 wire \tt_um_rejunity_ay8913.pwm_C.accumulator[3] ;
 wire \tt_um_rejunity_ay8913.pwm_C.accumulator[4] ;
 wire \tt_um_rejunity_ay8913.pwm_C.accumulator[5] ;
 wire \tt_um_rejunity_ay8913.pwm_C.accumulator[6] ;
 wire \tt_um_rejunity_ay8913.pwm_C.accumulator[7] ;
 wire \tt_um_rejunity_ay8913.pwm_C.accumulator[8] ;
 wire \tt_um_rejunity_ay8913.pwm_C.accumulator[9] ;
 wire \tt_um_rejunity_ay8913.pwm_master.accumulator[10] ;
 wire \tt_um_rejunity_ay8913.pwm_master.accumulator[2] ;
 wire \tt_um_rejunity_ay8913.pwm_master.accumulator[3] ;
 wire \tt_um_rejunity_ay8913.pwm_master.accumulator[4] ;
 wire \tt_um_rejunity_ay8913.pwm_master.accumulator[5] ;
 wire \tt_um_rejunity_ay8913.pwm_master.accumulator[6] ;
 wire \tt_um_rejunity_ay8913.pwm_master.accumulator[7] ;
 wire \tt_um_rejunity_ay8913.pwm_master.accumulator[8] ;
 wire \tt_um_rejunity_ay8913.pwm_master.accumulator[9] ;
 wire \tt_um_rejunity_ay8913.restart_envelope ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.counter[0] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.counter[1] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.counter[2] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.counter[3] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.counter[4] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[10] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[11] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[2] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[3] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[4] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[5] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[6] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[7] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[8] ;
 wire \tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[9] ;
 wire \tt_um_rejunity_ay8913.tone_A ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[0] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[10] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[11] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[1] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[2] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[3] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[4] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[5] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[6] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[7] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[8] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.counter[9] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[0] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[10] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[11] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[1] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[2] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[3] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[4] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[5] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[6] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[7] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[8] ;
 wire \tt_um_rejunity_ay8913.tone_A_generator.period[9] ;
 wire \tt_um_rejunity_ay8913.tone_B ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[0] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[10] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[11] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[1] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[2] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[3] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[4] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[5] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[6] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[7] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[8] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.counter[9] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[0] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[10] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[11] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[1] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[2] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[3] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[4] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[5] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[6] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[7] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[8] ;
 wire \tt_um_rejunity_ay8913.tone_B_generator.period[9] ;
 wire \tt_um_rejunity_ay8913.tone_C ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[0] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[10] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[11] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[1] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[2] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[3] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[4] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[5] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[6] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[7] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[8] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.counter[9] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[0] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[10] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[11] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[1] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[2] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[3] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[4] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[5] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[6] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[7] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[8] ;
 wire \tt_um_rejunity_ay8913.tone_C_generator.period[9] ;
 wire \tt_um_rejunity_ay8913.tone_disable_A ;
 wire \tt_um_rejunity_ay8913.tone_disable_B ;
 wire \tt_um_rejunity_ay8913.tone_disable_C ;

 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1272__S (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net3));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1274__S (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net3));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1276__S (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net3));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1278__S (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net3));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1331__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0966_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1341__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0973_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1393__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0966_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1397__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0973_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1421__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0973_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1432__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0973_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1457__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0966_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1460__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1461__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1066_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1466__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net9));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1467__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net8));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1467__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net10));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1470__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1075_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1471__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net10));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1473__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1078_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1475__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1075_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1477__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1067_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1479__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[1]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1480__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1084_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1482__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[2]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1483__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1086_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1485__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[3]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1488__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net4));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1490__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1091_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1490__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1075_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1494__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1094_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1495__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1078_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1497__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1097_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1497__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1094_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1498__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1067_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1500__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1084_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1502__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1086_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1507__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1103_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1510__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1104_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1514__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net10));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1515__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1110_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1517__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1111_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1523__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1104_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1527__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1104_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1531__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1110_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1537__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1128_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1541__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1111_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1544__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1133_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1550__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1110_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1551__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1139_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1553__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net10));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1554__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1141_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1562__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1142_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1566__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1142_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1617__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1139_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1649__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1139_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1654__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1078_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1655__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1214_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1657__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1067_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1659__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1084_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1661__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1086_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1667__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1091_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1669__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net5));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1670__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1224_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1672__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net6));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1673__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1226_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1676__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1228_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1681__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1232_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1682__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1097_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1682__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1232_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1683__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1067_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1685__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1084_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1687__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1086_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1691__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1694__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1214_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1696__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1239_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1698__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[1]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1699__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1245_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1701__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[2]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1702__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1247_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1704__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[3]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1705__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1249_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1709__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1091_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1711__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1224_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1713__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1226_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1715__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1228_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1734__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1133_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1761__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1142_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1762__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0276_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1763__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0277_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1767__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1128_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1768__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1239_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1770__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1091_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1775__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1214_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1777__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1239_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1779__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1245_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1781__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1247_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1783__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1249_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1788__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0293_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1790__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1224_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1792__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1226_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1794__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1228_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1798__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1214_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1800__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1239_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1802__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1245_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1804__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1247_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1806__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1249_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1810__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0293_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1812__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1224_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1814__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1226_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1816__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1228_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1818__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1139_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1821__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0276_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1823__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1142_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1825__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1830__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0318_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1832__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1245_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1834__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1247_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1836__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1249_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1838__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0293_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1840__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net5));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1926__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net2));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1929__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net1));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1930__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0410_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1933__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net1));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1933__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net2));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1935__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0415_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1937__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0417_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1938__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1078_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1939__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0419_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1941__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0419_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1945__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0417_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1946__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0425_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1947__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0424_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1952__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0430_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1980__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0424_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1998__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0424_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2002__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0424_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2014__S (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0419_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2032__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0492_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2037__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0492_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2053__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1133_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2068__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1133_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2082__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1128_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2097__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0542_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2111__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1141_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2114__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0425_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2118__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0542_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2186__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0624_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2187__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1141_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2189__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0425_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2193__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0410_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2193__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0415_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2194__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0430_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2235__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1097_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2236__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0318_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2238__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[1]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2241__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[2]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2244__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[3]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2304__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0542_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2306__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0425_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2310__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0410_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2310__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0415_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2311__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0430_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2349__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0492_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2403__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0417_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2404__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1141_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2404__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0812_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2406__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0417_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2410__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0410_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2410__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0415_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2411__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0430_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2417__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0821_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2437__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0821_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2444__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0821_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2446__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0821_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2447__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0812_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2450__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1104_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2460__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1111_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2464__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1111_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2468__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1110_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2472__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0276_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2474__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net9));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2474__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net8));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2475__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net6));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2475__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net5));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2476__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net4));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2479__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0276_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2483__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1066_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2490__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1103_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2495__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1103_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2500__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1103_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2504__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0966_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2509__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0318_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2519__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0293_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2521__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net5));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2523__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net6));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2528__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1128_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2529__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0318_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2534__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1097_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2535__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1066_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2539__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0492_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2540__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1066_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_2_0__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_2_1__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_2_2__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_2_3__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_38_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_39_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_40_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_41_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_42_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_43_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload0_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload1_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input10_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(rst_n));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input1_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input2_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[1]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input3_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[3]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input4_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[4]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input5_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[5]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input6_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[6]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input7_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[7]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input8_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_2[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input9_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_2[1]));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_0_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_0_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_0_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_0_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_14_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_420 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_1_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_22_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_27_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_28_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_28_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_421 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_31_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_31_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_32_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_32_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_32_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_32_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_32_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_32_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_32_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_34_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_34_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_34_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_34_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_35_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_35_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_35_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_35_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_35_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_35_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_36_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_180 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_39_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_39_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_40_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_40_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_41_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_41_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_41_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_42_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_43_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_45_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_180 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_45_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_46_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_46_145 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_46_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_46_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_46_355 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_47_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_47_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_47_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_47_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_48_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_48_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_48_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_71 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_49_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_49_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_49_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_50_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_50_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_50_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_50_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_50_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_51_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_51_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_51_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_52_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_52_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_52_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_52_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_52_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_52_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_53_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_53_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_53_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_53_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_53_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_53_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_53_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_53_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_54_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_54_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_54_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_54_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_54_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_54_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_54_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_55_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_55_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_55_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_55_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_55_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_55_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_55_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_55_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_55_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_55_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_55_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_55_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_55_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_55_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_55_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_55_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_55_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_55_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_55_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_55_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_55_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_55_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_56_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_56_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_56_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_56_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_56_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_56_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_56_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_56_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_56_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_56_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_56_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_56_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_56_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_56_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_56_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_56_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_56_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_56_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_56_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_56_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_56_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_320 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Left_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Left_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Left_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Left_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Left_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Left_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Left_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Left_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Left_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Left_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Left_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Left_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Left_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Left_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_22_Left_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_23_Left_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_24_Left_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_25_Left_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_26_Left_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_27_Left_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_28_Left_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_29_Left_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Left_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_30_Left_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_31_Left_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_32_Left_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_33_Left_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_34_Left_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_35_Left_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_36_Left_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_37_Left_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_38_Left_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_39_Left_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Left_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_40_Left_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_41_Left_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_42_Left_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_43_Left_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_44_Left_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_45_Left_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_45_Right_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_46_Left_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_46_Right_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_47_Left_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_47_Right_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_48_Left_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_48_Right_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_49_Left_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_49_Right_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Left_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_50_Left_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_50_Right_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_51_Left_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_51_Right_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_52_Left_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_52_Right_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_53_Left_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_53_Right_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_54_Left_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_54_Right_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_55_Left_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_55_Right_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_56_Left_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_56_Right_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Left_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Left_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Left_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Left_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Left_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_55_450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_55_451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_55_452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_55_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_55_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_55_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_56_467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1271_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.LED ),
    .Y(_0915_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _1272_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(net3),
    .B(_0915_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[9] ),
    .Y(_0916_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1273_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0916_),
    .Y(net18));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _1274_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(net3),
    .B(_0915_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[9] ),
    .Y(_0917_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1275_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0917_),
    .Y(net19));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _1276_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(net3),
    .B(_0915_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[9] ),
    .Y(_0918_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1277_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0918_),
    .Y(net11));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _1278_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(net3),
    .B(_0915_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[10] ),
    .Y(_0919_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1279_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0919_),
    .Y(net12));
 gf180mcu_as_sc_mcu7t3v3__xnor2_4 _1280_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.envelope_generator.invert_output ),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[0] ),
    .Y(_0920_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1281_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0921_),
    .B(\tt_um_rejunity_ay8913.noise_generator.lfsr[0] ),
    .A(\tt_um_rejunity_ay8913.noise_disable_C ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1282_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_disable_C ),
    .A(\tt_um_rejunity_ay8913.tone_C ),
    .Y(_0922_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1283_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.envelope_C ),
    .A(\tt_um_rejunity_ay8913.amplitude_C[0] ),
    .Y(_0923_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _1284_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0921_),
    .B(_0922_),
    .C(_0923_),
    .Y(_0924_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_4 _1285_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0925_),
    .C(_0924_),
    .B(_0920_),
    .A(\tt_um_rejunity_ay8913.envelope_C ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1286_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.envelope_B ),
    .A(\tt_um_rejunity_ay8913.amplitude_B[0] ),
    .Y(_0926_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1287_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_disable_B ),
    .A(\tt_um_rejunity_ay8913.tone_B ),
    .Y(_0927_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1288_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[0] ),
    .Y(_0928_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1289_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0929_),
    .B(_0928_),
    .A(\tt_um_rejunity_ay8913.noise_disable_B ));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _1290_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0926_),
    .B(_0927_),
    .C(_0929_),
    .Y(_0930_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_4 _1291_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0931_),
    .C(_0930_),
    .B(_0920_),
    .A(\tt_um_rejunity_ay8913.envelope_B ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1292_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.envelope_A ),
    .A(\tt_um_rejunity_ay8913.amplitude_A[0] ),
    .Y(_0932_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1293_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_disable_A ),
    .A(\tt_um_rejunity_ay8913.tone_A ),
    .Y(_0933_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1294_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0934_),
    .B(_0928_),
    .A(\tt_um_rejunity_ay8913.noise_disable_A ));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _1295_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0932_),
    .B(_0933_),
    .C(_0934_),
    .Y(_0935_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1296_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0936_),
    .C(_0935_),
    .B(_0920_),
    .A(\tt_um_rejunity_ay8913.envelope_A ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1297_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0936_),
    .A(_0931_),
    .Y(_0937_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1298_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0937_),
    .A(_0925_),
    .Y(_0938_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1299_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0938_),
    .Y(net16));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1300_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0939_),
    .A(_0925_),
    .B(_0931_),
    .C(_0936_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1301_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0939_),
    .Y(net17));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1302_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[0] ),
    .Y(_0940_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _1303_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[22] ),
    .B(\blink.counter[21] ),
    .C(\blink.counter[20] ),
    .Y(_0941_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1304_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0942_),
    .B(_0941_),
    .A(\blink.counter[19] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1305_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0943_),
    .A(\blink.counter[18] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1306_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0944_),
    .A(\blink.counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1307_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0945_),
    .A(\blink.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1308_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0946_),
    .A(\blink.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1309_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0947_),
    .A(\blink.counter[12] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1310_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0947_),
    .A(_0944_),
    .B(_0945_),
    .C(_0946_),
    .Y(_0948_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1311_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0949_),
    .B(\blink.counter[15] ),
    .A(\blink.counter[13] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1312_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0950_),
    .B(\blink.counter[16] ),
    .A(\blink.counter[14] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1313_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0951_),
    .A(\blink.counter[17] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1314_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0951_),
    .A(_0948_),
    .B(_0949_),
    .C(_0950_),
    .Y(_0952_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1315_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0953_),
    .B(_0952_),
    .A(_0943_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1316_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0954_),
    .B(_0953_),
    .A(_0942_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1317_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\blink.counter[30] ),
    .A(\blink.counter[28] ),
    .Y(_0955_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1318_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[26] ),
    .B(\blink.counter[29] ),
    .C(_0955_),
    .Y(_0956_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1319_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\blink.counter[25] ),
    .A(\blink.counter[23] ),
    .Y(_0957_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1320_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[24] ),
    .B(\blink.counter[27] ),
    .C(_0957_),
    .Y(_0958_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _1321_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0954_),
    .B(_0956_),
    .C(_0958_),
    .Y(_0959_),
    .D(\blink.counter[31] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1322_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0959_),
    .Y(_0960_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1323_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0960_),
    .Y(_0961_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1324_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0000_),
    .B(_0961_),
    .A(_0940_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1325_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0940_),
    .A(\blink.counter[1] ),
    .Y(_0962_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1326_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0963_),
    .B(_0940_),
    .A(\blink.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1327_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0961_),
    .B(_0962_),
    .C(_0963_),
    .Y(_0964_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1328_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0964_),
    .Y(_0001_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1329_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0959_),
    .Y(_0965_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1330_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0965_),
    .Y(_0966_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1331_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0966_),
    .Y(_0967_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1332_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0962_),
    .A(\blink.counter[2] ),
    .Y(_0968_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1333_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0002_),
    .B(_0968_),
    .A(_0967_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1334_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[1] ),
    .B(\blink.counter[0] ),
    .C(\blink.counter[3] ),
    .D(\blink.counter[2] ),
    .Y(_0969_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1335_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\blink.counter[3] ),
    .A(\blink.counter[1] ),
    .B(_0940_),
    .C(\blink.counter[2] ),
    .Y(_0970_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1336_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0971_),
    .B(_0970_),
    .A(_0969_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1337_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0003_),
    .B(_0971_),
    .A(_0967_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1338_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0972_),
    .A(\blink.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1339_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0965_),
    .Y(_0973_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1340_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0974_),
    .B(_0969_),
    .A(_0972_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1341_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0974_),
    .A(_0973_),
    .Y(_0975_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1342_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0004_),
    .C(_0975_),
    .B(_0969_),
    .A(_0972_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1343_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0974_),
    .A(\blink.counter[5] ),
    .Y(_0976_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1344_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0005_),
    .B(_0976_),
    .A(_0967_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1345_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0977_),
    .A(\blink.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1346_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0977_),
    .B(_0972_),
    .C(_0969_),
    .Y(_0978_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1347_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0979_),
    .B(_0978_),
    .A(\blink.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1348_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0978_),
    .A(\blink.counter[6] ),
    .Y(_0980_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1349_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0961_),
    .B(_0979_),
    .C(_0980_),
    .Y(_0981_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1350_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0981_),
    .Y(_0006_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1351_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0960_),
    .Y(_0982_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1352_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0980_),
    .A(\blink.counter[7] ),
    .Y(_0983_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1353_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0984_),
    .B(_0980_),
    .A(\blink.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1354_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0982_),
    .B(_0983_),
    .C(_0984_),
    .Y(_0985_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1355_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0985_),
    .Y(_0007_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1356_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0983_),
    .A(\blink.counter[8] ),
    .Y(_0986_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1357_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0008_),
    .B(_0986_),
    .A(_0967_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1358_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0983_),
    .A(\blink.counter[8] ),
    .Y(_0987_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1359_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0988_),
    .B(_0987_),
    .A(\blink.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1360_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0987_),
    .A(\blink.counter[9] ),
    .Y(_0989_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1361_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0982_),
    .B(_0988_),
    .C(_0989_),
    .Y(_0990_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1362_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0990_),
    .Y(_0009_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1363_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0991_),
    .B(_0989_),
    .A(\blink.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1364_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\blink.counter[8] ),
    .A(\blink.counter[10] ),
    .Y(_0992_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1365_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0992_),
    .A(\blink.counter[9] ),
    .Y(_0993_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1366_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0993_),
    .A(_0983_),
    .Y(_0994_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1367_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0982_),
    .B(_0991_),
    .C(_0994_),
    .Y(_0995_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1368_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0995_),
    .Y(_0010_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1369_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[7] ),
    .B(\blink.counter[6] ),
    .C(_0978_),
    .D(_0993_),
    .Y(_0996_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1370_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0996_),
    .A(_0944_),
    .Y(_0997_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1371_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0011_),
    .B(_0997_),
    .A(_0961_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1372_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0947_),
    .B(_0944_),
    .C(_0996_),
    .Y(_0998_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1373_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0998_),
    .Y(_0999_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1374_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1000_),
    .C(\blink.counter[12] ),
    .B(_0994_),
    .A(\blink.counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1375_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0982_),
    .B(_0999_),
    .C(_1000_),
    .Y(_1001_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1376_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1001_),
    .Y(_0012_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1377_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0960_),
    .Y(_1002_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1378_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1003_),
    .B(_0999_),
    .A(\blink.counter[13] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1379_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0999_),
    .A(\blink.counter[13] ),
    .Y(_1004_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1380_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1002_),
    .B(_1003_),
    .C(_1004_),
    .Y(_1005_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1381_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1005_),
    .Y(_0013_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1382_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1006_),
    .B(_1004_),
    .A(\blink.counter[14] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1383_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\blink.counter[14] ),
    .A(\blink.counter[13] ),
    .Y(_1007_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1384_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1007_),
    .A(_0999_),
    .Y(_1008_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1385_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1002_),
    .B(_1006_),
    .C(_1008_),
    .Y(_1009_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1386_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1009_),
    .Y(_0014_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1387_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1010_),
    .B(_1008_),
    .A(\blink.counter[15] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1388_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1008_),
    .A(\blink.counter[15] ),
    .Y(_1011_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1389_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1002_),
    .B(_1010_),
    .C(_1011_),
    .Y(_1012_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1390_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1012_),
    .Y(_0015_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1391_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[15] ),
    .B(\blink.counter[16] ),
    .C(_0998_),
    .D(_1007_),
    .Y(_1013_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1392_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1014_),
    .B(_1011_),
    .A(\blink.counter[16] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1393_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1015_),
    .B(_1014_),
    .A(_0966_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1394_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1015_),
    .A(_1013_),
    .Y(_1016_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1395_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1016_),
    .Y(_0016_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1396_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1017_),
    .B(_1013_),
    .A(_0951_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1397_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1017_),
    .A(_0973_),
    .Y(_1018_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1398_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0017_),
    .C(_1018_),
    .B(_1013_),
    .A(_0951_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1399_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1019_),
    .B(_1017_),
    .A(\blink.counter[18] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1400_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0943_),
    .B(_0951_),
    .C(_1013_),
    .Y(_1020_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1401_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1020_),
    .Y(_1021_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1402_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1002_),
    .B(_1019_),
    .C(_1021_),
    .Y(_1022_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1403_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1022_),
    .Y(_0018_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1404_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0960_),
    .Y(_1023_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1405_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1024_),
    .B(_1021_),
    .A(\blink.counter[19] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1406_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1021_),
    .A(\blink.counter[19] ),
    .Y(_1025_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1407_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1023_),
    .B(_1024_),
    .C(_1025_),
    .Y(_1026_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1408_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1026_),
    .Y(_0019_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1409_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1027_),
    .B(_1025_),
    .A(\blink.counter[20] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1410_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1025_),
    .A(\blink.counter[20] ),
    .Y(_1028_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1411_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1023_),
    .B(_1027_),
    .C(_1028_),
    .Y(_1029_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1412_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1029_),
    .Y(_0020_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1413_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1030_),
    .B(_1028_),
    .A(\blink.counter[21] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1414_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1028_),
    .A(\blink.counter[21] ),
    .Y(_1031_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1415_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1023_),
    .B(_1030_),
    .C(_1031_),
    .Y(_1032_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1416_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1032_),
    .Y(_0021_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1417_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1033_),
    .B(_1031_),
    .A(\blink.counter[22] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1418_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1020_),
    .A(_0942_),
    .Y(_1034_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1419_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1023_),
    .B(_1033_),
    .C(_1034_),
    .Y(_1035_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1420_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1035_),
    .Y(_0022_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1421_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0973_),
    .Y(_1036_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1422_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1037_),
    .B(_1034_),
    .A(\blink.counter[23] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1423_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1034_),
    .A(\blink.counter[23] ),
    .Y(_1038_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1424_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1036_),
    .B(_1037_),
    .C(_1038_),
    .Y(_1039_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1425_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1039_),
    .Y(_0023_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1426_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1040_),
    .B(_1038_),
    .A(\blink.counter[24] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1427_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1038_),
    .A(\blink.counter[24] ),
    .Y(_1041_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1428_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1036_),
    .B(_1040_),
    .C(_1041_),
    .Y(_1042_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1429_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1042_),
    .Y(_0024_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1430_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1043_),
    .A(\blink.counter[25] ));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1431_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[23] ),
    .B(\blink.counter[24] ),
    .C(_0942_),
    .D(_1021_),
    .Y(_1044_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1432_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1045_),
    .A(_1043_),
    .B(_1044_),
    .C(_0973_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1433_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0025_),
    .C(_1045_),
    .B(_1041_),
    .A(\blink.counter[25] ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1434_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1046_),
    .C(\blink.counter[26] ),
    .B(_1041_),
    .A(\blink.counter[25] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1435_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1047_),
    .A(\blink.counter[26] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1436_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1043_),
    .B(_1047_),
    .C(_1044_),
    .Y(_1048_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1437_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1048_),
    .Y(_1049_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1438_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1036_),
    .B(_1046_),
    .C(_1049_),
    .Y(_1050_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1439_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1050_),
    .Y(_0026_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1440_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[27] ),
    .Y(_1051_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1441_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1052_),
    .B(_1049_),
    .A(_1051_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1442_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1048_),
    .A(_1051_),
    .Y(_1053_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1443_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1036_),
    .B(_1052_),
    .C(_1053_),
    .Y(_1054_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1444_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1054_),
    .Y(_0027_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1445_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[28] ),
    .Y(_1055_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1446_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1056_),
    .B(_1053_),
    .A(_1055_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1447_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0965_),
    .A(_1051_),
    .B(_1055_),
    .C(_1049_),
    .Y(_1057_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1448_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0028_),
    .B(_1057_),
    .A(_1056_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1449_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\blink.counter[29] ),
    .Y(_1058_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1450_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1059_),
    .A(_1058_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _1451_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1051_),
    .B(\blink.counter[28] ),
    .C(_1049_),
    .Y(_1060_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1452_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0965_),
    .A(_1058_),
    .B(_1055_),
    .C(_1053_),
    .Y(_1061_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1453_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0029_),
    .C(_1061_),
    .B(_1060_),
    .A(_1059_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _1454_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1058_),
    .B(_1055_),
    .C(_1053_),
    .Y(_1062_),
    .D(\blink.counter[30] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1455_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1063_),
    .B(\blink.counter[30] ),
    .A(_1058_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1456_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1064_),
    .B(_1063_),
    .A(_1060_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1457_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0966_),
    .B(_1062_),
    .C(_1064_),
    .Y(_1065_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1458_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1065_),
    .Y(_0030_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1459_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0031_),
    .B(_1064_),
    .A(\blink.counter[31] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1460_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[0]),
    .Y(_1066_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1461_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1066_),
    .Y(_1067_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1462_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.latched_register[1] ),
    .Y(_1068_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1463_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.latched_register[0] ),
    .Y(_1069_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1464_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1070_),
    .B(_1069_),
    .A(_1068_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1465_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1071_),
    .A(\tt_um_rejunity_ay8913.latched_register[2] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1466_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1072_),
    .A(net9));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1467_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.active ),
    .B(_1072_),
    .C(net8),
    .D(net10),
    .Y(_1073_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1468_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.latched_register[3] ),
    .B(_1071_),
    .C(_1073_),
    .Y(_1074_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1469_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1074_),
    .A(_1070_),
    .Y(_1075_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1470_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1075_),
    .Y(_1076_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1471_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1077_),
    .A(net10));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1472_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1077_),
    .Y(_1078_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1473_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1078_),
    .Y(_1079_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1474_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1079_),
    .Y(_1080_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1475_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1081_),
    .B(_1075_),
    .A(_1080_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1476_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1081_),
    .Y(_1082_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1477_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1067_),
    .B(_1076_),
    .C(_1082_),
    .D(\tt_um_rejunity_ay8913.noise_generator.period[0] ),
    .Y(_1083_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1478_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1083_),
    .Y(_0032_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1479_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[1]),
    .Y(_1084_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1480_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1084_),
    .B(_1076_),
    .C(_1082_),
    .D(\tt_um_rejunity_ay8913.noise_generator.period[1] ),
    .Y(_1085_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1481_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1085_),
    .Y(_0033_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1482_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[2]),
    .Y(_1086_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1483_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1086_),
    .B(_1076_),
    .C(_1082_),
    .D(\tt_um_rejunity_ay8913.noise_generator.period[2] ),
    .Y(_1087_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1484_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1087_),
    .Y(_0034_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1485_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[3]),
    .Y(_1088_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1486_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1088_),
    .B(_1076_),
    .C(_1082_),
    .D(\tt_um_rejunity_ay8913.noise_generator.period[3] ),
    .Y(_1089_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1487_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1089_),
    .Y(_0035_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1488_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net4),
    .Y(_1090_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1489_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1090_),
    .Y(_1091_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1490_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1091_),
    .B(_1075_),
    .C(_1081_),
    .D(\tt_um_rejunity_ay8913.noise_generator.period[4] ),
    .Y(_1092_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1491_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1092_),
    .Y(_0036_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1492_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1093_),
    .B(_1068_),
    .A(_1069_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1493_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1093_),
    .A(_1074_),
    .Y(_1094_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1494_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1094_),
    .Y(_1095_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1495_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1078_),
    .Y(_1096_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1496_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1096_),
    .Y(_1097_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1497_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1098_),
    .B(_1094_),
    .A(_1097_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1498_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1067_),
    .B(_1095_),
    .C(_1098_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[8] ),
    .Y(_1099_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1499_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1099_),
    .Y(_0037_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1500_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1084_),
    .B(_1095_),
    .C(_1098_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[9] ),
    .Y(_1100_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1501_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1100_),
    .Y(_0038_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1502_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1086_),
    .B(_1095_),
    .C(_1098_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[10] ),
    .Y(_1101_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1503_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1101_),
    .Y(_0039_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1504_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1088_),
    .B(_1095_),
    .C(_1098_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[11] ),
    .Y(_1102_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1505_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1102_),
    .Y(_0040_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1506_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1080_),
    .Y(_1103_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1507_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1103_),
    .Y(_1104_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1508_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1105_),
    .B(net16),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1509_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net16),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[2] ),
    .Y(_1106_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1510_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1104_),
    .B(_1105_),
    .C(_1106_),
    .Y(_1107_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1511_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1107_),
    .Y(_0041_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1512_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1108_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1513_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net17),
    .A(_1108_),
    .Y(_1109_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1514_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net10),
    .Y(_1110_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1515_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1110_),
    .Y(_1111_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1516_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1109_),
    .A(_1106_),
    .Y(_1112_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1517_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1113_),
    .B(_1112_),
    .A(_1111_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1518_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0042_),
    .C(_1113_),
    .B(_1109_),
    .A(_1106_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1519_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net17),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[3] ),
    .Y(_1114_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1520_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1114_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[2] ),
    .B(_0938_),
    .C(_1109_),
    .Y(_1115_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1521_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1116_),
    .B(_1115_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1522_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1115_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[4] ),
    .Y(_1117_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1523_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1104_),
    .B(_1116_),
    .C(_1117_),
    .Y(_1118_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1524_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1118_),
    .Y(_0043_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1525_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1119_),
    .B(_1117_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1526_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1117_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[5] ),
    .Y(_1120_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1527_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1104_),
    .B(_1119_),
    .C(_1120_),
    .Y(_1121_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1528_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1121_),
    .Y(_0044_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1529_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1120_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[6] ),
    .Y(_1122_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1530_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[4] ),
    .B(\tt_um_rejunity_ay8913.pwm_master.accumulator[5] ),
    .C(\tt_um_rejunity_ay8913.pwm_master.accumulator[6] ),
    .D(_1115_),
    .Y(_1123_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1531_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1123_),
    .A(_1110_),
    .Y(_1124_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1532_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1124_),
    .A(_1122_),
    .Y(_1125_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1533_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1125_),
    .Y(_0045_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1534_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1126_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1535_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1127_),
    .B(_1123_),
    .A(_1126_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1536_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1080_),
    .Y(_1128_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1537_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1129_),
    .A(_1126_),
    .B(_1123_),
    .C(_1128_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1538_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0046_),
    .B(_1129_),
    .A(_1127_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1539_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1127_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[8] ),
    .Y(_1130_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1540_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1127_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[8] ),
    .Y(_1131_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1541_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1132_),
    .B(_1131_),
    .A(_1111_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1542_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0047_),
    .B(_1132_),
    .A(_1130_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1543_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1079_),
    .Y(_1133_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1544_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1133_),
    .Y(_1134_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1545_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1134_),
    .Y(_1135_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1546_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1136_),
    .B(_1130_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1547_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1130_),
    .A(\tt_um_rejunity_ay8913.pwm_master.accumulator[9] ),
    .Y(_1137_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1548_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1135_),
    .B(_1136_),
    .C(_1137_),
    .Y(_1138_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1549_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1138_),
    .Y(_0048_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1550_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1110_),
    .Y(_1139_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1551_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1137_),
    .A(_1139_),
    .Y(_1140_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1552_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1140_),
    .Y(_0049_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1553_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net10),
    .Y(_1141_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1554_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1141_),
    .Y(_1142_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1555_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[4] ),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[3] ),
    .Y(_1143_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1556_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1143_),
    .Y(_1144_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1557_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[0] ),
    .Y(_1145_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1558_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1143_),
    .A(_1077_),
    .Y(_1146_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1559_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1147_),
    .B(_1146_),
    .A(_1145_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1560_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1147_),
    .Y(_1148_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1561_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1148_),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[2] ),
    .Y(_1149_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1562_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1149_),
    .A(_1142_),
    .B(net16),
    .C(_1144_),
    .Y(_1150_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1563_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1150_),
    .Y(_0050_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1564_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1151_),
    .B(_1146_),
    .A(_1145_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1565_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[3] ),
    .B(_1147_),
    .C(_1151_),
    .D(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[2] ),
    .Y(_1152_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1566_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1152_),
    .A(_1142_),
    .B(net17),
    .C(_1144_),
    .Y(_1153_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1567_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1153_),
    .Y(_0051_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1568_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1148_),
    .Y(_0129_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1569_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1151_),
    .Y(_0096_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1570_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[4] ),
    .B(_0129_),
    .C(_0096_),
    .D(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[3] ),
    .Y(_1154_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1571_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1154_),
    .Y(_0052_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1572_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[5] ),
    .B(_0129_),
    .C(_0096_),
    .D(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[4] ),
    .Y(_1155_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1573_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1155_),
    .Y(_0053_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1574_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[6] ),
    .B(_0129_),
    .C(_0096_),
    .D(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[5] ),
    .Y(_1156_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1575_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1156_),
    .Y(_0054_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1576_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1148_),
    .Y(_1157_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1577_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1151_),
    .Y(_1158_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1578_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[7] ),
    .B(_1157_),
    .C(_1158_),
    .D(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[6] ),
    .Y(_1159_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1579_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1159_),
    .Y(_0055_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1580_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[8] ),
    .B(_1157_),
    .C(_1158_),
    .D(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[7] ),
    .Y(_1160_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1581_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1160_),
    .Y(_0056_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1582_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[9] ),
    .B(_1157_),
    .C(_1158_),
    .D(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[8] ),
    .Y(_1161_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1583_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1161_),
    .Y(_0057_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1584_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[10] ),
    .B(_1157_),
    .C(_1158_),
    .D(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[9] ),
    .Y(_1162_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1585_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1162_),
    .Y(_0058_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1586_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[11] ),
    .B(_1148_),
    .C(_1151_),
    .D(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[10] ),
    .Y(_1163_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1587_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1163_),
    .Y(_0059_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1588_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1164_),
    .B(_0925_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1589_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0925_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[2] ),
    .Y(_1165_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1590_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1135_),
    .B(_1164_),
    .C(_1165_),
    .Y(_1166_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1591_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1166_),
    .Y(_0060_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1592_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1167_),
    .B(_1165_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1593_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1165_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[3] ),
    .Y(_1168_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1594_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1135_),
    .B(_1167_),
    .C(_1168_),
    .Y(_1169_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1595_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1169_),
    .Y(_0061_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1596_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1170_),
    .B(_1168_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1597_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1168_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[4] ),
    .Y(_1171_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1598_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1135_),
    .B(_1170_),
    .C(_1171_),
    .Y(_1172_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1599_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1172_),
    .Y(_0062_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1600_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1134_),
    .Y(_1173_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1601_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1174_),
    .B(_1171_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1602_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1171_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[5] ),
    .Y(_1175_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1603_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1173_),
    .B(_1174_),
    .C(_1175_),
    .Y(_1176_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1604_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1176_),
    .Y(_0063_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1605_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1177_),
    .B(_1175_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1606_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1175_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[6] ),
    .Y(_1178_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1607_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1173_),
    .B(_1177_),
    .C(_1178_),
    .Y(_1179_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1608_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1179_),
    .Y(_0064_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1609_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1180_),
    .B(_1178_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1610_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1178_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[7] ),
    .Y(_1181_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1611_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1173_),
    .B(_1180_),
    .C(_1181_),
    .Y(_1182_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1612_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1182_),
    .Y(_0065_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1613_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1183_),
    .B(_1181_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1614_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1181_),
    .A(\tt_um_rejunity_ay8913.pwm_C.accumulator[8] ),
    .Y(_1184_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1615_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1173_),
    .B(_1183_),
    .C(_1184_),
    .Y(_1185_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1616_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1185_),
    .Y(_0066_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1617_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1184_),
    .A(_1139_),
    .Y(_1186_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1618_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1186_),
    .Y(_0067_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1619_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1134_),
    .Y(_1187_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1620_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1188_),
    .B(_0931_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1621_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0931_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[2] ),
    .Y(_1189_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1622_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1187_),
    .B(_1188_),
    .C(_1189_),
    .Y(_1190_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1623_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1190_),
    .Y(_0068_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1624_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1191_),
    .B(_1189_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1625_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1189_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[3] ),
    .Y(_1192_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1626_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1187_),
    .B(_1191_),
    .C(_1192_),
    .Y(_1193_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1627_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1193_),
    .Y(_0069_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1628_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1194_),
    .B(_1192_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1629_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1192_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[4] ),
    .Y(_1195_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1630_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1187_),
    .B(_1194_),
    .C(_1195_),
    .Y(_1196_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1631_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1196_),
    .Y(_0070_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1632_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1197_),
    .B(_1195_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1633_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1195_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[5] ),
    .Y(_1198_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1634_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1187_),
    .B(_1197_),
    .C(_1198_),
    .Y(_1199_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1635_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1199_),
    .Y(_0071_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1636_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1134_),
    .Y(_1200_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1637_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1201_),
    .B(_1198_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1638_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1198_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[6] ),
    .Y(_1202_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1639_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1200_),
    .B(_1201_),
    .C(_1202_),
    .Y(_1203_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1640_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1203_),
    .Y(_0072_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1641_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1204_),
    .B(_1202_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1642_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1202_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[7] ),
    .Y(_1205_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1643_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1200_),
    .B(_1204_),
    .C(_1205_),
    .Y(_1206_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1644_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1206_),
    .Y(_0073_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1645_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1207_),
    .B(_1205_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1646_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1205_),
    .A(\tt_um_rejunity_ay8913.pwm_B.accumulator[8] ),
    .Y(_1208_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1647_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1200_),
    .B(_1207_),
    .C(_1208_),
    .Y(_1209_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1648_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1209_),
    .Y(_0074_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1649_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1208_),
    .A(_1139_),
    .Y(_1210_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1650_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1210_),
    .Y(_0075_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1651_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1211_),
    .B(_1069_),
    .A(_1068_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1652_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1211_),
    .A(_1074_),
    .Y(_1212_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1653_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1212_),
    .Y(_1213_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1654_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1078_),
    .Y(_1214_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1655_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1215_),
    .B(_1212_),
    .A(_1214_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1656_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1215_),
    .Y(_1216_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1657_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1067_),
    .B(_1213_),
    .C(_1216_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[0] ),
    .Y(_1217_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1658_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1217_),
    .Y(_0076_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1659_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1084_),
    .B(_1213_),
    .C(_1216_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[1] ),
    .Y(_1218_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1660_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1218_),
    .Y(_0077_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1661_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1086_),
    .B(_1213_),
    .C(_1216_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[2] ),
    .Y(_1219_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1662_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1219_),
    .Y(_0078_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1663_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1088_),
    .B(_1213_),
    .C(_1216_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[3] ),
    .Y(_1220_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1664_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1220_),
    .Y(_0079_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1665_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1212_),
    .Y(_1221_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1666_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1215_),
    .Y(_1222_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1667_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1091_),
    .B(_1221_),
    .C(_1222_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[4] ),
    .Y(_1223_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1668_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1223_),
    .Y(_0080_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1669_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net5),
    .Y(_1224_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1670_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1224_),
    .B(_1221_),
    .C(_1222_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[5] ),
    .Y(_1225_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1671_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1225_),
    .Y(_0081_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1672_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net6),
    .Y(_1226_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1673_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1226_),
    .B(_1221_),
    .C(_1222_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[6] ),
    .Y(_1227_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1674_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1227_),
    .Y(_0082_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1675_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net7),
    .Y(_1228_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1676_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1228_),
    .B(_1221_),
    .C(_1222_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.period[7] ),
    .Y(_1229_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1677_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1229_),
    .Y(_0083_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1678_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.latched_register[0] ),
    .A(\tt_um_rejunity_ay8913.latched_register[1] ),
    .Y(_1230_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1679_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.latched_register[3] ),
    .B(\tt_um_rejunity_ay8913.latched_register[2] ),
    .C(_1073_),
    .Y(_1231_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1680_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1231_),
    .A(_1230_),
    .Y(_1232_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1681_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1232_),
    .Y(_1233_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1682_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1234_),
    .B(_1232_),
    .A(_1097_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1683_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1067_),
    .B(_1233_),
    .C(_1234_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[8] ),
    .Y(_1235_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1684_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1235_),
    .Y(_0084_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1685_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1084_),
    .B(_1233_),
    .C(_1234_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[9] ),
    .Y(_1236_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1686_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1236_),
    .Y(_0085_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1687_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1086_),
    .B(_1233_),
    .C(_1234_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[10] ),
    .Y(_1237_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1688_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1237_),
    .Y(_0086_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1689_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1088_),
    .B(_1233_),
    .C(_1234_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[11] ),
    .Y(_1238_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1690_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1238_),
    .Y(_0087_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1691_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[0]),
    .Y(_1239_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1692_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1231_),
    .A(_1070_),
    .Y(_1240_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1693_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1240_),
    .Y(_1241_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1694_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1242_),
    .B(_1240_),
    .A(_1214_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1695_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1242_),
    .Y(_1243_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1696_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1239_),
    .B(_1241_),
    .C(_1243_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[0] ),
    .Y(_1244_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1697_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1244_),
    .Y(_0088_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1698_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[1]),
    .Y(_1245_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1699_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1245_),
    .B(_1241_),
    .C(_1243_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[1] ),
    .Y(_1246_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1700_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1246_),
    .Y(_0089_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1701_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[2]),
    .Y(_1247_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1702_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1247_),
    .B(_1241_),
    .C(_1243_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[2] ),
    .Y(_1248_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1703_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1248_),
    .Y(_0090_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1704_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[3]),
    .Y(_1249_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1705_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1249_),
    .B(_1241_),
    .C(_1243_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[3] ),
    .Y(_1250_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1706_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1250_),
    .Y(_0091_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1707_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1240_),
    .Y(_1251_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1708_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1242_),
    .Y(_1252_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1709_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1091_),
    .B(_1251_),
    .C(_1252_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[4] ),
    .Y(_1253_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1710_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1253_),
    .Y(_0092_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1711_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1224_),
    .B(_1251_),
    .C(_1252_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[5] ),
    .Y(_1254_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1712_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1254_),
    .Y(_0093_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1713_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1226_),
    .B(_1251_),
    .C(_1252_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[6] ),
    .Y(_1255_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1714_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1255_),
    .Y(_0094_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1715_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1228_),
    .B(_1251_),
    .C(_1252_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.period[7] ),
    .Y(_1256_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1716_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1256_),
    .Y(_0095_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1717_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1146_),
    .Y(_1257_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1718_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1258_),
    .B(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[1] ),
    .A(_1145_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1719_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[1] ),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[0] ),
    .Y(_1259_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1720_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1257_),
    .B(_1258_),
    .C(_1259_),
    .Y(_1260_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1721_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1260_),
    .Y(_0097_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1722_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1261_),
    .B(_1259_),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1723_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1259_),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[2] ),
    .Y(_1262_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1724_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1257_),
    .B(_1261_),
    .C(_1262_),
    .Y(_1263_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1725_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1263_),
    .Y(_0098_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1726_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1262_),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[3] ),
    .Y(_1264_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1727_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0099_),
    .B(_1264_),
    .A(_1257_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1728_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1265_),
    .C(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[4] ),
    .B(_1262_),
    .A(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1729_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0100_),
    .B(_1265_),
    .A(_1257_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1730_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1266_),
    .B(_0936_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1731_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0936_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[2] ),
    .Y(_1267_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1732_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1200_),
    .B(_1266_),
    .C(_1267_),
    .Y(_1268_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1733_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1268_),
    .Y(_0101_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1734_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1133_),
    .Y(_1269_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1735_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1269_),
    .Y(_1270_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1736_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0257_),
    .B(_1267_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1737_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1267_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[3] ),
    .Y(_0258_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1738_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1270_),
    .B(_0257_),
    .C(_0258_),
    .Y(_0259_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1739_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0259_),
    .Y(_0102_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1740_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0260_),
    .B(_0258_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1741_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0258_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[4] ),
    .Y(_0261_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1742_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1270_),
    .B(_0260_),
    .C(_0261_),
    .Y(_0262_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1743_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0262_),
    .Y(_0103_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1744_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0263_),
    .B(_0261_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1745_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0261_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[5] ),
    .Y(_0264_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1746_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1270_),
    .B(_0263_),
    .C(_0264_),
    .Y(_0265_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1747_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0265_),
    .Y(_0104_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1748_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0266_),
    .B(_0264_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1749_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0264_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[6] ),
    .Y(_0267_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1750_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1270_),
    .B(_0266_),
    .C(_0267_),
    .Y(_0268_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1751_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0268_),
    .Y(_0105_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1752_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1269_),
    .Y(_0269_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1753_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0270_),
    .B(_0267_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1754_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0267_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[7] ),
    .Y(_0271_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1755_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0269_),
    .B(_0270_),
    .C(_0271_),
    .Y(_0272_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1756_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0272_),
    .Y(_0106_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1757_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0273_),
    .B(_0271_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1758_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0271_),
    .A(\tt_um_rejunity_ay8913.pwm_A.accumulator[8] ),
    .Y(_0274_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1759_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0269_),
    .B(_0273_),
    .C(_0274_),
    .Y(_0275_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1760_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0275_),
    .Y(_0107_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1761_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1142_),
    .Y(_0276_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1762_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0274_),
    .A(_0276_),
    .Y(_0277_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1763_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0277_),
    .Y(_0108_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1764_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0278_),
    .A(\tt_um_rejunity_ay8913.latched_register[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1765_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0278_),
    .B(\tt_um_rejunity_ay8913.latched_register[2] ),
    .C(_1073_),
    .Y(_0279_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1766_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0279_),
    .A(_1211_),
    .Y(_0280_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1767_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0281_),
    .B(_0280_),
    .A(_1128_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1768_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1239_),
    .B(_0280_),
    .C(_0281_),
    .D(\tt_um_rejunity_ay8913.amplitude_A[0] ),
    .Y(_0282_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1769_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0282_),
    .Y(_0109_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1770_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1091_),
    .B(_0280_),
    .C(_0281_),
    .D(\tt_um_rejunity_ay8913.envelope_A ),
    .Y(_0283_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1771_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0283_),
    .Y(_0110_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1772_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0278_),
    .B(_1071_),
    .C(_1073_),
    .Y(_0284_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1773_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0284_),
    .A(_1211_),
    .Y(_0285_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1774_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0285_),
    .Y(_0286_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1775_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0287_),
    .B(_0285_),
    .A(_1214_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1776_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0287_),
    .Y(_0288_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1777_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1239_),
    .B(_0286_),
    .C(_0288_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[8] ),
    .Y(_0289_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1778_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0289_),
    .Y(_0111_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1779_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1245_),
    .B(_0286_),
    .C(_0288_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[9] ),
    .Y(_0290_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1780_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0290_),
    .Y(_0112_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1781_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1247_),
    .B(_0286_),
    .C(_0288_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[10] ),
    .Y(_0291_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1782_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0291_),
    .Y(_0113_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1783_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1249_),
    .B(_0286_),
    .C(_0288_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[11] ),
    .Y(_0292_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1784_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0292_),
    .Y(_0114_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1785_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1090_),
    .Y(_0293_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1786_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0285_),
    .Y(_0294_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1787_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0287_),
    .Y(_0295_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1788_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0293_),
    .B(_0294_),
    .C(_0295_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[12] ),
    .Y(_0296_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1789_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0296_),
    .Y(_0115_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1790_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1224_),
    .B(_0294_),
    .C(_0295_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[13] ),
    .Y(_0297_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1791_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0297_),
    .Y(_0116_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1792_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1226_),
    .B(_0294_),
    .C(_0295_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[14] ),
    .Y(_0298_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1793_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0298_),
    .Y(_0117_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1794_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1228_),
    .B(_0294_),
    .C(_0295_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[15] ),
    .Y(_0299_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1795_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0299_),
    .Y(_0118_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1796_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1231_),
    .A(_1211_),
    .Y(_0300_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1797_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0300_),
    .Y(_0301_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1798_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0302_),
    .B(_0300_),
    .A(_1214_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1799_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0302_),
    .Y(_0303_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1800_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1239_),
    .B(_0301_),
    .C(_0303_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[0] ),
    .Y(_0304_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1801_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0304_),
    .Y(_0119_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1802_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1245_),
    .B(_0301_),
    .C(_0303_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[1] ),
    .Y(_0305_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1803_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0305_),
    .Y(_0120_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1804_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1247_),
    .B(_0301_),
    .C(_0303_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[2] ),
    .Y(_0306_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1805_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0306_),
    .Y(_0121_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1806_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1249_),
    .B(_0301_),
    .C(_0303_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[3] ),
    .Y(_0307_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1807_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0307_),
    .Y(_0122_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1808_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0300_),
    .Y(_0308_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1809_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0302_),
    .Y(_0309_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1810_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0293_),
    .B(_0308_),
    .C(_0309_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[4] ),
    .Y(_0310_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1811_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0310_),
    .Y(_0123_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1812_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1224_),
    .B(_0308_),
    .C(_0309_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[5] ),
    .Y(_0311_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1813_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0311_),
    .Y(_0124_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1814_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1226_),
    .B(_0308_),
    .C(_0309_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[6] ),
    .Y(_0312_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1815_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0312_),
    .Y(_0125_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1816_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1228_),
    .B(_0308_),
    .C(_0309_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[7] ),
    .Y(_0313_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1817_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0313_),
    .Y(_0126_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1818_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0127_),
    .B(_1144_),
    .A(_1139_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1819_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0314_),
    .B(_1144_),
    .A(_1145_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _1820_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_0314_),
    .B(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[11] ),
    .A(\tt_um_rejunity_ay8913.DAC_dat ),
    .Y(_0315_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1821_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0315_),
    .A(_0276_),
    .Y(_0316_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1822_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0316_),
    .Y(_0128_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1823_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0317_),
    .B(_1142_),
    .A(\tt_um_rejunity_ay8913.noise_generator.signal_edge.signal ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1824_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0130_),
    .A(_0317_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1825_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[0]),
    .Y(_0318_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1826_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1230_),
    .A(_1074_),
    .Y(_0319_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1827_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0319_),
    .Y(_0320_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1828_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0321_),
    .B(_0319_),
    .A(_1096_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1829_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0321_),
    .Y(_0322_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1830_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0318_),
    .B(_0320_),
    .C(_0322_),
    .D(\tt_um_rejunity_ay8913.tone_disable_A ),
    .Y(_0323_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1831_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0323_),
    .Y(_0131_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1832_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1245_),
    .B(_0320_),
    .C(_0322_),
    .D(\tt_um_rejunity_ay8913.tone_disable_B ),
    .Y(_0324_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1833_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0324_),
    .Y(_0132_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1834_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1247_),
    .B(_0320_),
    .C(_0322_),
    .D(\tt_um_rejunity_ay8913.tone_disable_C ),
    .Y(_0325_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1835_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0325_),
    .Y(_0133_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1836_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1249_),
    .B(_0320_),
    .C(_0322_),
    .D(\tt_um_rejunity_ay8913.noise_disable_A ),
    .Y(_0326_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1837_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0326_),
    .Y(_0134_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1838_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0293_),
    .B(_0319_),
    .C(_0321_),
    .D(\tt_um_rejunity_ay8913.noise_disable_B ),
    .Y(_0327_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1839_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0327_),
    .Y(_0135_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1840_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net5),
    .B(_0319_),
    .C(_0321_),
    .D(\tt_um_rejunity_ay8913.noise_disable_C ),
    .Y(_0328_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1841_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0328_),
    .Y(_0136_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1842_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0284_),
    .A(_1093_),
    .Y(_0329_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1843_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0329_),
    .Y(_0137_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1844_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0330_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0 ),
    .A(\tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1845_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0331_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.hold ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1846_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0332_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.stop ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1847_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0332_),
    .A(\tt_um_rejunity_ay8913.envelope_continue ),
    .B(_0331_),
    .C(_0330_),
    .Y(_0333_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1848_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0333_),
    .A(_0330_),
    .Y(_0334_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1849_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0334_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[0] ),
    .Y(_0335_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1850_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0336_),
    .B(_0334_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1851_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.restart_envelope ),
    .A(_1096_),
    .Y(_0337_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1852_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0337_),
    .Y(_0338_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1853_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0335_),
    .B(_0336_),
    .C(_0338_),
    .Y(_0339_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1854_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0339_),
    .Y(_0138_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1855_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0340_),
    .B(_0335_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1856_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0335_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[1] ),
    .Y(_0341_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1857_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0338_),
    .B(_0340_),
    .C(_0341_),
    .Y(_0342_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1858_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0342_),
    .Y(_0139_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1859_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0343_),
    .B(_0341_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1860_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0341_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[2] ),
    .Y(_0344_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1861_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0338_),
    .B(_0343_),
    .C(_0344_),
    .Y(_0345_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1862_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0345_),
    .Y(_0140_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1863_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0344_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[3] ),
    .Y(_0346_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1864_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0347_),
    .C(_0337_),
    .B(_0344_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1865_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0347_),
    .A(_0346_),
    .Y(_0348_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1866_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0348_),
    .Y(_0141_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1867_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[0] ),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[1] ),
    .Y(_0349_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1868_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[3] ),
    .B(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[2] ),
    .C(_0330_),
    .D(_0349_),
    .Y(_0350_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1869_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0142_),
    .C(_0338_),
    .B(_0350_),
    .A(_0333_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1870_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0351_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[15] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1871_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0352_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[15] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1872_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0353_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[14] ));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _1873_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0354_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[15] ),
    .B(_0352_),
    .C(_0353_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[14] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1874_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0355_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[14] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1875_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0356_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[13] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1876_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0355_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[14] ),
    .C(\tt_um_rejunity_ay8913.envelope_generator.period[13] ),
    .D(_0356_),
    .Y(_0357_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1877_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0358_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[12] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1878_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0359_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[12] ),
    .A(_0358_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1879_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0360_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[9] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1880_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0361_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[8] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1881_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[9] ),
    .B(_0360_),
    .C(_0361_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[8] ),
    .Y(_0362_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1882_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0360_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[9] ),
    .Y(_0363_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1883_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[10] ),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[10] ),
    .Y(_0364_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1884_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[11] ),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[11] ),
    .Y(_0365_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1885_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0365_),
    .A(_0364_),
    .Y(_0366_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1886_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0367_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[11] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1887_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[10] ),
    .Y(_0368_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1888_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0369_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[10] ),
    .A(_0368_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1889_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0370_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[11] ),
    .B(_0367_),
    .C(_0369_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1890_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0370_),
    .A(_0362_),
    .B(_0363_),
    .C(_0366_),
    .Y(_0371_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1891_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0372_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[13] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1892_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0373_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[12] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1893_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[13] ),
    .B(_0372_),
    .C(_0373_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[12] ),
    .Y(_0374_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1894_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0375_),
    .C(_0374_),
    .B(_0371_),
    .A(_0359_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1895_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0375_),
    .A(_0357_),
    .Y(_0376_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1896_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0351_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[15] ),
    .C(_0354_),
    .D(_0376_),
    .Y(_0377_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1897_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0378_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[7] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1898_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0379_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[6] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1899_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[5] ),
    .Y(_0380_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1900_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0381_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[5] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1901_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0382_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1902_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0383_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[3] ),
    .A(_0382_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1903_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0384_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[2] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1904_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0385_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1905_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0386_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[0] ),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1906_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0387_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[1] ),
    .B(_0385_),
    .C(_0386_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1907_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0388_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[2] ),
    .B(_0384_),
    .C(_0387_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1908_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0389_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[3] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1909_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0390_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.period[4] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1910_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[3] ),
    .B(_0389_),
    .C(_0390_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[4] ),
    .Y(_0391_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1911_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0392_),
    .A(_0383_),
    .B(_0388_),
    .C(_0391_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1912_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0393_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1913_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0394_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _1914_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0395_),
    .A(_0393_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[5] ),
    .C(\tt_um_rejunity_ay8913.envelope_generator.period[4] ),
    .D(_0394_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1915_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0380_),
    .B(_0381_),
    .C(_0392_),
    .D(_0395_),
    .Y(_0396_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1916_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0397_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[6] ),
    .B(_0379_),
    .C(_0396_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1917_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0398_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[7] ),
    .B(_0378_),
    .C(_0397_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1918_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0357_),
    .B(_0362_),
    .C(_0374_),
    .Y(_0399_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1919_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0354_),
    .B(_0359_),
    .C(_0363_),
    .D(_0366_),
    .Y(_0400_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1920_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0401_),
    .A(_0400_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1921_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0402_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1922_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0403_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1923_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0403_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[7] ),
    .C(\tt_um_rejunity_ay8913.envelope_generator.period[15] ),
    .D(_0351_),
    .Y(_0404_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1924_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0405_),
    .C(_0404_),
    .B(\tt_um_rejunity_ay8913.envelope_generator.period[8] ),
    .A(_0402_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1925_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0398_),
    .B(_0399_),
    .C(_0401_),
    .D(_0405_),
    .Y(_0406_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1926_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0407_),
    .A(net2));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1927_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0408_),
    .B(\tt_um_rejunity_ay8913.clk_counter[1] ),
    .A(\tt_um_rejunity_ay8913.clk_counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1928_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0409_),
    .A(\tt_um_rejunity_ay8913.clk_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_4 _1929_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0407_),
    .B(net1),
    .C(_0408_),
    .D(_0409_),
    .Y(_0410_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1930_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0410_),
    .Y(_0411_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1931_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0412_),
    .B(\tt_um_rejunity_ay8913.clk_counter[5] ),
    .A(\tt_um_rejunity_ay8913.clk_counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1932_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0413_),
    .B(\tt_um_rejunity_ay8913.clk_counter[6] ),
    .A(\tt_um_rejunity_ay8913.clk_counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1933_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0414_),
    .B(net2),
    .A(net1));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1934_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0415_),
    .A(_0412_),
    .B(_0413_),
    .C(_0414_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1935_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0415_),
    .Y(_0416_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1936_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0417_),
    .B(_0416_),
    .A(_0411_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1937_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0418_),
    .A(_0377_),
    .B(_0406_),
    .C(_0417_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1938_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0419_),
    .B(\tt_um_rejunity_ay8913.restart_envelope ),
    .A(_1078_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1939_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0420_),
    .B(_0418_),
    .A(_0419_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1940_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0420_),
    .Y(_0421_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1941_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0422_),
    .B(_0419_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1942_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal ),
    .B(_0418_),
    .C(_0421_),
    .D(_0422_),
    .Y(_0423_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1943_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0423_),
    .Y(_0143_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1944_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0420_),
    .Y(_0424_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1945_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0417_),
    .Y(_0425_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1946_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0425_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[0] ),
    .Y(_0426_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1947_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0426_),
    .A(_0424_),
    .Y(_0427_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1948_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0427_),
    .Y(_0144_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1949_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0421_),
    .Y(_0428_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1950_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0411_),
    .Y(_0429_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1951_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0416_),
    .Y(_0430_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1952_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[1] ),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[0] ),
    .B(_0429_),
    .C(_0430_),
    .Y(_0431_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1953_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[1] ),
    .B(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[0] ),
    .C(_0411_),
    .D(_0416_),
    .Y(_0432_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1954_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0433_),
    .B(_0432_),
    .A(_0431_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1955_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0145_),
    .B(_0433_),
    .A(_0428_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1956_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0421_),
    .Y(_0434_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1957_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0435_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1958_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0436_),
    .B(_0432_),
    .A(_0435_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1959_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0432_),
    .A(_0435_),
    .Y(_0437_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1960_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0434_),
    .B(_0436_),
    .C(_0437_),
    .Y(_0438_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1961_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0438_),
    .Y(_0146_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1962_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0439_),
    .B(_0436_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1963_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0382_),
    .B(_0435_),
    .C(_0432_),
    .Y(_0440_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1964_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0440_),
    .Y(_0441_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1965_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0434_),
    .B(_0439_),
    .C(_0441_),
    .Y(_0442_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1966_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0442_),
    .Y(_0147_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1967_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[4] ),
    .Y(_0443_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1968_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0441_),
    .A(_0443_),
    .Y(_0444_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1969_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0445_),
    .B(_0441_),
    .A(_0443_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1970_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0434_),
    .B(_0444_),
    .C(_0445_),
    .Y(_0446_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1971_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0446_),
    .Y(_0148_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1972_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0444_),
    .A(_0380_),
    .Y(_0447_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1973_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0149_),
    .B(_0447_),
    .A(_0428_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1974_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[6] ),
    .A(_0380_),
    .B(_0443_),
    .C(_0441_),
    .Y(_0448_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1975_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[6] ),
    .B(_0380_),
    .C(_0443_),
    .D(_0440_),
    .Y(_0449_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1976_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0450_),
    .B(_0449_),
    .A(_0448_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1977_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0150_),
    .B(_0450_),
    .A(_0428_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1978_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0449_),
    .A(_0403_),
    .Y(_0451_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1979_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0452_),
    .B(_0449_),
    .A(_0403_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1980_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0424_),
    .B(_0451_),
    .C(_0452_),
    .Y(_0453_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1981_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0453_),
    .Y(_0151_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1982_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0452_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[8] ),
    .Y(_0454_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1983_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0152_),
    .B(_0454_),
    .A(_0428_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1984_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0421_),
    .Y(_0455_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1985_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[9] ),
    .Y(_0456_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1986_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0402_),
    .B(_0403_),
    .C(_0449_),
    .Y(_0457_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1987_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0457_),
    .A(_0456_),
    .Y(_0458_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1988_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0153_),
    .B(_0458_),
    .A(_0455_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1989_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0457_),
    .A(_0456_),
    .Y(_0459_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1990_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0459_),
    .A(_0368_),
    .Y(_0460_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1991_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0154_),
    .B(_0460_),
    .A(_0455_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1992_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[11] ),
    .A(_0368_),
    .B(_0456_),
    .C(_0457_),
    .Y(_0461_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _1993_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[11] ),
    .B(_0368_),
    .C(_0456_),
    .D(_0457_),
    .Y(_0462_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1994_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0463_),
    .B(_0462_),
    .A(_0461_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1995_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0155_),
    .B(_0463_),
    .A(_0455_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1996_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0462_),
    .A(_0358_),
    .Y(_0464_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1997_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0465_),
    .B(_0462_),
    .A(_0358_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1998_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0424_),
    .B(_0464_),
    .C(_0465_),
    .Y(_0466_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1999_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0466_),
    .Y(_0156_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2000_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0467_),
    .B(_0465_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[13] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2001_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0465_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[13] ),
    .Y(_0468_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2002_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0424_),
    .B(_0467_),
    .C(_0468_),
    .Y(_0469_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2003_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0469_),
    .Y(_0157_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2004_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0468_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[14] ),
    .Y(_0470_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2005_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0158_),
    .B(_0470_),
    .A(_0455_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2006_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0471_),
    .C(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[15] ),
    .B(_0468_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[14] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2007_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0159_),
    .B(_0471_),
    .A(_0434_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2008_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0472_),
    .A(\tt_um_rejunity_ay8913.envelope_attack ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2009_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0473_),
    .A(\tt_um_rejunity_ay8913.envelope_continue ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2010_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.envelope_alternate ),
    .A(\tt_um_rejunity_ay8913.envelope_generator.hold ),
    .Y(_0474_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2011_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0475_),
    .A(\tt_um_rejunity_ay8913.envelope_continue ),
    .B(_0474_),
    .C(_0350_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2012_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0476_),
    .A(_0473_),
    .B(\tt_um_rejunity_ay8913.envelope_attack ),
    .C(_0475_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2013_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0476_),
    .A(\tt_um_rejunity_ay8913.envelope_generator.invert_output ),
    .Y(_0477_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _2014_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_0419_),
    .B(_0477_),
    .A(_0472_),
    .Y(_0478_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2015_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0478_),
    .Y(_0160_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2016_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0479_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[1] ));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _2017_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0480_),
    .B(\tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0 ),
    .A(\tt_um_rejunity_ay8913.noise_generator.signal_edge.signal ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2018_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0480_),
    .Y(_0481_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2019_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0481_),
    .Y(_0482_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2020_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0482_),
    .Y(_0483_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2021_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0484_),
    .A(_0928_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _2022_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0485_),
    .B(\tt_um_rejunity_ay8913.noise_generator.signal_edge.signal ),
    .A(\tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0 ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2023_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0485_),
    .Y(_0486_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2024_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0487_),
    .A(_0484_),
    .B(_0486_),
    .C(_1269_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2025_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0161_),
    .C(_0487_),
    .B(_0483_),
    .A(_0479_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2026_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0488_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[2] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2027_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0489_),
    .A(_0479_),
    .B(_0486_),
    .C(_1269_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2028_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0162_),
    .C(_0489_),
    .B(_0483_),
    .A(_0488_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2029_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0490_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2030_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0491_),
    .B(_0481_),
    .A(_0490_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2031_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1079_),
    .Y(_0492_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2032_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0492_),
    .Y(_0493_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2033_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0494_),
    .C(_0493_),
    .B(_0486_),
    .A(_0488_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2034_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0494_),
    .A(_0491_),
    .Y(_0495_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2035_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0495_),
    .Y(_0163_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2036_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0496_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[4] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2037_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0492_),
    .Y(_0497_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2038_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0498_),
    .A(_0490_),
    .B(_0486_),
    .C(_0497_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2039_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0164_),
    .C(_0498_),
    .B(_0483_),
    .A(_0496_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2040_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0499_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[5] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2041_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0485_),
    .Y(_0500_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2042_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0500_),
    .Y(_0501_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2043_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0502_),
    .A(_0496_),
    .B(_0501_),
    .C(_0497_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2044_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0165_),
    .C(_0502_),
    .B(_0483_),
    .A(_0499_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2045_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0503_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[6] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2046_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0481_),
    .Y(_0504_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2047_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0505_),
    .A(_0499_),
    .B(_0501_),
    .C(_0497_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2048_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0166_),
    .C(_0505_),
    .B(_0504_),
    .A(_0503_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2049_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0506_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[7] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2050_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0507_),
    .A(_0503_),
    .B(_0501_),
    .C(_0497_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2051_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0167_),
    .C(_0507_),
    .B(_0504_),
    .A(_0506_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2052_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0508_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[8] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2053_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1133_),
    .Y(_0509_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2054_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0510_),
    .A(_0506_),
    .B(_0501_),
    .C(_0509_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2055_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0168_),
    .C(_0510_),
    .B(_0504_),
    .A(_0508_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2056_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0511_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[9] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2057_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0500_),
    .Y(_0512_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2058_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0513_),
    .A(_0508_),
    .B(_0512_),
    .C(_0509_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2059_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0169_),
    .C(_0513_),
    .B(_0504_),
    .A(_0511_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2060_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0514_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[10] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2061_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0481_),
    .Y(_0515_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2062_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0516_),
    .A(_0511_),
    .B(_0512_),
    .C(_0509_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2063_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0170_),
    .C(_0516_),
    .B(_0515_),
    .A(_0514_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2064_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0517_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[11] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2065_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0518_),
    .A(_0514_),
    .B(_0512_),
    .C(_0509_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2066_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0171_),
    .C(_0518_),
    .B(_0515_),
    .A(_0517_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2067_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0519_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[12] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2068_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1133_),
    .Y(_0520_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2069_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0521_),
    .A(_0517_),
    .B(_0512_),
    .C(_0520_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2070_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0172_),
    .C(_0521_),
    .B(_0515_),
    .A(_0519_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2071_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0522_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[13] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2072_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0500_),
    .Y(_0523_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2073_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0524_),
    .A(_0519_),
    .B(_0523_),
    .C(_0520_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2074_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0173_),
    .C(_0524_),
    .B(_0515_),
    .A(_0522_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2075_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0525_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[14] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2076_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0526_),
    .A(_0522_),
    .B(_0523_),
    .C(_0520_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2077_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0174_),
    .C(_0526_),
    .B(_0482_),
    .A(_0525_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2078_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0527_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[15] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2079_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0528_),
    .A(_0525_),
    .B(_0523_),
    .C(_0520_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2080_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0175_),
    .C(_0528_),
    .B(_0482_),
    .A(_0527_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2081_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0529_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[16] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2082_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0530_),
    .A(_0527_),
    .B(_0523_),
    .C(_1128_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2083_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0176_),
    .C(_0530_),
    .B(_0482_),
    .A(_0529_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2084_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[12] ),
    .B(\tt_um_rejunity_ay8913.noise_generator.lfsr[11] ),
    .C(\tt_um_rejunity_ay8913.noise_generator.lfsr[10] ),
    .Y(_0531_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2085_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0531_),
    .A(_0511_),
    .Y(_0532_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2086_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[16] ),
    .B(\tt_um_rejunity_ay8913.noise_generator.lfsr[15] ),
    .C(\tt_um_rejunity_ay8913.noise_generator.lfsr[14] ),
    .Y(_0533_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2087_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0533_),
    .A(_0522_),
    .Y(_0534_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2088_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0534_),
    .A(_0532_),
    .Y(_0535_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2089_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[8] ),
    .B(\tt_um_rejunity_ay8913.noise_generator.lfsr[7] ),
    .C(\tt_um_rejunity_ay8913.noise_generator.lfsr[6] ),
    .Y(_0536_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2090_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0536_),
    .A(_0499_),
    .Y(_0537_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2091_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[4] ),
    .B(\tt_um_rejunity_ay8913.noise_generator.lfsr[2] ),
    .C(\tt_um_rejunity_ay8913.noise_generator.lfsr[1] ),
    .Y(_0538_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2092_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0535_),
    .B(_0537_),
    .C(_0538_),
    .Y(_0539_),
    .D(_0491_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2093_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1080_),
    .A(\tt_um_rejunity_ay8913.noise_generator.lfsr[3] ),
    .B(_0928_),
    .C(_0480_),
    .Y(_0540_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2094_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0541_),
    .A(_0529_),
    .B(_0500_),
    .C(_0540_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2095_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0177_),
    .C(_0541_),
    .B(_0539_),
    .A(_0484_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2096_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0416_),
    .A(_0411_),
    .Y(_0542_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2097_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0542_),
    .Y(_0543_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2098_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0544_),
    .A(\tt_um_rejunity_ay8913.noise_generator.period[2] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2099_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0545_),
    .A(\tt_um_rejunity_ay8913.noise_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _2100_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0546_),
    .B(\tt_um_rejunity_ay8913.noise_generator.period[0] ),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2101_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0547_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[1] ),
    .B(_0545_),
    .C(_0546_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2102_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0548_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[2] ),
    .B(_0544_),
    .C(_0547_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2103_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0549_),
    .A(\tt_um_rejunity_ay8913.noise_generator.period[3] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2104_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0549_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[3] ),
    .Y(_0550_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2105_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0544_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[2] ),
    .Y(_0551_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2106_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0552_),
    .A(\tt_um_rejunity_ay8913.noise_generator.period[4] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2107_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[4] ),
    .B(_0552_),
    .C(_0549_),
    .D(\tt_um_rejunity_ay8913.noise_generator.tone.counter[3] ),
    .Y(_0553_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2108_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0553_),
    .A(_0548_),
    .B(_0550_),
    .C(_0551_),
    .Y(_0554_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2109_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0552_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[4] ),
    .Y(_0555_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _2110_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0543_),
    .B(_0554_),
    .C(_0555_),
    .Y(_0556_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2111_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0557_),
    .B(_0556_),
    .A(_1141_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2112_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.noise_generator.signal_edge.signal ),
    .B(_0556_),
    .C(_0557_),
    .D(_0317_),
    .Y(_0558_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2113_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0558_),
    .Y(_0178_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2114_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0425_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[0] ),
    .Y(_0559_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2115_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0559_),
    .A(_0557_),
    .Y(_0560_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2116_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0560_),
    .Y(_0179_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2117_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0557_),
    .Y(_0561_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2118_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0542_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[0] ),
    .Y(_0562_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2119_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0562_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[1] ),
    .Y(_0563_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2120_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0180_),
    .B(_0563_),
    .A(_0561_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2121_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0562_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[1] ),
    .Y(_0564_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2122_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0565_),
    .B(_0564_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2123_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0564_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[2] ),
    .Y(_0566_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2124_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0561_),
    .B(_0565_),
    .C(_0566_),
    .Y(_0567_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2125_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0567_),
    .Y(_0181_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2126_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0566_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[3] ),
    .Y(_0568_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2127_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0182_),
    .B(_0568_),
    .A(_0561_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2128_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0569_),
    .C(\tt_um_rejunity_ay8913.noise_generator.tone.counter[4] ),
    .B(_0566_),
    .A(\tt_um_rejunity_ay8913.noise_generator.tone.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2129_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0183_),
    .B(_0569_),
    .A(_0561_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2130_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0184_),
    .A(_0422_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2131_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0570_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2132_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[8] ),
    .Y(_0571_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2133_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0572_),
    .A(_0571_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _2134_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0573_),
    .A(_0570_),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.period[9] ),
    .C(\tt_um_rejunity_ay8913.tone_C_generator.period[8] ),
    .D(_0572_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2135_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0574_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.period[5] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2136_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0574_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[5] ),
    .Y(_0575_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2137_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0576_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.period[0] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2138_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0577_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2139_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[0] ),
    .B(_0576_),
    .C(_0577_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.counter[1] ),
    .Y(_0578_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2140_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0577_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[1] ),
    .Y(_0579_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _2141_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0580_),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.counter[3] ),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.period[3] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2142_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.period[2] ),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[2] ),
    .Y(_0581_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2143_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0582_),
    .B(_0581_),
    .A(_0580_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2144_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0583_),
    .A(_0578_),
    .B(_0579_),
    .C(_0582_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2145_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0584_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2146_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0585_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2147_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0586_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2148_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0585_),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.period[3] ),
    .C(\tt_um_rejunity_ay8913.tone_C_generator.period[4] ),
    .D(_0586_),
    .Y(_0587_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2149_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0584_),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.period[2] ),
    .C(_0580_),
    .Y(_0588_),
    .D(_0587_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2150_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0589_),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.period[4] ),
    .A(_0586_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2151_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0590_),
    .A(_0583_),
    .B(_0588_),
    .C(_0589_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2152_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0591_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.period[6] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2153_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[6] ),
    .B(_0591_),
    .C(_0574_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.counter[5] ),
    .Y(_0592_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2154_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0593_),
    .A(_0575_),
    .B(_0590_),
    .C(_0592_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2155_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0594_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2156_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0595_),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.period[6] ),
    .A(_0594_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2157_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0596_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.period[7] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2158_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0596_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[7] ),
    .Y(_0597_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2159_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[7] ),
    .Y(_0598_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2160_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0599_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.period[8] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2161_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0598_),
    .B(_0596_),
    .C(_0599_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.counter[8] ),
    .Y(_0600_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2162_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0600_),
    .A(_0593_),
    .B(_0595_),
    .C(_0597_),
    .Y(_0601_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2163_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.period[9] ),
    .A(_0570_),
    .Y(_0602_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2164_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0603_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.period[11] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2165_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0604_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.period[10] ));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _2166_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0605_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[11] ),
    .B(_0603_),
    .C(_0604_),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2167_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0604_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[10] ),
    .Y(_0606_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2168_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0606_),
    .A(_0605_),
    .Y(_0607_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2169_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0608_),
    .B(_0607_),
    .A(_0602_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2170_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0609_),
    .A(_0573_),
    .B(_0601_),
    .C(_0608_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2171_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0610_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[11] ),
    .B(_0603_),
    .C(_0606_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2172_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0570_),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.period[9] ),
    .C(\tt_um_rejunity_ay8913.tone_C_generator.period[8] ),
    .D(_0572_),
    .Y(_0611_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2173_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0603_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[11] ),
    .Y(_0612_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2174_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0575_),
    .B(_0579_),
    .C(_0597_),
    .D(_0612_),
    .Y(_0613_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2175_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0614_),
    .B(_0599_),
    .A(_0571_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2176_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[0] ),
    .Y(_0615_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2177_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0616_),
    .A(_0615_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2178_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0617_),
    .C(_0589_),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.period[0] ),
    .A(_0616_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _2179_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0614_),
    .B(_0602_),
    .C(_0617_),
    .Y(_0618_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2180_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0578_),
    .B(_0587_),
    .C(_0618_),
    .Y(_0619_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2181_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0580_),
    .B(_0581_),
    .C(_0607_),
    .D(_0619_),
    .Y(_0620_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2182_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0611_),
    .B(_0613_),
    .C(_0620_),
    .Y(_0621_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2183_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0598_),
    .B(_0596_),
    .C(\tt_um_rejunity_ay8913.tone_C_generator.period[6] ),
    .D(_0594_),
    .Y(_0622_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2184_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0623_),
    .B(_0622_),
    .A(_0592_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2185_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0609_),
    .B(_0610_),
    .C(_0621_),
    .D(_0623_),
    .Y(_0624_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2186_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0625_),
    .B(_0624_),
    .A(_0543_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2187_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0626_),
    .B(_0625_),
    .A(_1141_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2188_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0626_),
    .Y(_0627_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2189_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0425_),
    .A(_0615_),
    .Y(_0628_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2190_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0628_),
    .A(_0627_),
    .Y(_0629_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2191_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0629_),
    .Y(_0185_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2192_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0626_),
    .Y(_0630_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2193_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[1] ),
    .B(_0615_),
    .C(_0410_),
    .D(_0415_),
    .Y(_0631_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2194_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\tt_um_rejunity_ay8913.tone_C_generator.counter[1] ),
    .A(_0615_),
    .B(_0429_),
    .C(_0430_),
    .Y(_0632_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2195_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0633_),
    .B(_0632_),
    .A(_0631_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2196_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0186_),
    .B(_0633_),
    .A(_0630_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2197_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0626_),
    .Y(_0634_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2198_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0635_),
    .B(_0631_),
    .A(_0584_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2199_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0631_),
    .A(_0584_),
    .Y(_0636_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2200_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0634_),
    .B(_0635_),
    .C(_0636_),
    .Y(_0637_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2201_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0637_),
    .Y(_0187_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2202_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0585_),
    .B(_0584_),
    .C(_0631_),
    .Y(_0638_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2203_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0639_),
    .B(_0635_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2204_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0627_),
    .B(_0638_),
    .C(_0639_),
    .Y(_0640_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2205_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0640_),
    .Y(_0188_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2206_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0638_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[4] ),
    .Y(_0641_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2207_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0642_),
    .B(_0638_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2208_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0627_),
    .B(_0641_),
    .C(_0642_),
    .Y(_0643_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2209_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0643_),
    .Y(_0189_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2210_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0641_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[5] ),
    .Y(_0644_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2211_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0190_),
    .B(_0644_),
    .A(_0630_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _2212_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[5] ),
    .B(\tt_um_rejunity_ay8913.tone_C_generator.counter[4] ),
    .C(_0638_),
    .Y(_0645_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2213_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0645_),
    .A(_0594_),
    .Y(_0646_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2214_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0191_),
    .B(_0646_),
    .A(_0630_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2215_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0647_),
    .B(_0645_),
    .A(_0594_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2216_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0647_),
    .A(_0598_),
    .Y(_0648_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2217_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0192_),
    .B(_0648_),
    .A(_0630_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2218_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0647_),
    .A(_0598_),
    .Y(_0649_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2219_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0649_),
    .A(_0571_),
    .Y(_0650_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2220_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0193_),
    .B(_0650_),
    .A(_0634_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2221_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0649_),
    .A(_0571_),
    .Y(_0651_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2222_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0651_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[9] ),
    .Y(_0652_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2223_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0653_),
    .B(_0651_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2224_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0627_),
    .B(_0652_),
    .C(_0653_),
    .Y(_0654_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2225_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0654_),
    .Y(_0194_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2226_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0652_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[10] ),
    .Y(_0655_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2227_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0195_),
    .B(_0655_),
    .A(_0634_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2228_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0656_),
    .C(\tt_um_rejunity_ay8913.tone_C_generator.counter[11] ),
    .B(_0652_),
    .A(\tt_um_rejunity_ay8913.tone_C_generator.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2229_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0196_),
    .B(_0656_),
    .A(_0634_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2230_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0625_),
    .A(\tt_um_rejunity_ay8913.tone_C ),
    .Y(_0657_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2231_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0657_),
    .A(_0493_),
    .Y(_0658_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2232_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0658_),
    .Y(_0197_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2233_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1231_),
    .A(_1093_),
    .Y(_0659_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2234_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0659_),
    .Y(_0660_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2235_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0661_),
    .B(_0659_),
    .A(_1097_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2236_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0318_),
    .B(_0660_),
    .C(_0661_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[8] ),
    .Y(_0662_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2237_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0662_),
    .Y(_0198_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2238_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[1]),
    .Y(_0663_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2239_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0663_),
    .B(_0660_),
    .C(_0661_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[9] ),
    .Y(_0664_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2240_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0664_),
    .Y(_0199_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2241_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[2]),
    .Y(_0665_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2242_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0665_),
    .B(_0660_),
    .C(_0661_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[10] ),
    .Y(_0666_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2243_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0666_),
    .Y(_0200_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2244_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[3]),
    .Y(_0667_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2245_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0667_),
    .B(_0660_),
    .C(_0661_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.period[11] ),
    .Y(_0668_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2246_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0668_),
    .Y(_0201_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2247_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0669_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2248_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0670_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _2249_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0671_),
    .A(_0669_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[11] ),
    .C(\tt_um_rejunity_ay8913.tone_B_generator.period[10] ),
    .D(_0670_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2250_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0672_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[9] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2251_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0672_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[9] ),
    .Y(_0673_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2252_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[8] ),
    .Y(_0674_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2253_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0675_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[8] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2254_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0676_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2255_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0677_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _2256_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0678_),
    .A(_0676_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[7] ),
    .C(\tt_um_rejunity_ay8913.tone_B_generator.period[8] ),
    .D(_0677_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2257_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[7] ),
    .Y(_0679_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2258_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0680_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[7] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2259_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0681_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2260_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0682_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[6] ),
    .A(_0681_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2261_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0683_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[5] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2262_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0683_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[5] ),
    .Y(_0684_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2263_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0685_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[4] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2264_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0686_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2265_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0686_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[1] ),
    .Y(_0687_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2266_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0688_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[0] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2267_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[0] ),
    .B(_0688_),
    .C(_0686_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.counter[1] ),
    .Y(_0689_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _2268_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0690_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.counter[3] ),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[3] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2269_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[2] ),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[2] ),
    .Y(_0691_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2270_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0692_),
    .B(_0691_),
    .A(_0690_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2271_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0693_),
    .A(_0687_),
    .B(_0689_),
    .C(_0692_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2272_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0694_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2273_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0695_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2274_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0696_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2275_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0695_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[3] ),
    .C(\tt_um_rejunity_ay8913.tone_B_generator.period[4] ),
    .D(_0696_),
    .Y(_0697_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2276_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0694_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[2] ),
    .C(_0690_),
    .Y(_0698_),
    .D(_0697_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2277_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[4] ),
    .B(_0685_),
    .C(_0693_),
    .D(_0698_),
    .Y(_0699_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2278_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0700_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[6] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2279_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[6] ),
    .B(_0700_),
    .C(_0683_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.counter[5] ),
    .Y(_0701_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2280_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0702_),
    .A(_0684_),
    .B(_0699_),
    .C(_0701_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2281_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0679_),
    .B(_0680_),
    .C(_0682_),
    .D(_0702_),
    .Y(_0703_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2282_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0674_),
    .B(_0675_),
    .C(_0678_),
    .D(_0703_),
    .Y(_0704_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2283_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0705_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.period[10] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2284_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[10] ),
    .B(_0705_),
    .C(_0672_),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.counter[9] ),
    .Y(_0706_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2285_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0707_),
    .A(_0673_),
    .B(_0704_),
    .C(_0706_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2286_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0708_),
    .B(_0687_),
    .A(_0684_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2287_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0709_),
    .B(_0708_),
    .A(_0706_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2288_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[4] ),
    .Y(_0710_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _2289_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0711_),
    .A(_0681_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[6] ),
    .C(_0685_),
    .D(_0710_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2290_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0711_),
    .A(_0671_),
    .Y(_0712_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2291_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0712_),
    .A(_0709_),
    .Y(_0713_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2292_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0676_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[7] ),
    .C(\tt_um_rejunity_ay8913.tone_B_generator.period[8] ),
    .D(_0677_),
    .Y(_0714_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2293_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0701_),
    .A(_0714_),
    .Y(_0715_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2294_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0689_),
    .B(_0697_),
    .C(_0715_),
    .Y(_0716_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2295_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[0] ),
    .Y(_0717_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2296_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0718_),
    .A(_0717_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2297_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0718_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[0] ),
    .C(_0680_),
    .D(_0679_),
    .Y(_0719_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2298_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0720_),
    .A(_0674_),
    .B(_0675_),
    .C(_0719_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2299_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0721_),
    .B(_0720_),
    .A(_0692_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2300_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0721_),
    .A(_0716_),
    .Y(_0722_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2301_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0723_),
    .B(\tt_um_rejunity_ay8913.tone_B_generator.period[11] ),
    .A(_0669_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2302_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0723_),
    .A(_0673_),
    .B(_0713_),
    .C(_0722_),
    .Y(_0724_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2303_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0725_),
    .A(_0671_),
    .B(_0707_),
    .C(_0724_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2304_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0726_),
    .A(_0542_),
    .B(_0725_),
    .C(_1079_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2305_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0726_),
    .Y(_0727_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2306_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0425_),
    .A(_0717_),
    .Y(_0728_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2307_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0728_),
    .A(_0727_),
    .Y(_0729_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2308_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0729_),
    .Y(_0202_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2309_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0726_),
    .Y(_0730_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2310_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[1] ),
    .B(_0717_),
    .C(_0410_),
    .D(_0415_),
    .Y(_0731_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2311_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\tt_um_rejunity_ay8913.tone_B_generator.counter[1] ),
    .A(_0717_),
    .B(_0429_),
    .C(_0430_),
    .Y(_0732_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2312_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0733_),
    .B(_0732_),
    .A(_0731_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2313_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0203_),
    .B(_0733_),
    .A(_0730_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2314_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0726_),
    .Y(_0734_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2315_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0735_),
    .B(_0731_),
    .A(_0694_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2316_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0731_),
    .A(_0694_),
    .Y(_0736_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2317_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0734_),
    .B(_0735_),
    .C(_0736_),
    .Y(_0737_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2318_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0737_),
    .Y(_0204_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2319_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0695_),
    .B(_0694_),
    .C(_0731_),
    .Y(_0738_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2320_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0739_),
    .B(_0735_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2321_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0727_),
    .B(_0738_),
    .C(_0739_),
    .Y(_0740_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2322_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0740_),
    .Y(_0205_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2323_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0738_),
    .A(_0710_),
    .Y(_0741_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2324_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0742_),
    .B(_0738_),
    .A(_0710_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2325_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0727_),
    .B(_0741_),
    .C(_0742_),
    .Y(_0743_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2326_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0743_),
    .Y(_0206_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2327_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0741_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[5] ),
    .Y(_0744_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2328_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0207_),
    .B(_0744_),
    .A(_0730_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _2329_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[5] ),
    .B(_0710_),
    .C(_0738_),
    .Y(_0745_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2330_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0745_),
    .A(_0681_),
    .Y(_0746_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2331_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0208_),
    .B(_0746_),
    .A(_0730_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2332_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0747_),
    .B(_0745_),
    .A(_0681_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2333_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0747_),
    .A(_0679_),
    .Y(_0748_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2334_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0209_),
    .B(_0748_),
    .A(_0730_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2335_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0747_),
    .A(_0679_),
    .Y(_0749_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2336_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0749_),
    .A(_0674_),
    .Y(_0750_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2337_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0210_),
    .B(_0750_),
    .A(_0734_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2338_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0749_),
    .A(_0674_),
    .Y(_0751_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2339_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0751_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[9] ),
    .Y(_0752_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2340_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0753_),
    .B(_0751_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2341_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0727_),
    .B(_0752_),
    .C(_0753_),
    .Y(_0754_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2342_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0754_),
    .Y(_0211_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2343_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0752_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[10] ),
    .Y(_0755_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2344_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0212_),
    .B(_0755_),
    .A(_0734_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2345_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0756_),
    .C(\tt_um_rejunity_ay8913.tone_B_generator.counter[11] ),
    .B(_0752_),
    .A(\tt_um_rejunity_ay8913.tone_B_generator.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2346_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0213_),
    .B(_0756_),
    .A(_0734_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2347_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0757_),
    .A(\tt_um_rejunity_ay8913.tone_B ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2348_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0758_),
    .C(_0757_),
    .B(_0725_),
    .A(_0543_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2349_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0492_),
    .A(_0757_),
    .B(_0543_),
    .C(_0725_),
    .Y(_0759_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2350_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0759_),
    .A(_0758_),
    .Y(_0760_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2351_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0760_),
    .Y(_0214_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2352_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0761_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2353_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0762_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2354_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[4] ),
    .A(_0762_),
    .Y(_0763_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2355_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0764_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2356_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[3] ),
    .A(_0764_),
    .Y(_0765_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2357_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[2] ),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[2] ),
    .Y(_0766_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2358_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0766_),
    .A(_0765_),
    .Y(_0767_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2359_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0768_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.period[0] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2360_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0769_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2361_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[0] ),
    .B(_0768_),
    .C(_0769_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.counter[1] ),
    .Y(_0770_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2362_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0769_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[1] ),
    .Y(_0771_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2363_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0772_),
    .B(_0771_),
    .A(_0770_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2364_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0773_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2365_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0764_),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[3] ),
    .C(\tt_um_rejunity_ay8913.tone_A_generator.period[4] ),
    .D(_0762_),
    .Y(_0774_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2366_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0774_),
    .A(_0773_),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[2] ),
    .C(_0765_),
    .Y(_0775_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2367_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0776_),
    .A(_0767_),
    .B(_0772_),
    .C(_0775_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2368_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0761_),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[5] ),
    .C(_0763_),
    .D(_0776_),
    .Y(_0777_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2369_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[5] ),
    .A(_0761_),
    .Y(_0778_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2370_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0779_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2371_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[6] ),
    .A(_0779_),
    .Y(_0780_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2372_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0781_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2373_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0781_),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[7] ),
    .C(\tt_um_rejunity_ay8913.tone_A_generator.period[6] ),
    .D(_0779_),
    .Y(_0782_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2374_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0782_),
    .A(_0777_),
    .B(_0778_),
    .C(_0780_),
    .Y(_0783_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2375_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0784_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2376_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[8] ),
    .A(_0784_),
    .Y(_0785_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2377_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[7] ),
    .A(_0781_),
    .Y(_0786_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2378_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0787_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2379_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0787_),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[9] ),
    .C(\tt_um_rejunity_ay8913.tone_A_generator.period[8] ),
    .D(_0784_),
    .Y(_0788_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2380_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0788_),
    .A(_0783_),
    .B(_0785_),
    .C(_0786_),
    .Y(_0789_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2381_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[9] ),
    .A(_0787_),
    .Y(_0790_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2382_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0791_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.period[10] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2383_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0792_),
    .B(_0791_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2384_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0793_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.period[11] ));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2385_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[11] ),
    .B(_0793_),
    .C(_0791_),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.counter[10] ),
    .Y(_0794_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2386_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0795_),
    .B(_0794_),
    .A(_0792_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2387_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0796_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2388_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0797_),
    .A(_0796_),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[11] ),
    .C(_0792_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2389_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0797_),
    .A(_0789_),
    .B(_0790_),
    .C(_0795_),
    .Y(_0798_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2390_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[0] ),
    .Y(_0799_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2391_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0800_),
    .A(_0799_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2392_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0801_),
    .B(_0771_),
    .A(_0763_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2393_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0802_),
    .C(_0801_),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[0] ),
    .A(_0800_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2394_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0767_),
    .B(_0790_),
    .C(_0795_),
    .D(_0802_),
    .Y(_0803_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2395_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0770_),
    .B(_0774_),
    .C(_0782_),
    .Y(_0804_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2396_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0805_),
    .B(_0780_),
    .A(_0778_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2397_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0806_),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[11] ),
    .A(_0796_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2398_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0807_),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.period[5] ),
    .A(_0761_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2399_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0806_),
    .B(_0807_),
    .C(_0785_),
    .D(_0786_),
    .Y(_0808_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2400_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0788_),
    .B(_0805_),
    .C(_0808_),
    .Y(_0809_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2401_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0810_),
    .B(_0809_),
    .A(_0804_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2402_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0810_),
    .A(_0803_),
    .Y(_0811_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2403_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0812_),
    .A(_0798_),
    .B(_0811_),
    .C(_0417_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2404_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0813_),
    .B(_0812_),
    .A(_1141_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2405_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0813_),
    .Y(_0814_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2406_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0417_),
    .A(_0799_),
    .Y(_0815_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2407_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0815_),
    .A(_0814_),
    .Y(_0816_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2408_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0816_),
    .Y(_0215_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2409_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0813_),
    .Y(_0817_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2410_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[1] ),
    .B(_0799_),
    .C(_0410_),
    .D(_0415_),
    .Y(_0818_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2411_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\tt_um_rejunity_ay8913.tone_A_generator.counter[1] ),
    .A(_0799_),
    .B(_0429_),
    .C(_0430_),
    .Y(_0819_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2412_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0820_),
    .B(_0819_),
    .A(_0818_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2413_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0216_),
    .B(_0820_),
    .A(_0817_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2414_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0813_),
    .Y(_0821_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2415_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0822_),
    .B(_0818_),
    .A(_0773_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2416_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0818_),
    .A(_0773_),
    .Y(_0823_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2417_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0821_),
    .B(_0822_),
    .C(_0823_),
    .Y(_0824_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2418_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0824_),
    .Y(_0217_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2419_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0764_),
    .B(_0773_),
    .C(_0818_),
    .Y(_0825_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2420_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0826_),
    .B(_0822_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2421_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0814_),
    .B(_0825_),
    .C(_0826_),
    .Y(_0827_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2422_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0827_),
    .Y(_0218_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2423_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0825_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[4] ),
    .Y(_0828_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2424_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0829_),
    .B(_0825_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2425_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0814_),
    .B(_0828_),
    .C(_0829_),
    .Y(_0830_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2426_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0830_),
    .Y(_0219_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2427_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0828_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[5] ),
    .Y(_0831_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2428_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0220_),
    .B(_0831_),
    .A(_0817_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _2429_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[5] ),
    .B(\tt_um_rejunity_ay8913.tone_A_generator.counter[4] ),
    .C(_0825_),
    .Y(_0832_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2430_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0832_),
    .A(_0779_),
    .Y(_0833_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2431_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0221_),
    .B(_0833_),
    .A(_0817_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2432_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0834_),
    .B(_0832_),
    .A(_0779_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2433_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0834_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[7] ),
    .Y(_0835_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2434_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0222_),
    .B(_0835_),
    .A(_0817_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2435_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0834_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[7] ),
    .Y(_0836_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2436_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0836_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[8] ),
    .Y(_0837_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2437_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0223_),
    .B(_0837_),
    .A(_0821_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2438_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0836_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[8] ),
    .Y(_0838_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2439_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0838_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[9] ),
    .Y(_0839_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2440_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0840_),
    .B(_0838_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2441_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0814_),
    .B(_0839_),
    .C(_0840_),
    .Y(_0841_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2442_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0841_),
    .Y(_0224_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2443_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0839_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[10] ),
    .Y(_0842_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2444_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0225_),
    .B(_0842_),
    .A(_0821_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2445_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0843_),
    .C(\tt_um_rejunity_ay8913.tone_A_generator.counter[11] ),
    .B(_0839_),
    .A(\tt_um_rejunity_ay8913.tone_A_generator.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2446_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0226_),
    .B(_0843_),
    .A(_0821_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2447_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0812_),
    .A(\tt_um_rejunity_ay8913.tone_A ),
    .Y(_0844_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2448_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0844_),
    .A(_0493_),
    .Y(_0845_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2449_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0845_),
    .Y(_0227_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2450_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0228_),
    .B(_1104_),
    .A(\tt_um_rejunity_ay8913.clk_counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2451_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_ay8913.clk_counter[1] ),
    .A(\tt_um_rejunity_ay8913.clk_counter[0] ),
    .Y(_0846_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2452_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0269_),
    .B(_0408_),
    .C(_0846_),
    .Y(_0847_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2453_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0847_),
    .Y(_0229_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2454_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0848_),
    .B(_0846_),
    .A(\tt_um_rejunity_ay8913.clk_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2455_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0846_),
    .A(\tt_um_rejunity_ay8913.clk_counter[2] ),
    .Y(_0849_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2456_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0269_),
    .B(_0848_),
    .C(_0849_),
    .Y(_0850_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2457_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0850_),
    .Y(_0230_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2458_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0849_),
    .A(\tt_um_rejunity_ay8913.clk_counter[3] ),
    .Y(_0851_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2459_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0849_),
    .A(\tt_um_rejunity_ay8913.clk_counter[3] ),
    .Y(_0852_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2460_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0853_),
    .B(_0852_),
    .A(_1111_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2461_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0231_),
    .B(_0853_),
    .A(_0851_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2462_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0851_),
    .A(\tt_um_rejunity_ay8913.clk_counter[4] ),
    .Y(_0854_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2463_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0851_),
    .A(\tt_um_rejunity_ay8913.clk_counter[4] ),
    .Y(_0855_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2464_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0856_),
    .B(_0855_),
    .A(_1111_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2465_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0232_),
    .B(_0856_),
    .A(_0854_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2466_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0857_),
    .B(_0854_),
    .A(\tt_um_rejunity_ay8913.clk_counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2467_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0854_),
    .A(\tt_um_rejunity_ay8913.clk_counter[5] ),
    .Y(_0858_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2468_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0858_),
    .A(_1110_),
    .Y(_0859_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2469_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0859_),
    .A(_0857_),
    .Y(_0860_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2470_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0860_),
    .Y(_0233_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2471_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0857_),
    .A(\tt_um_rejunity_ay8913.clk_counter[6] ),
    .Y(_0861_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2472_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0861_),
    .A(_0276_),
    .Y(_0862_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2473_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0862_),
    .Y(_0234_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2474_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0863_),
    .B(net8),
    .A(net9));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2475_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net5),
    .A(net6),
    .Y(_0864_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2476_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net7),
    .A(net4),
    .Y(_0865_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2477_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0863_),
    .B(_0864_),
    .C(_0865_),
    .Y(_0866_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2478_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0867_),
    .A(\tt_um_rejunity_ay8913.active ),
    .B(_0863_),
    .C(_0866_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2479_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0867_),
    .A(_0276_),
    .Y(_0868_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2480_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0868_),
    .Y(_0235_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2481_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0866_),
    .Y(_0869_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2482_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0869_),
    .A(_1069_),
    .Y(_0870_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2483_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0871_),
    .A(_1066_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2484_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0866_),
    .Y(_0872_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2485_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0873_),
    .C(_0493_),
    .B(_0872_),
    .A(_0871_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2486_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0873_),
    .A(_0870_),
    .Y(_0874_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2487_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0874_),
    .Y(_0236_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2488_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0869_),
    .A(_1068_),
    .Y(_0875_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2489_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0876_),
    .A(_0663_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2490_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0877_),
    .C(_1103_),
    .B(_0872_),
    .A(_0876_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2491_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0877_),
    .A(_0875_),
    .Y(_0878_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2492_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0878_),
    .Y(_0237_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2493_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0869_),
    .A(\tt_um_rejunity_ay8913.latched_register[2] ),
    .Y(_0879_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2494_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0880_),
    .A(_0665_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2495_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0881_),
    .C(_1103_),
    .B(_0872_),
    .A(_0880_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2496_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0881_),
    .A(_0879_),
    .Y(_0882_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2497_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0882_),
    .Y(_0238_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2498_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0869_),
    .A(\tt_um_rejunity_ay8913.latched_register[3] ),
    .Y(_0883_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2499_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0884_),
    .A(_0667_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2500_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0885_),
    .C(_1103_),
    .B(_0872_),
    .A(_0884_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2501_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0885_),
    .A(_0883_),
    .Y(_0886_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2502_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0886_),
    .Y(_0239_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2503_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0887_),
    .A(\blink.LED ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2504_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0966_),
    .A(_0887_),
    .Y(_0240_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2505_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0279_),
    .A(_1230_),
    .Y(_0888_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2506_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0888_),
    .Y(_0889_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2507_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0890_),
    .B(_0888_),
    .A(_1096_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2508_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0890_),
    .Y(_0891_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2509_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0318_),
    .B(_0889_),
    .C(_0891_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[0] ),
    .Y(_0892_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2510_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0892_),
    .Y(_0241_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2511_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0663_),
    .B(_0889_),
    .C(_0891_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[1] ),
    .Y(_0893_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2512_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0893_),
    .Y(_0242_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2513_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0665_),
    .B(_0889_),
    .C(_0891_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[2] ),
    .Y(_0894_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2514_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0894_),
    .Y(_0243_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2515_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0667_),
    .B(_0889_),
    .C(_0891_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[3] ),
    .Y(_0895_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2516_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0895_),
    .Y(_0244_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2517_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0888_),
    .Y(_0896_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2518_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0890_),
    .Y(_0897_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2519_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0293_),
    .B(_0896_),
    .C(_0897_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[4] ),
    .Y(_0898_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2520_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0898_),
    .Y(_0245_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2521_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net5),
    .B(_0896_),
    .C(_0897_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[5] ),
    .Y(_0899_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2522_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0899_),
    .Y(_0246_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2523_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net6),
    .B(_0896_),
    .C(_0897_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[6] ),
    .Y(_0900_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2524_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0900_),
    .Y(_0247_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2525_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net7),
    .B(_0896_),
    .C(_0897_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.period[7] ),
    .Y(_0901_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2526_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0901_),
    .Y(_0248_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2527_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0279_),
    .A(_1070_),
    .Y(_0902_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2528_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0903_),
    .B(_0902_),
    .A(_1128_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2529_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0318_),
    .B(_0902_),
    .C(_0903_),
    .D(\tt_um_rejunity_ay8913.amplitude_C[0] ),
    .Y(_0904_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2530_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0904_),
    .Y(_0249_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2531_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1090_),
    .B(_0902_),
    .C(_0903_),
    .D(\tt_um_rejunity_ay8913.envelope_C ),
    .Y(_0905_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2532_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0905_),
    .Y(_0250_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2533_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0279_),
    .A(_1093_),
    .Y(_0906_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2534_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0907_),
    .B(_0906_),
    .A(_1097_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2535_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1066_),
    .B(_0906_),
    .C(_0907_),
    .D(\tt_um_rejunity_ay8913.amplitude_B[0] ),
    .Y(_0908_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2536_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0908_),
    .Y(_0251_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2537_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1090_),
    .B(_0906_),
    .C(_0907_),
    .D(\tt_um_rejunity_ay8913.envelope_B ),
    .Y(_0909_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2538_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0909_),
    .Y(_0252_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2539_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0910_),
    .B(_0329_),
    .A(_0492_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2540_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1066_),
    .B(_0137_),
    .C(_0910_),
    .D(\tt_um_rejunity_ay8913.envelope_generator.hold ),
    .Y(_0911_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2541_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0911_),
    .Y(_0253_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2542_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0663_),
    .B(_0137_),
    .C(_0910_),
    .D(\tt_um_rejunity_ay8913.envelope_alternate ),
    .Y(_0912_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2543_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0912_),
    .Y(_0254_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2544_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0665_),
    .B(_0137_),
    .C(_0910_),
    .D(\tt_um_rejunity_ay8913.envelope_attack ),
    .Y(_0913_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2545_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0913_),
    .Y(_0255_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2546_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0667_),
    .B(_0329_),
    .C(_0910_),
    .D(\tt_um_rejunity_ay8913.envelope_continue ),
    .Y(_0914_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2547_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0914_),
    .Y(_0256_));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2548_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_6_wb_clk_i),
    .D(_0000_),
    .Q(\blink.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2549_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_6_wb_clk_i),
    .D(_0001_),
    .Q(\blink.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2550_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_5_wb_clk_i),
    .D(_0002_),
    .Q(\blink.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2551_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_7_wb_clk_i),
    .D(_0003_),
    .Q(\blink.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2552_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_6_wb_clk_i),
    .D(_0004_),
    .Q(\blink.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2553_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_6_wb_clk_i),
    .D(_0005_),
    .Q(\blink.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2554_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_2_wb_clk_i),
    .D(_0006_),
    .Q(\blink.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2555_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_1_wb_clk_i),
    .D(_0007_),
    .Q(\blink.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2556_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_2_wb_clk_i),
    .D(_0008_),
    .Q(\blink.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2557_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_1_wb_clk_i),
    .D(_0009_),
    .Q(\blink.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2558_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_1_wb_clk_i),
    .D(_0010_),
    .Q(\blink.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2559_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_2_wb_clk_i),
    .D(_0011_),
    .Q(\blink.counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2560_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_1_wb_clk_i),
    .D(_0012_),
    .Q(\blink.counter[12] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2561_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_1_wb_clk_i),
    .D(_0013_),
    .Q(\blink.counter[13] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2562_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_1_wb_clk_i),
    .D(_0014_),
    .Q(\blink.counter[14] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2563_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_43_wb_clk_i),
    .D(_0015_),
    .Q(\blink.counter[15] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2564_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_0_wb_clk_i),
    .D(_0016_),
    .Q(\blink.counter[16] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2565_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_0_wb_clk_i),
    .D(_0017_),
    .Q(\blink.counter[17] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2566_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_43_wb_clk_i),
    .D(_0018_),
    .Q(\blink.counter[18] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2567_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_43_wb_clk_i),
    .D(_0019_),
    .Q(\blink.counter[19] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2568_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_0_wb_clk_i),
    .D(_0020_),
    .Q(\blink.counter[20] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2569_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_40_wb_clk_i),
    .D(_0021_),
    .Q(\blink.counter[21] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2570_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_43_wb_clk_i),
    .D(_0022_),
    .Q(\blink.counter[22] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2571_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_43_wb_clk_i),
    .D(_0023_),
    .Q(\blink.counter[23] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2572_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_43_wb_clk_i),
    .D(_0024_),
    .Q(\blink.counter[24] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2573_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_42_wb_clk_i),
    .D(_0025_),
    .Q(\blink.counter[25] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2574_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_42_wb_clk_i),
    .D(_0026_),
    .Q(\blink.counter[26] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2575_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_42_wb_clk_i),
    .D(_0027_),
    .Q(\blink.counter[27] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2576_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_42_wb_clk_i),
    .D(_0028_),
    .Q(\blink.counter[28] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2577_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_42_wb_clk_i),
    .D(_0029_),
    .Q(\blink.counter[29] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2578_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_41_wb_clk_i),
    .D(_0030_),
    .Q(\blink.counter[30] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2579_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_41_wb_clk_i),
    .D(_0031_),
    .Q(\blink.counter[31] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2580_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_3_wb_clk_i),
    .D(_0032_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.period[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2581_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_2_wb_clk_i),
    .D(_0033_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2582_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_3_wb_clk_i),
    .D(_0034_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.period[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2583_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_3_wb_clk_i),
    .D(_0035_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.period[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2584_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_37_wb_clk_i),
    .D(_0036_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.period[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2585_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_7_wb_clk_i),
    .D(_0037_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2586_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_7_wb_clk_i),
    .D(_0038_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2587_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_7_wb_clk_i),
    .D(_0039_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2588_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_7_wb_clk_i),
    .D(_0040_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2589_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_34_wb_clk_i),
    .D(_0041_),
    .Q(\tt_um_rejunity_ay8913.pwm_master.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2590_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_31_wb_clk_i),
    .D(_0042_),
    .Q(\tt_um_rejunity_ay8913.pwm_master.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2591_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_33_wb_clk_i),
    .D(_0043_),
    .Q(\tt_um_rejunity_ay8913.pwm_master.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2592_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_30_wb_clk_i),
    .D(_0044_),
    .Q(\tt_um_rejunity_ay8913.pwm_master.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2593_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_33_wb_clk_i),
    .D(_0045_),
    .Q(\tt_um_rejunity_ay8913.pwm_master.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2594_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_33_wb_clk_i),
    .D(_0046_),
    .Q(\tt_um_rejunity_ay8913.pwm_master.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2595_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_34_wb_clk_i),
    .D(_0047_),
    .Q(\tt_um_rejunity_ay8913.pwm_master.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2596_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_34_wb_clk_i),
    .D(_0048_),
    .Q(\tt_um_rejunity_ay8913.pwm_master.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2597_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_34_wb_clk_i),
    .D(_0049_),
    .Q(\tt_um_rejunity_ay8913.pwm_master.accumulator[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2598_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_32_wb_clk_i),
    .D(_0050_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2599_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_32_wb_clk_i),
    .D(_0051_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2600_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_31_wb_clk_i),
    .D(_0052_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2601_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_32_wb_clk_i),
    .D(_0053_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2602_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_31_wb_clk_i),
    .D(_0054_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2603_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_31_wb_clk_i),
    .D(_0055_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2604_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_31_wb_clk_i),
    .D(_0056_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2605_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_31_wb_clk_i),
    .D(_0057_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2606_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_31_wb_clk_i),
    .D(_0058_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2607_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_30_wb_clk_i),
    .D(_0059_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2608_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_35_wb_clk_i),
    .D(_0060_),
    .Q(\tt_um_rejunity_ay8913.pwm_C.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2609_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_34_wb_clk_i),
    .D(_0061_),
    .Q(\tt_um_rejunity_ay8913.pwm_C.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2610_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_34_wb_clk_i),
    .D(_0062_),
    .Q(\tt_um_rejunity_ay8913.pwm_C.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2611_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_40_wb_clk_i),
    .D(_0063_),
    .Q(\tt_um_rejunity_ay8913.pwm_C.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2612_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_40_wb_clk_i),
    .D(_0064_),
    .Q(\tt_um_rejunity_ay8913.pwm_C.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2613_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_40_wb_clk_i),
    .D(_0065_),
    .Q(\tt_um_rejunity_ay8913.pwm_C.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2614_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_40_wb_clk_i),
    .D(_0066_),
    .Q(\tt_um_rejunity_ay8913.pwm_C.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2615_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_39_wb_clk_i),
    .D(_0067_),
    .Q(\tt_um_rejunity_ay8913.pwm_C.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2616_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_36_wb_clk_i),
    .D(_0068_),
    .Q(\tt_um_rejunity_ay8913.pwm_B.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2617_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_36_wb_clk_i),
    .D(_0069_),
    .Q(\tt_um_rejunity_ay8913.pwm_B.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2618_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_35_wb_clk_i),
    .D(_0070_),
    .Q(\tt_um_rejunity_ay8913.pwm_B.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2619_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_35_wb_clk_i),
    .D(_0071_),
    .Q(\tt_um_rejunity_ay8913.pwm_B.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2620_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_35_wb_clk_i),
    .D(_0072_),
    .Q(\tt_um_rejunity_ay8913.pwm_B.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2621_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_39_wb_clk_i),
    .D(_0073_),
    .Q(\tt_um_rejunity_ay8913.pwm_B.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2622_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_39_wb_clk_i),
    .D(_0074_),
    .Q(\tt_um_rejunity_ay8913.pwm_B.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2623_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_34_wb_clk_i),
    .D(_0075_),
    .Q(\tt_um_rejunity_ay8913.pwm_B.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2624_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_5_wb_clk_i),
    .D(_0076_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2625_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_13_wb_clk_i),
    .D(_0077_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2626_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_8_wb_clk_i),
    .D(_0078_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2627_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_7_wb_clk_i),
    .D(_0079_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2628_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_12_wb_clk_i),
    .D(_0080_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2629_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_11_wb_clk_i),
    .D(_0081_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2630_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_11_wb_clk_i),
    .D(_0082_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2631_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_10_wb_clk_i),
    .D(_0083_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.period[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2632_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_4_wb_clk_i),
    .D(_0084_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2633_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_2_wb_clk_i),
    .D(_0085_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2634_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_2_wb_clk_i),
    .D(_0086_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2635_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_2_wb_clk_i),
    .D(_0087_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2636_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_14_wb_clk_i),
    .D(_0088_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2637_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_13_wb_clk_i),
    .D(_0089_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2638_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_25_wb_clk_i),
    .D(_0090_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2639_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_14_wb_clk_i),
    .D(_0091_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2640_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_13_wb_clk_i),
    .D(_0092_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2641_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_13_wb_clk_i),
    .D(_0093_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2642_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_14_wb_clk_i),
    .D(_0094_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2643_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_14_wb_clk_i),
    .D(_0095_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.period[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2644_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_30_wb_clk_i),
    .D(_0096_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2645_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_30_wb_clk_i),
    .D(_0097_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2646_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_30_wb_clk_i),
    .D(_0098_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2647_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_29_wb_clk_i),
    .D(_0099_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2648_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_29_wb_clk_i),
    .D(_0100_),
    .Q(\tt_um_rejunity_ay8913.spi_dac_i_2.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2649_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_35_wb_clk_i),
    .D(_0101_),
    .Q(\tt_um_rejunity_ay8913.pwm_A.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2650_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_35_wb_clk_i),
    .D(_0102_),
    .Q(\tt_um_rejunity_ay8913.pwm_A.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2651_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_35_wb_clk_i),
    .D(_0103_),
    .Q(\tt_um_rejunity_ay8913.pwm_A.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2652_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_33_wb_clk_i),
    .D(_0104_),
    .Q(\tt_um_rejunity_ay8913.pwm_A.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2653_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_36_wb_clk_i),
    .D(_0105_),
    .Q(\tt_um_rejunity_ay8913.pwm_A.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2654_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_26_wb_clk_i),
    .D(_0106_),
    .Q(\tt_um_rejunity_ay8913.pwm_A.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2655_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_29_wb_clk_i),
    .D(_0107_),
    .Q(\tt_um_rejunity_ay8913.pwm_A.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2656_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_34_wb_clk_i),
    .D(_0108_),
    .Q(\tt_um_rejunity_ay8913.pwm_A.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2657_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_37_wb_clk_i),
    .D(_0109_),
    .Q(\tt_um_rejunity_ay8913.amplitude_A[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2658_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_36_wb_clk_i),
    .D(_0110_),
    .Q(\tt_um_rejunity_ay8913.envelope_A ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2659_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_18_wb_clk_i),
    .D(_0111_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2660_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_18_wb_clk_i),
    .D(_0112_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2661_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_18_wb_clk_i),
    .D(_0113_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2662_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_18_wb_clk_i),
    .D(_0114_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2663_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_17_wb_clk_i),
    .D(_0115_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[12] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2664_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_19_wb_clk_i),
    .D(_0116_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[13] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2665_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_18_wb_clk_i),
    .D(_0117_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[14] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2666_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_18_wb_clk_i),
    .D(_0118_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[15] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2667_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_14_wb_clk_i),
    .D(_0119_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2668_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_15_wb_clk_i),
    .D(_0120_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2669_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_14_wb_clk_i),
    .D(_0121_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2670_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_13_wb_clk_i),
    .D(_0122_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2671_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_18_wb_clk_i),
    .D(_0123_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2672_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_18_wb_clk_i),
    .D(_0124_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2673_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_16_wb_clk_i),
    .D(_0125_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2674_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_11_wb_clk_i),
    .D(_0126_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2675_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_34_wb_clk_i),
    .D(_0127_),
    .Q(\tt_um_rejunity_ay8913.DAC_le ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2676_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_30_wb_clk_i),
    .D(_0128_),
    .Q(\tt_um_rejunity_ay8913.DAC_dat ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2677_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_32_wb_clk_i),
    .D(_0129_),
    .Q(\tt_um_rejunity_ay8913.DAC_clk ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2678_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_37_wb_clk_i),
    .D(_0130_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0 ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2679_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_26_wb_clk_i),
    .D(_0131_),
    .Q(\tt_um_rejunity_ay8913.tone_disable_A ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2680_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_37_wb_clk_i),
    .D(_0132_),
    .Q(\tt_um_rejunity_ay8913.tone_disable_B ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2681_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_37_wb_clk_i),
    .D(_0133_),
    .Q(\tt_um_rejunity_ay8913.tone_disable_C ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2682_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_25_wb_clk_i),
    .D(_0134_),
    .Q(\tt_um_rejunity_ay8913.noise_disable_A ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2683_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_26_wb_clk_i),
    .D(_0135_),
    .Q(\tt_um_rejunity_ay8913.noise_disable_B ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2684_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0136_),
    .Q(\tt_um_rejunity_ay8913.noise_disable_C ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2685_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0137_),
    .Q(\tt_um_rejunity_ay8913.restart_envelope ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2686_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_28_wb_clk_i),
    .D(_0138_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2687_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_28_wb_clk_i),
    .D(_0139_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2688_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0140_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2689_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_28_wb_clk_i),
    .D(_0141_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.envelope_counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2690_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_23_wb_clk_i),
    .D(_0142_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.stop ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2691_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_22_wb_clk_i),
    .D(_0143_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2692_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_15_wb_clk_i),
    .D(_0144_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2693_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_24_wb_clk_i),
    .D(_0145_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2694_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_24_wb_clk_i),
    .D(_0146_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2695_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_21_wb_clk_i),
    .D(_0147_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2696_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_22_wb_clk_i),
    .D(_0148_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2697_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_22_wb_clk_i),
    .D(_0149_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2698_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_21_wb_clk_i),
    .D(_0150_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2699_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_20_wb_clk_i),
    .D(_0151_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2700_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_21_wb_clk_i),
    .D(_0152_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2701_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_19_wb_clk_i),
    .D(_0153_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2702_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_19_wb_clk_i),
    .D(_0154_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2703_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_19_wb_clk_i),
    .D(_0155_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2704_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_19_wb_clk_i),
    .D(_0156_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[12] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2705_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_20_wb_clk_i),
    .D(_0157_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[13] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2706_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_20_wb_clk_i),
    .D(_0158_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[14] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2707_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_20_wb_clk_i),
    .D(_0159_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.tone.counter[15] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2708_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0160_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.invert_output ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2709_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_36_wb_clk_i),
    .D(_0161_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2710_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_36_wb_clk_i),
    .D(_0162_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2711_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_35_wb_clk_i),
    .D(_0163_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2712_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_38_wb_clk_i),
    .D(_0164_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2713_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_38_wb_clk_i),
    .D(_0165_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2714_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_38_wb_clk_i),
    .D(_0166_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2715_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_3_wb_clk_i),
    .D(_0167_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2716_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_0_wb_clk_i),
    .D(_0168_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2717_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_41_wb_clk_i),
    .D(_0169_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2718_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_41_wb_clk_i),
    .D(_0170_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2719_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_40_wb_clk_i),
    .D(_0171_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2720_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_40_wb_clk_i),
    .D(_0172_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2721_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_40_wb_clk_i),
    .D(_0173_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[12] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2722_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_39_wb_clk_i),
    .D(_0174_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[13] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2723_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_39_wb_clk_i),
    .D(_0175_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[14] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2724_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_39_wb_clk_i),
    .D(_0176_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[15] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2725_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_38_wb_clk_i),
    .D(_0177_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.lfsr[16] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2726_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_37_wb_clk_i),
    .D(_0178_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.signal_edge.signal ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2727_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_4_wb_clk_i),
    .D(_0179_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.tone.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2728_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_3_wb_clk_i),
    .D(_0180_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.tone.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2729_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_0_wb_clk_i),
    .D(_0181_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.tone.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2730_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_3_wb_clk_i),
    .D(_0182_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.tone.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2731_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_3_wb_clk_i),
    .D(_0183_),
    .Q(\tt_um_rejunity_ay8913.noise_generator.tone.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2732_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_22_wb_clk_i),
    .D(_0184_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0 ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2733_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_10_wb_clk_i),
    .D(_0185_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2734_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_12_wb_clk_i),
    .D(_0186_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2735_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_9_wb_clk_i),
    .D(_0187_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2736_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_9_wb_clk_i),
    .D(_0188_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2737_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_9_wb_clk_i),
    .D(_0189_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2738_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_10_wb_clk_i),
    .D(_0190_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2739_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_10_wb_clk_i),
    .D(_0191_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2740_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_10_wb_clk_i),
    .D(_0192_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2741_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_8_wb_clk_i),
    .D(_0193_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2742_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_8_wb_clk_i),
    .D(_0194_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2743_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_8_wb_clk_i),
    .D(_0195_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2744_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_8_wb_clk_i),
    .D(_0196_),
    .Q(\tt_um_rejunity_ay8913.tone_C_generator.counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2745_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_4_wb_clk_i),
    .D(_0197_),
    .Q(\tt_um_rejunity_ay8913.tone_C ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2746_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_14_wb_clk_i),
    .D(_0198_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2747_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_14_wb_clk_i),
    .D(_0199_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2748_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_24_wb_clk_i),
    .D(_0200_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2749_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_24_wb_clk_i),
    .D(_0201_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.period[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2750_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_5_wb_clk_i),
    .D(_0202_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2751_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_13_wb_clk_i),
    .D(_0203_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2752_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_4_wb_clk_i),
    .D(_0204_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2753_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_4_wb_clk_i),
    .D(_0205_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2754_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_5_wb_clk_i),
    .D(_0206_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2755_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_5_wb_clk_i),
    .D(_0207_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2756_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_5_wb_clk_i),
    .D(_0208_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2757_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_5_wb_clk_i),
    .D(_0209_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2758_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_6_wb_clk_i),
    .D(_0210_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2759_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_5_wb_clk_i),
    .D(_0211_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2760_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_6_wb_clk_i),
    .D(_0212_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2761_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_6_wb_clk_i),
    .D(_0213_),
    .Q(\tt_um_rejunity_ay8913.tone_B_generator.counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2762_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_4_wb_clk_i),
    .D(_0214_),
    .Q(\tt_um_rejunity_ay8913.tone_B ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2763_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_16_wb_clk_i),
    .D(_0215_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2764_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_12_wb_clk_i),
    .D(_0216_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2765_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_12_wb_clk_i),
    .D(_0217_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2766_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_12_wb_clk_i),
    .D(_0218_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2767_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_11_wb_clk_i),
    .D(_0219_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2768_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_11_wb_clk_i),
    .D(_0220_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2769_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_11_wb_clk_i),
    .D(_0221_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2770_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_11_wb_clk_i),
    .D(_0222_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2771_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_17_wb_clk_i),
    .D(_0223_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2772_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_17_wb_clk_i),
    .D(_0224_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2773_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_17_wb_clk_i),
    .D(_0225_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2774_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_17_wb_clk_i),
    .D(_0226_),
    .Q(\tt_um_rejunity_ay8913.tone_A_generator.counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2775_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_25_wb_clk_i),
    .D(_0227_),
    .Q(\tt_um_rejunity_ay8913.tone_A ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2776_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_26_wb_clk_i),
    .D(_0228_),
    .Q(\tt_um_rejunity_ay8913.clk_counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2777_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0229_),
    .Q(\tt_um_rejunity_ay8913.clk_counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2778_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_26_wb_clk_i),
    .D(_0230_),
    .Q(\tt_um_rejunity_ay8913.clk_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2779_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_29_wb_clk_i),
    .D(_0231_),
    .Q(\tt_um_rejunity_ay8913.clk_counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2780_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_29_wb_clk_i),
    .D(_0232_),
    .Q(\tt_um_rejunity_ay8913.clk_counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2781_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_28_wb_clk_i),
    .D(_0233_),
    .Q(\tt_um_rejunity_ay8913.clk_counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2782_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0234_),
    .Q(\tt_um_rejunity_ay8913.clk_counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2783_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_23_wb_clk_i),
    .D(_0235_),
    .Q(\tt_um_rejunity_ay8913.active ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2784_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_25_wb_clk_i),
    .D(_0236_),
    .Q(\tt_um_rejunity_ay8913.latched_register[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2785_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_14_wb_clk_i),
    .D(_0237_),
    .Q(\tt_um_rejunity_ay8913.latched_register[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2786_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0238_),
    .Q(\tt_um_rejunity_ay8913.latched_register[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2787_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_23_wb_clk_i),
    .D(_0239_),
    .Q(\tt_um_rejunity_ay8913.latched_register[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2788_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_41_wb_clk_i),
    .D(_0240_),
    .Q(\blink.LED ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2789_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_24_wb_clk_i),
    .D(_0241_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2790_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_24_wb_clk_i),
    .D(_0242_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2791_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_23_wb_clk_i),
    .D(_0243_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2792_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_23_wb_clk_i),
    .D(_0244_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2793_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_23_wb_clk_i),
    .D(_0245_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2794_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_22_wb_clk_i),
    .D(_0246_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2795_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_22_wb_clk_i),
    .D(_0247_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2796_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_23_wb_clk_i),
    .D(_0248_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.period[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2797_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_26_wb_clk_i),
    .D(_0249_),
    .Q(\tt_um_rejunity_ay8913.amplitude_C[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2798_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_26_wb_clk_i),
    .D(_0250_),
    .Q(\tt_um_rejunity_ay8913.envelope_C ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2799_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_37_wb_clk_i),
    .D(_0251_),
    .Q(\tt_um_rejunity_ay8913.amplitude_B[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2800_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_37_wb_clk_i),
    .D(_0252_),
    .Q(\tt_um_rejunity_ay8913.envelope_B ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2801_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0253_),
    .Q(\tt_um_rejunity_ay8913.envelope_generator.hold ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2802_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0254_),
    .Q(\tt_um_rejunity_ay8913.envelope_alternate ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2803_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_27_wb_clk_i),
    .D(_0255_),
    .Q(\tt_um_rejunity_ay8913.envelope_attack ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2804_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_leaf_23_wb_clk_i),
    .D(_0256_),
    .Q(\tt_um_rejunity_ay8913.envelope_continue ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2824_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.DAC_dat ),
    .Y(net13));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2825_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.DAC_le ),
    .Y(net14));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2826_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_ay8913.DAC_clk ),
    .Y(net15));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(wb_clk_i),
    .Y(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_2_0__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_2_1__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_2_2__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_2_3__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_10_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i),
    .Y(clknet_leaf_10_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_11_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i),
    .Y(clknet_leaf_11_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_12_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i),
    .Y(clknet_leaf_12_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_13_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i),
    .Y(clknet_leaf_13_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_14_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_14_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_15_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_15_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_16_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_16_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_17_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_17_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_18_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_18_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_19_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_19_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_1_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_1_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_20_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_20_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_21_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_21_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_22_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_22_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_23_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_23_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_24_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i),
    .Y(clknet_leaf_24_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_25_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_25_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_26_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_26_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_27_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_27_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_28_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_28_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_29_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_29_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_2_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_2_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_30_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_30_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_31_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_31_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_32_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_32_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_33_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_33_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_34_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_34_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_35_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_35_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_36_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_2__leaf_wb_clk_i),
    .Y(clknet_leaf_36_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_37_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_37_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_38_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_38_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_39_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_39_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_3_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_3_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_40_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_40_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_41_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_41_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_42_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_42_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_43_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_43_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_4_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i),
    .Y(clknet_leaf_4_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_5_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i),
    .Y(clknet_leaf_5_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_6_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i),
    .Y(clknet_leaf_6_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_7_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i),
    .Y(clknet_leaf_7_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_8_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i),
    .Y(clknet_leaf_8_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_leaf_9_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i),
    .Y(clknet_leaf_9_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload0 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkload1 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_42_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_43_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 clkload12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_6_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_7_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_8_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_9_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_10_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 clkload17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_11_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_12_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_13_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_25_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_26_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_28_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_29_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkload24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_30_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_31_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_32_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_33_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 clkload28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_34_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_35_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload3 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_1_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkload30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_36_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_15_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_16_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkload33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_17_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 clkload34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_18_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkload35 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_19_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_20_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_21_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_22_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 clkload39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_23_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 clkload4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_2_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_24_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 clkload5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_3_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_4_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkload7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_38_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_39_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_leaf_41_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input1 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[0]),
    .Y(net1));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(rst_n),
    .Y(net10));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[1]),
    .Y(net2));
 gf180mcu_as_sc_mcu7t3v3__buff_4 input3 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[3]),
    .Y(net3));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[4]),
    .Y(net4));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[5]),
    .Y(net5));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[6]),
    .Y(net6));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[7]),
    .Y(net7));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_2[0]),
    .Y(net8));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_2[1]),
    .Y(net9));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net11),
    .Y(io_out[10]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net12),
    .Y(io_out[11]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net13),
    .Y(io_out[17]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net14),
    .Y(io_out[18]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net15),
    .Y(io_out[19]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net16),
    .Y(io_out[20]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net17),
    .Y(io_out[21]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net18),
    .Y(io_out[8]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net19),
    .Y(io_out[9]));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net20));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net21));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net22));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net23));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net24));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net25));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net26));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net27));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net28));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net29));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net30));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net31));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net32));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net33));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net34));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_35 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net35));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net36));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net37));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_ay8913_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net38));
 assign io_out[0] = net20;
 assign io_out[12] = net28;
 assign io_out[13] = net29;
 assign io_out[14] = net30;
 assign io_out[15] = net31;
 assign io_out[16] = net32;
 assign io_out[1] = net21;
 assign io_out[22] = net38;
 assign io_out[23] = net33;
 assign io_out[24] = net34;
 assign io_out[25] = net35;
 assign io_out[26] = net36;
 assign io_out[27] = net37;
 assign io_out[2] = net22;
 assign io_out[3] = net23;
 assign io_out[4] = net24;
 assign io_out[5] = net25;
 assign io_out[6] = net26;
 assign io_out[7] = net27;
endmodule
