* NGSPICE file created from wrapped_sn76489.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

.subckt wrapped_sn76489 custom_settings[0] custom_settings[1] io_in_1[0] io_in_1[1]
+ io_in_1[2] io_in_1[3] io_in_1[4] io_in_1[5] io_in_1[6] io_in_1[7] io_in_2 io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[17] io_out[18] io_out[19] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i io_out[15] io_out[14]
+ io_out[13] io_out[3] io_out[2] io_out[1] io_out[16]
X_2037_ _0328_ _0329_ _0331_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1343__B _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2106_ _0373_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2084__B _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer7 _0820_ net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1270_ _0715_ _0716_ _0718_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2655_ _0129_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1606_ _1048_ _1049_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_22_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1537_ _0951_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1468_ _0916_ _0911_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1399_ _0839_ _0847_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2586_ _0060_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1978__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2672__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2079__B _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1666__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\] _0648_ _0646_ _0649_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2371_ _0599_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1322_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _0771_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__1672__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1409__A1 _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2569_ _0043_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2545__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2707_ _0181_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2638_ _0112_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2695__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1887__A1 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1871_ _0194_ _0202_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2568__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1940_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\] _0252_ _0255_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2119__A2 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2423_ _1104_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2285_ tt_um_rejunity_sn76489.pwm.accumulator\[4\] net19 _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2354_ _0587_ _0137_ _0588_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1305_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\] _0754_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2447__B _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2710__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2070_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\] _0358_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
+ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_44_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1785_ _1195_ _1197_ _1157_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1854_ _1252_ _1253_ _1254_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1260__A2 _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\] _0238_ _0243_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2406_ _0614_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2276__A1 _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2268_ tt_um_rejunity_sn76489.pwm.accumulator\[2\] _0521_ _0522_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2337_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\] tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\]
+ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\] _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2199_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\] _0465_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
+ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1315__A3 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2200__A1 _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1570_ _1006_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2606__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2053_ _0343_ _0344_ _0330_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xrebuffer17 _0898_ net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2122_ _0280_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1768_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\] _0818_ _1183_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1837_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\] _0892_ _1240_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1906_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\] tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
+ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\] _0952_ tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
+ tt_um_rejunity_sn76489.control_noise\[0\]\[1\] _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__2430__A1 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2497__A1 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1699_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\] _1122_ _1127_ _1128_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2249__A1 _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2629__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput20 net20 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2488__A1 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1622_ _1063_ _1064_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2671_ _0145_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1553_ _0997_ _0998_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1484_ _0909_ _0910_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2479__A1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2036_ _0328_ _0329_ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2105_ _0388_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2403__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer8 _0779_ net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2654_ _0128_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1536_ _0976_ _0979_ _0981_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1605_ _0960_ _0844_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2585_ _0059_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1467_ _0830_ _0912_ _0915_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1398_ _0840_ net50 _0843_ _0844_ _0846_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_54_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2019_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\] _0869_ _0316_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2526__D _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2114__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2370_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\] _0596_ _0593_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\]
+ _0597_ net22 _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1321_ _0767_ _0769_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_19_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2706_ _0180_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_2568_ _0042_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1345__B2 _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1519_ _0963_ _0936_ _0835_ _0965_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2637_ _0111_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2499_ _0690_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1870_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\] _1026_ _0201_ _0202_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_36_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2353_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\] _0000_ _0132_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\]
+ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2422_ _0634_ _0629_ _0636_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2284_ _0533_ _0535_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1304_ _0750_ _0751_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__2055__A2 _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2662__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1999_ _0299_ _0296_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\] _0301_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1557__A1 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1922_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\] _0241_ _0242_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2535__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1784_ _1196_ _1032_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1853_ _1252_ _1253_ _1238_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2685__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2336_ _0575_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\] tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\]
+ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2405_ _0622_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2267_ _0824_ _0864_ _0821_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2198_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
+ _0463_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_35_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2193__B _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2558__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2122__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2052_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\] _1018_ _0344_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xrebuffer18 _0847_ net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2121_ _0365_ _0398_ _0401_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1905_ _0220_ _0227_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1767_ _1171_ _1182_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1698_ _1126_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1836_ _1236_ _1237_ _1239_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2319_ _0560_ _0563_ _0564_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2700__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input11_I io_in_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput21 net21 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1621_ _1046_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2670_ _0144_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1552_ _0966_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1483_ _0928_ _0930_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2104_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\] _0384_ _0386_ _0387_ _0377_
+ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA_input3_I io_in_1[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2035_ _0209_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1819_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\] _1051_ _1224_ _1226_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1914__A1 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer9 _0848_ net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_8_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2653_ _0127_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1535_ _0971_ _0975_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1604_ _0777_ _0815_ _0781_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_22_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2584_ _0058_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1466_ _0913_ _0914_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2321__A1 _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1397_ _0840_ _0841_ _0845_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_49_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2018_ _1210_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_19_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1320_ _0768_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_11_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _0179_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2636_ _0110_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2567_ _0041_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1449_ _0867_ _0896_ _0897_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1518_ _0964_ _0936_ _0825_ _0963_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2498_ _0690_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_25_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2283_ _0224_ net56 _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2352_ net47 _0515_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2524__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2421_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\] _0635_ _0624_ _0636_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1303_ tt_um_rejunity_sn76489.chan\[0\].attenuation.in _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_51_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2035__I _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1998_ _0299_ _0296_ _0300_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2619_ _0093_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2506__A1 _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1852_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\] _1028_ _1253_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1921_ _0231_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1783_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[4\] _1196_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_24_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2335_ _0575_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\] _0576_ _0133_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2266_ _0513_ _0518_ _0519_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2404_ net8 _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2197_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
+ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
+ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_35_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1728__B _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2120_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\] _0389_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
+ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2051_ _0341_ _0342_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2652__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer19 _0782_ net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1835_ _1236_ _1237_ _1238_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1904_ tt_um_rejunity_sn76489.clk_counter\[6\] _0225_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1766_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\] _0818_ _1181_ _1182_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1697_ _1097_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2194__A2 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2318_ tt_um_rejunity_sn76489.pwm.accumulator\[9\] net24 _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2249_ _0286_ _0492_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_33_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2185__A2 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput22 net22 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2675__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1696__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1620_ _1045_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2289__B _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1551_ _0962_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1482_ _0735_ _0929_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2103_ _0380_ _0385_ _0381_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1687__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2034_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\] _0973_ _0329_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1439__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ _1211_ _1225_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2548__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1749_ _1165_ _1167_ _1168_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2218__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1841__A1 _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2652_ _0126_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1534_ _0980_ net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1603_ _1045_ _1046_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1465_ _0889_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2583_ _0057_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2017_ _0312_ _0313_ _0314_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1396_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _0754_ _0756_ _0845_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_13_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2713__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2379__A2 _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_36_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1697__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2704_ _0178_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2635_ _0109_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2566_ _0040_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1448_ _0872_ _0895_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1517_ _0780_ _0833_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2497_ _0655_ _0689_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1379_ _0808_ _0810_ _0826_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2297__A1 _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2609__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2420_ _0628_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2282_ _0530_ _0532_ _0531_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2351_ _0586_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1302_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _0751_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_1997_ _0299_ _0296_ _0210_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2549_ _0023_ clknet_4_7_0_wb_clk_i net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_30_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2618_ _0092_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1851_ _1247_ _1031_ _1251_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1920_ _0236_ _0239_ _0240_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1782_ _1191_ _1193_ _1194_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2581__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2403_ _0620_ _0612_ _0621_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2334_ _0575_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\] _1077_ _0223_ _0576_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2265_ tt_um_rejunity_sn76489.pwm.accumulator\[1\] _0516_ _0519_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2196_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
+ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
+ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2050_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\] _1015_ _0338_ _0342_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2415__A1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1765_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\] _1179_ _1181_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1834_ _1126_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1903_ _0222_ _0226_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1696_ _1102_ _1121_ _1125_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2317_ tt_um_rejunity_sn76489.pwm.accumulator\[8\] net23 _1062_ tt_um_rejunity_sn76489.pwm.accumulator\[9\]
+ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2179_ _0396_ _0449_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2248_ _0504_ _0506_ _1132_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput23 net23 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ _0992_ _0995_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1481_ _0850_ _0906_ _0747_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_1_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2033_ _0323_ _0924_ _0327_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_27_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2102_ _0380_ _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1817_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\] _1051_ _1224_ _1225_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1748_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\] _1014_ _1168_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1679_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\] _1112_ _1099_ _1114_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2642__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2651_ _0125_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1602_ _0953_ _0721_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2582_ _0056_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_14_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1533_ _0976_ _0979_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1464_ _0885_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1395_ _0760_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_54_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2016_ _0312_ _0313_ _0210_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1379__B _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1520__A1 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2538__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2565_ _0039_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1516_ _0813_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2703_ _0177_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2634_ _0108_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1447_ _0872_ _0895_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1378_ _0808_ _0810_ _0826_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_4_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2477__C _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2496_ _0627_ _0669_ _0679_ _0668_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_45_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2350_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\] _0000_ _0511_ _0585_
+ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2281_ _0530_ _0531_ _0532_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1301_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\] _0750_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_30_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1996_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\] _0299_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2548_ _0022_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2617_ _0091_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2479_ _0634_ _0672_ _0677_ _0676_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1781_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\] _0913_ _1194_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1850_ _1246_ _1250_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2333_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\] _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2402_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\] _0617_ _0615_ _0621_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2264_ tt_um_rejunity_sn76489.pwm.accumulator\[1\] _0516_ _0518_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2195_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\] _0403_ _0462_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ _0276_ _0277_ _0284_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2121__A1 _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2188__A1 _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1760__B _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1902_ _0224_ _0225_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\] _1179_ _1180_ _0024_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1833_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\] _0892_ _1237_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2179__A1 _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2316_ _0558_ _0561_ _0562_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1654__C _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1695_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\] _1122_ _1115_ _1125_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2178_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] _0444_ _0448_ _0449_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2247_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\] _0396_ _0505_ _0506_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2006__B _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput13 net13 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput24 net24 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2571__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1480_ _0719_ _0927_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2032_ _0322_ _0326_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1439__A3 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2101_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\] _0373_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
+ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1816_ _1219_ _1055_ _1223_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1747_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\] _1014_ _1167_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1375__A2 _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1678_ _1107_ _1111_ _1113_ _1093_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2594__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2650_ _0124_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1532_ _0922_ _0977_ _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1601_ _0797_ _0851_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2581_ _0055_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input1_I custom_settings[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1463_ _0891_ net58 net52 _0889_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1394_ _0750_ _0804_ _0842_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_2015_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\] _0869_ _0313_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2702_ _0176_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2564_ _0038_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1515_ _0809_ _0959_ _0961_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2633_ _0107_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_2495_ _1104_ _0682_ _0688_ _0686_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1446_ _0882_ _0890_ _0894_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1377_ _0774_ _0778_ _0816_ _0814_ _0825_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_4_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1763__B _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2655__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2280_ _0524_ _0525_ _0527_ _0529_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1300_ _0722_ _0728_ _0743_ _0748_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_47_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1995_ _0296_ _0298_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2616_ _0090_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2547_ _0021_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1429_ _0715_ _0877_ _0726_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2478_ _0715_ _0673_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2488__C _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2528__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2678__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1780_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\] _0913_ _1193_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1650__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2332_ _0574_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2401_ _1108_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2263_ _0456_ _0517_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2194_ _0833_ _0457_ _0461_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ _0275_ net1 _0279_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2360__A2 _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1871__A1 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1832_ _1232_ _1234_ _1235_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1901_ tt_um_rejunity_sn76489.clk_counter\[5\] tt_um_rejunity_sn76489.clk_counter\[4\]
+ _0219_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_8_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1763_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\] _1179_ _1157_ _1180_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1694_ _1096_ _1121_ _1124_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2315_ _0558_ _0561_ _0539_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2246_ _0281_ _0500_ _0503_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2177_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\] _0441_ _0448_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_50_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2073__I _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput14 net14 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput25 net25 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2716__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2100_ _0361_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2031_ _0323_ _0924_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1815_ _1218_ _1222_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1746_ _1142_ _1166_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1677_ net3 _1112_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2229_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\] _0355_ _0489_ _0490_ _0482_
+ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__2012__A1 _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1600_ _1024_ _1037_ _1021_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1531_ _0926_ _0944_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1462_ _0909_ _0910_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_10_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2580_ _0054_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1393_ tt_um_rejunity_sn76489.chan\[0\].attenuation.in _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2014_ _0307_ _0801_ _0310_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2561__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1729_ _1149_ _1151_ _1152_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2481__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2701_ _0175_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2584__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2632_ _0106_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1445_ _0830_ _0848_ _0893_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2563_ _0037_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1514_ _0960_ net45 _0888_ _0809_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_10_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ _0777_ _0683_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1376_ _0773_ _0767_ _0775_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_4_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1994_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\] _0293_ _0297_ _0298_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2166__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2445__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ _0089_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2546_ _0020_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1428_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\] tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
+ _0717_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2477_ _1095_ _0672_ _0675_ _0676_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_38_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1359_ _0805_ _0806_ _0760_ _0807_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_21_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _1105_ _0611_ _0619_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2331_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\] _0573_ _0574_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2262_ tt_um_rejunity_sn76489.pwm.accumulator\[1\] _0513_ _0516_ _0517_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_35_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2418__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2193_ _0833_ _0457_ _0460_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1977_ _1140_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2529_ _0003_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1703__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1831_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\] _0811_ _1235_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1900_ _0223_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1762_ _0779_ _0784_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1693_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\] _1122_ _1115_ _1124_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2314_ _0559_ _0560_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_27_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2176_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2245_ _0287_ _0500_ _0503_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_11_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2303__B _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput15 net15 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput26 net26 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ _0322_ _0324_ _0325_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1814_ _1219_ _1055_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1745_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\] _1014_ _1165_ _1166_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1676_ _1110_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2159_ _0428_ _0432_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2228_ _0485_ _0488_ _0475_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2260__A2 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ _0944_ _0926_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1461_ _0778_ _0834_ _0779_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1392_ _0751_ _0762_ _0752_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_22_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1801__I _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ _0309_ _0311_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1728_ _1149_ _1151_ _1127_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2706__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1659_ _1097_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_48_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2562_ _0036_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2700_ _0174_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2631_ _0105_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1444_ _0891_ _0892_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1375_ _0802_ _0819_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1513_ _0750_ _0842_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2493_ _1101_ _0682_ _0687_ _0686_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_2_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2551__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1993_ _1098_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2545_ _0019_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1708__A1 _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2614_ _0088_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1427_ _0732_ _0873_ _0874_ _0742_ _0875_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1358_ _0758_ _0762_ _0752_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2476_ _1092_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_41_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1289_ tt_um_rejunity_sn76489.chan\[3\].attenuation.in _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2330_ _1078_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2261_ _0802_ _0819_ _0515_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2192_ _0209_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ _0220_ _0282_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2528_ _0002_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2459_ _0654_ _0661_ _0663_ _1093_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2036__B _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1785__B _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1761_ _1177_ _1175_ _1178_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1830_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\] _0811_ _1234_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2313_ _0553_ _0554_ _0556_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1692_ _1118_ _1121_ _1123_ _1093_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1311__A2 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2175_ _0446_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2244_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\] _0492_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
+ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_7_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1959_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\] _0260_ _0269_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput16 net16 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput27 net27 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_3_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2612__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1813_ _1218_ _1220_ _1221_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1744_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\] _0984_ _1164_ _1165_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1675_ _1110_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2158_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\] _0426_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
+ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2635__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2227_ _0485_ _0488_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2089_ _0370_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2658__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1460_ _0844_ net46 _0761_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1391_ _0758_ _0763_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_54_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2012_ _0224_ _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1727_ _1150_ _0923_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1692__C _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1658_ net12 _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1589_ _1030_ _0967_ _1033_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_5_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1680__A1 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2561_ _0035_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1512_ _0806_ _0807_ _0843_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2630_ _0104_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2492_ _0815_ _0683_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1443_ net58 _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1374_ _0822_ _0796_ _0799_ _0800_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1662__A1 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1992_ _0295_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2544_ _0018_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2613_ _0087_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2475_ _0716_ _0673_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1357_ _0750_ _0754_ _0752_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_1426_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _0737_ _0730_ _0875_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1288_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _0737_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__1717__I _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2124__A2 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2260_ net41 _0786_ _0514_ _0749_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2191_ _0456_ _0459_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1975_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\] _0281_ _0282_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2354__A2 _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1409_ _0716_ _0723_ _0718_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2458_ _0795_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2527_ _0001_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1272__I _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2389_ _0610_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2042__A1 _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2541__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2691__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1760_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\] _1064_ _1157_ _1178_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_40_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1691_ net3 _1122_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2312_ tt_um_rejunity_sn76489.pwm.accumulator\[8\] net23 _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2174_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\] _0425_ _0443_ _0445_ _0439_
+ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2243_ _0498_ _0353_ _0501_ _0502_ _1141_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput17 net17 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 net28 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_rebuffer10_I _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1378__A3 _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2564__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1889_ _0212_ tt_um_rejunity_sn76489.clk_counter\[1\] tt_um_rejunity_sn76489.clk_counter\[2\]
+ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1958_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\] _0263_ _0268_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2047__B _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2263__A1 _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2510__B _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1829__A1 _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2587__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2254__A1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1812_ _1218_ _1220_ _1203_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1743_ _1161_ _1163_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1674_ _1086_ _1109_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2226_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\] _0478_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
+ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2157_ _0431_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2493__A1 _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2088_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\] _0373_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
+ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2245__A1 _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2381__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2484__A1 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1390_ _0832_ _0835_ _0837_ _0838_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_54_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ _0305_ _0308_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2475__A1 _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1588_ _1031_ _1032_ _0968_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1726_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[4\] _1150_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1657_ _1095_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2209_ _0470_ _0473_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2466__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2560_ _0034_ clknet_4_5_0_wb_clk_i net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1511_ _0951_ _0957_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1442_ _0839_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2625__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2491_ _1095_ _0682_ _0685_ _0686_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_49_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1373_ _0794_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2448__A1 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1709_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\] _0822_ _1135_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2689_ _0163_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1991_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\] _0293_ _0295_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2612_ _0086_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2543_ _0017_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1425_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _0731_ _0874_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2474_ _0654_ _0672_ _0674_ _0665_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1356_ _0803_ _0804_ _0763_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1287_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _0736_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_21_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1580__A1 _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1643__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2190_ _0453_ _0458_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1974_ _0280_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2526_ _0000_ clknet_4_13_0_wb_clk_i net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1408_ _0712_ _0724_ _0713_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2457_ _0660_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2388_ _0610_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1339_ _0722_ _0728_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1690_ _1120_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2311_ tt_um_rejunity_sn76489.pwm.accumulator\[9\] net24 _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1544__A1 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2242_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] _0499_ _0495_ _0502_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2173_ _0289_ _0444_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1957_ _0266_ _0267_ _0262_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2709__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput18 net18 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1888_ _1140_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2509_ _1085_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1811_ _1219_ _1055_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1742_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\] _0984_ _1163_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1673_ _1081_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1317__B _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2225_ _0487_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1296__A3 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2531__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2156_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\] _0425_ _0428_ _0430_ _0419_
+ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2087_ _0358_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2681__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2236__A2 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ _0305_ _0308_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1651__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2554__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1725_ _1145_ _1147_ _1148_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1587_ _0910_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1656_ _1094_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2139_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\] _0413_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
+ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2208_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\] _0465_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
+ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2392__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1441_ _0885_ _0889_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1510_ _0727_ _0955_ _0956_ _0861_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_4_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2490_ _0223_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1372_ _0749_ _0791_ _0820_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1330__B _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1708_ _1132_ _1134_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2688_ _0162_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1639_ _1079_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_18_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1990_ _0293_ _0294_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2611_ _0085_ clknet_4_7_0_wb_clk_i net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2542_ _0016_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1424_ _0850_ _0741_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1355_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _0804_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2473_ _0723_ _0673_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1286_ _0732_ _0733_ _0734_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_21_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2615__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2348__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2520__A1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _0275_ net1 _0278_ _0279_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__2490__I _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1834__I _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2525_ _0706_ _0703_ _0707_ _0695_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1338_ net41 _0786_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1407_ _0715_ _0718_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2638__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2511__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ _0606_ _0607_ _0608_ _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2456_ _0660_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1269_ _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2508__C _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2502__A1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2243__C _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2310_ _0541_ _0557_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2172_ _0437_ _0442_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2241_ _0396_ _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2485__I _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1887_ _0194_ _0214_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1956_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\] _0260_ _0267_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput19 net54 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2508_ _1104_ _0691_ _0697_ _0695_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2439_ _0642_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_54_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2519__B _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1810_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[8\] _1219_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1741_ _1142_ _1162_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1672_ net7 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2155_ _0422_ _0427_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2224_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\] _0468_ _0485_ _0486_ _0482_
+ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_0_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2086_ _0372_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1939_ _0253_ _0254_ _0251_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2181__A2 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1435__A1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1683__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1724_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\] _0901_ _1148_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1586_ _0909_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1655_ net4 _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2207_ _0472_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2138_ _0410_ _0415_ _0213_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2069_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
+ _0356_ _0357_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1752__I _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1701__B _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1371_ _0819_ _0802_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1440_ _0803_ _0886_ _0887_ _0888_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_4_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2671__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1638_ _1076_ _1078_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1707_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\] _0822_ _1133_ _1134_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2687_ _0161_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1569_ _1004_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2544__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2694__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2610_ _0084_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2541_ _0015_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2472_ _0671_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1657__I _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1877__A1 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1423_ _0868_ _0863_ _0871_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1285_ _0729_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1354_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\] _0803_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_46_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2567__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ tt_um_rejunity_sn76489.clk_counter\[0\] tt_um_rejunity_sn76489.clk_counter\[1\]
+ tt_um_rejunity_sn76489.clk_counter\[3\] tt_um_rejunity_sn76489.clk_counter\[2\]
+ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_7_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2455_ _0655_ _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2524_ net5 _0703_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1337_ _0761_ _0766_ net48 _0784_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1406_ _0849_ _0850_ _0851_ _0852_ _0854_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1268_ _0708_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2386_ tt_um_rejunity_sn76489.latch_control_reg\[2\] _1084_ _0609_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_46_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2171_ _0437_ _0442_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2240_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] _0495_ _0499_ _0500_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_43_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1886_ _0212_ tt_um_rejunity_sn76489.clk_counter\[1\] _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1955_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\] _0263_ _0266_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2605__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2438_ _0632_ _0643_ _0647_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2507_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _0692_ _0697_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2369_ _0598_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1740_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\] _0984_ _1161_ _1162_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_40_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2628__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1671_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\] _1107_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input8_I io_in_1[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2223_ _0480_ _0484_ _0475_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2154_ _0288_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2085_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\] _0362_ _0370_ _0371_ _0297_
+ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_16_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1869_ _0197_ _0199_ _0200_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1938_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\] _0249_ _0254_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2090__B _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1723_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\] _0901_ _1147_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1654_ _1080_ _1088_ _1090_ _1093_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1585_ _1028_ _1029_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1371__A1 _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2206_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\] _0468_ _0470_ _0471_ _0439_
+ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_0_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2137_ _0355_ _0414_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2068_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
+ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
+ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_48_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1370_ _0811_ _0818_ _0785_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1637_ net12 _1077_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1706_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\] _0788_ _1133_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2686_ _0160_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1568_ _1011_ _1012_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1499_ _0946_ net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__1344__A1 _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1422_ _0869_ _0870_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2540_ _0014_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2471_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1353_ _0794_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1284_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _0733_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_46_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2669_ _0143_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1971_ _0276_ _0277_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1668__I _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1405_ _0849_ _0850_ _0853_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2523_ tt_um_rejunity_sn76489.control_noise\[0\]\[2\] _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2385_ net11 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_11_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2454_ _0656_ _0657_ _0658_ _0609_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xinput1 custom_settings[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1336_ _0761_ _0766_ _0779_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_1267_ _0711_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2534__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2202__I _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2684__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2557__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2170_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\] _0441_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
+ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1954_ _0264_ _0265_ _0262_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1885_ _0212_ _0213_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2368_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\] _0596_ _0593_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\]
+ _0597_ net21 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1861__I _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2437_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\] _0644_ _0646_ _0647_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2506_ _1101_ _0691_ _0696_ _0695_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_54_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2299_ tt_um_rejunity_sn76489.pwm.accumulator\[6\] _0980_ _0543_ _0544_ _0548_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1319_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_34_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2184__A1 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ _1105_ _1088_ _1106_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2222_ _0480_ _0484_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1681__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2153_ _0422_ _0427_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2084_ _0364_ _0369_ _0366_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1937_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\] _0252_ _0253_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1868_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\] _0994_ _0200_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1799_ _1207_ _1208_ _1209_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1722_ _1142_ _1146_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1584_ _0939_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ _1092_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2205_ _0466_ _0469_ _0429_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2136_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\] _0413_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
+ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2067_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
+ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
+ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_36_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2210__I _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2618__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2085__C _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1705_ _1131_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1567_ _0976_ _0979_ _0987_ _1009_ _0981_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1636_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\] tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
+ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2685_ _0159_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1498_ _0922_ _0945_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_1_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2186__B _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2119_ _0395_ _0353_ _0399_ _0400_ _0283_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1271__A1 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1421_ _0862_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2470_ _0655_ _0670_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_50_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1352_ _0796_ _0799_ _0800_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1283_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _0732_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_46_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2668_ _0142_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1619_ _1062_ net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2599_ _0073_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2505__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ _0275_ net1 _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2522_ _0632_ _0703_ _0705_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1335_ _0782_ _0776_ _0783_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1404_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _0795_ _0734_ _0853_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2453_ _0606_ tt_um_rejunity_sn76489.latch_control_reg\[0\] _0658_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2384_ tt_um_rejunity_sn76489.latch_control_reg\[0\] _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput2 custom_settings[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1266_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\] _0715_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1884_ _1131_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1953_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\] _0260_ _0265_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2193__A2 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2505_ _0803_ _0692_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2298_ tt_um_rejunity_sn76489.pwm.accumulator\[6\] net21 _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2367_ _0581_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1318_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _0767_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2436_ _0614_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_54_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2651__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2674__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2221_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\] _0478_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
+ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2152_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\] _0426_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
+ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1438__A1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2083_ _0364_ _0369_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1867_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\] _0994_ _0199_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1936_ _0231_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1798_ _1207_ _1208_ _1203_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1677__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2419_ _1101_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2547__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1721_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\] _0901_ _1145_ _1146_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1583_ _0935_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1652_ _1091_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2204_ _0466_ _0469_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2135_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
+ _0411_ _0412_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2066_ _0288_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1919_ _0235_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_27_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2712__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _1130_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2684_ _0158_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1566_ _0987_ _1009_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1497_ _0926_ _0944_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1635_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\] _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2049_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\] _1015_ _0341_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2118_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] _0397_ _0392_ _0400_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1271__A2 _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1420_ _0855_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1351_ _0733_ _0746_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1282_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\] _0730_ _0731_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1618_ _1043_ _1061_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2608__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2667_ _0141_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1549_ _0993_ _0994_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2598_ _0072_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1880__I _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_39_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2441__A1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2521_ tt_um_rejunity_sn76489.control_noise\[0\]\[1\] _0702_ _1092_ _0705_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1265_ _0710_ _0712_ _0713_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1403_ _0736_ _0733_ _0739_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1334_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\] _0768_ _0783_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2452_ net9 net10 _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2383_ tt_um_rejunity_sn76489.latch_control_reg\[1\] _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 io_in_1[0] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output15_I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2390__B _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1883_ tt_um_rejunity_sn76489.clk_counter\[0\] _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1952_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\] _0263_ _0264_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2504_ _1095_ _0691_ _0694_ _0695_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_3_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2435_ _0605_ _0643_ _0645_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2366_ _1079_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2297_ _0541_ _0546_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1317_ _0753_ _0764_ _0765_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_2_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2459__C _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2404__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ _0483_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2151_ _0413_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2082_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\] _0358_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
+ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1866_ _0194_ _0198_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1797_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\] _0998_ _1208_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_26_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1935_ _0248_ _0250_ _0251_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2418_ _0632_ _0629_ _0633_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_10_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2349_ _0581_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1720_ _1143_ _1144_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1651_ net12 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1582_ _0963_ _0832_ _0836_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1356__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2641__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I io_in_1[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2203_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\] _0465_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
+ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2134_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
+ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
+ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2065_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\] _0353_ _0354_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1831__A2 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1849_ _1247_ _1031_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1918_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\] _0238_ _0239_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1968__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1634_ _1075_ net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_41_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1703_ net12 _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2683_ _0157_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1565_ _1010_ net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1496_ _0931_ _0943_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2048_ _0338_ _0339_ _0340_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_1_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2537__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2117_ _0396_ _0398_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2687__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1559__A1 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1350_ _0797_ _0742_ _0798_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1281_ _0729_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_46_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1698__I _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1617_ _1044_ _1060_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2666_ _0140_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2597_ _0071_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1548_ _0991_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1479_ _0857_ _0904_ _0727_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_49_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2702__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1402_ _0742_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1981__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2142__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2451_ _1081_ _1082_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2520_ _0605_ _0703_ _0704_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1264_ tt_um_rejunity_sn76489.chan\[2\].attenuation.in _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1333_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _0780_ _0781_ _0782_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xinput4 io_in_1[1] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2382_ _0604_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2718_ _0192_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.control_noise\[0\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2649_ _0123_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_40_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1882_ _0208_ _0206_ _0211_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1951_ _0230_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_47_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2365_ _0595_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2434_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\] _0644_ _0638_ _0645_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2503_ _0223_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_54_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2296_ tt_um_rejunity_sn76489.pwm.accumulator\[6\] net21 _0545_ _0546_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1316_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _0755_ _0765_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_2_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2150_ _0361_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2081_ _0368_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2570__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1934_ _0234_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1865_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\] _0994_ _0197_ _0198_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1796_ _1205_ _1206_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2348_ _0283_ _0582_ _0584_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_3_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2417_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\] _0630_ _0624_ _0633_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2279_ tt_um_rejunity_sn76489.pwm.accumulator\[4\] _0898_ net53 _0531_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1581_ _1025_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1650_ net3 _1089_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1356__A2 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2202_ _0361_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2150__I _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2133_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
+ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
+ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2064_ _0280_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1292__A1 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1917_ _0237_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1779_ _1171_ _1192_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1848_ _1246_ _1248_ _1249_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1338__A2 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ _1067_ _1069_ _1074_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1564_ _0982_ _0987_ _1009_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1702_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\] _0788_ _1129_ _0013_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2682_ _0156_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1495_ _0941_ _0942_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2047_ _0338_ _0339_ _0330_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2116_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] _0392_ _0397_ _0398_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_12_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2508__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1280_ tt_um_rejunity_sn76489.chan\[3\].attenuation.in _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1616_ _1047_ _1059_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1547_ _0989_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2665_ _0139_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1970__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2596_ _0070_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2654__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1478_ _0923_ _0924_ _0925_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_37_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2423__I _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2450_ _0608_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1401_ _0737_ _0744_ _0738_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__2527__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2381_ net3 _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1263_ _0711_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1332_ _0768_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xinput5 io_in_1[2] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2717_ _0191_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.control_noise\[0\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2648_ _0122_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2579_ _0053_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1950_ _0259_ _0261_ _0262_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1881_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\] _1052_ _0210_ _0211_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2502_ _0804_ _0692_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2364_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\] _0589_ _0593_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\]
+ _0585_ net20 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2350__A2 _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1315_ _0758_ _0762_ _0763_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2433_ _0642_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_54_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2295_ _0543_ _0544_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2080_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\] _0362_ _0364_ _0367_ _0297_
+ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1933_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\] _0249_ _0250_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1864_ _0195_ _0196_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1795_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\] _1029_ _1201_ _1206_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_12_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2278_ _0529_ _0527_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2347_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\] _0575_ _0583_ _0584_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2416_ _1094_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1580_ _0843_ _0886_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2201_ _0462_ _0467_ _1132_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2132_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\] _0403_ _0410_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2063_ _0352_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1847_ _1246_ _1248_ _1238_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1916_ tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
+ _0229_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2241__A1 _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1778_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\] _0913_ _1191_ _1192_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_8_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2663__D _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2480__A1 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2560__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1701_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\] _0788_ _1127_ _1129_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2681_ _0155_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1632_ _1070_ _1072_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1563_ _1002_ _1008_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1494_ _0932_ _0933_ _0940_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_30_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2115_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\] _0389_ _0397_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2046_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\] _1015_ _0339_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2462__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2583__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_sn76489_40 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2664_ _0138_ clknet_4_14_0_wb_clk_i net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1615_ _1054_ _1058_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1546_ _0989_ _0991_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1477_ _0908_ _0917_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2595_ _0069_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_37_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2029_ _0322_ _0324_ _0210_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2435__A1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2426__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1400_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _0730_ _0849_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2380_ _0215_ _0229_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1331_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _0780_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_36_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1262_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\] _0711_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput6 io_in_1[3] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2647_ _0121_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2716_ _0190_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1529_ _0971_ _0975_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2578_ _0052_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2408__A1 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ _0209_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2501_ _0654_ _0691_ _0693_ _0686_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_3_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2363_ _0594_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2294_ _0542_ _0946_ _0536_ _0534_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1314_ _0755_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_2432_ _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_54_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2667__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1863_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\] _0997_ _1257_ _0196_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1932_ _0237_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1794_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\] _1029_ _1205_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2415_ _0605_ _0629_ _0631_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2346_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\] tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
+ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2277_ tt_um_rejunity_sn76489.pwm.accumulator\[3\] _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2074__I _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2062_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\] _1063_ _0351_ _1228_
+ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2131_ _0952_ _0406_ _0409_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2200_ _0289_ _0466_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1777_ _1185_ _1186_ _1190_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1846_ _1247_ _1031_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1915_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\] _0232_ _0236_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2329_ _0571_ net42 _0572_ _0215_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input12_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2705__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1631_ _1073_ net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2680_ _0154_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1700_ _1105_ _1121_ _1128_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1562_ _1007_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1493_ _0932_ _0933_ _0940_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2045_ _0334_ _0336_ _0337_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input4_I io_in_1[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2114_ _0280_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1829_ _1211_ _1233_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_sn76489_30 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2663_ _0137_ clknet_4_13_0_wb_clk_i net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1614_ _1025_ _1055_ _1057_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2594_ _0068_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1476_ _0907_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1545_ _0764_ _0844_ _0846_ _0990_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_22_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2380__A1 _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2028_ _0323_ _0924_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_37_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2550__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2123__A1 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1330_ _0770_ _0772_ _0776_ _0778_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_1261_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\] _0710_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 io_in_1[4] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2646_ _0120_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2577_ _0051_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2715_ _0189_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1528_ _0931_ _0943_ _0974_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1459_ _0905_ _0907_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2077__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2500_ _0754_ _0692_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2431_ _0606_ _0607_ _0608_ _0627_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_47_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2293_ _0542_ _0946_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2362_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\] _0589_ _0593_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\]
+ _0585_ net54 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_1313_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\] _0762_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_44_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1377__A2 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2326__A1 _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2629_ _0103_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2611__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1862_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\] _0997_ _0195_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput10 io_in_1[7] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1793_ _1201_ _1202_ _1204_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1931_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\] _0241_ _0248_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2414_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\] _0630_ _0624_ _0631_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2345_ _1076_ _1077_ net16 _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2276_ _0456_ _0528_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2634__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2061_ _0346_ _0350_ _0347_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1513__A2 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2130_ _0952_ _0406_ _0330_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1277__A1 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1914_ _0734_ _0232_ _0233_ _0235_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1776_ _1187_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1845_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[4\] _1247_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2328_ tt_um_rejunity_sn76489.pwm.accumulator\[11\] net26 _0572_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2657__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2259_ _0722_ _0728_ _0743_ _0748_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1440__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1630_ net55 _1070_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1431__A1 _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1561_ _1004_ _1006_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1492_ _0935_ _0939_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_49_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2044_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\] _0983_ _0337_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2113_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1670__A1 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1759_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\] _1064_ _1177_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1828_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\] _0811_ _1232_ _1233_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1973__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2029__B _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_sn76489_31 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1613_ _1034_ _1035_ _0995_ _1056_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2662_ _0136_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1544_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] net51 _0990_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2593_ _0067_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1475_ _0905_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2132__A2 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[4\] _0323_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_37_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1891__A1 _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1398__B1 _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 io_in_1[5] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1260_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\] _0708_ _0709_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_34_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2714_ _0188_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.latch_control_reg\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2353__A2 _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1527_ _0972_ _0973_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2645_ _0119_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2576_ _0050_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1389_ _0812_ _0780_ _0775_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1458_ _0906_ _0851_ _0743_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1881__B _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1900__I _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2361_ _0574_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2430_ _0623_ _0630_ _0641_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2292_ tt_um_rejunity_sn76489.pwm.accumulator\[5\] _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1312_ _0753_ _0757_ _0759_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__2690__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2023__A1 _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2559_ _0033_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2628_ _0102_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2563__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ _0246_ _0247_ _0240_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2253__A1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput11 io_in_2 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1792_ _1201_ _1202_ _1203_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1861_ _1210_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2344_ _0581_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2413_ _0628_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2275_ tt_um_rejunity_sn76489.pwm.accumulator\[3\] _0526_ _0527_ _0528_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2586__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__A1 _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2060_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\] _1063_ _0350_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_53_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1360__I _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2474__A1 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1913_ _0234_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1775_ _1171_ _1189_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1844_ _1242_ _1244_ _1245_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_8_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2327_ tt_um_rejunity_sn76489.pwm.accumulator\[11\] net26 _0571_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2258_ tt_um_rejunity_sn76489.pwm.accumulator\[0\] _0511_ _0513_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2465__A1 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2189_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\] _0457_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
+ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2315__B _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_18_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ _0854_ _0851_ _0745_ _1005_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_1491_ _0825_ _0936_ _0938_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2112_ _0394_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2043_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\] _0983_ _0336_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2119__C _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\] _1230_ _1232_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1758_ _1171_ _1176_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2624__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1689_ _1120_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2438__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_sn76489_32 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2661_ _0135_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1612_ _1025_ _1027_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1474_ _0898_ _0919_ _0921_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1543_ _0936_ _0988_ _0963_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2592_ _0066_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_37_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2026_ _0318_ _0320_ _0321_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_9_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 io_in_1[6] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2644_ _0118_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_2713_ _0187_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.latch_control_reg\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1526_ _0930_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1457_ _0853_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2575_ _0049_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1388_ _0813_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1699__B _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2009_ _0307_ _0801_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _0527_ _0137_ _0592_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1311_ _0756_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _0760_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
X_2291_ _1131_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2627_ _0101_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2558_ _0032_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1509_ _0953_ _0904_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2489_ _0812_ _0683_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2053__B _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2708__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1828__A2 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1860_ _1257_ _1258_ _0193_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1791_ _1126_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput12 rst_n net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2274_ _0867_ _0896_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_2343_ _1130_ _1077_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2412_ _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2138__B _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1821__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1268__I _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1989_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\] _0292_ _1228_ _0294_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer20_I _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1286__A3 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2530__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2680__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1641__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\] _0914_ _1245_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1912_ _1130_ tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise _0234_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1774_ _1185_ _1188_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2326_ _0541_ _0570_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1551__I _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2257_ tt_um_rejunity_sn76489.pwm.accumulator\[0\] _0511_ _0512_ _0119_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_4_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2553__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2188_ _0286_ _0441_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1490_ _0832_ _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2042_ _0315_ _0335_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2111_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\] _0384_ _0391_ _0393_ _0377_
+ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_49_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1826_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\] _1230_ _1231_ _0035_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1757_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\] _1064_ _1175_ _1176_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_40_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1688_ _1081_ _1082_ _1119_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2309_ _0555_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input10_I io_in_1[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2126__A1 _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_sn76489_33 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_46_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1611_ _1027_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2660_ _0134_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1404__A3 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1473_ _0903_ _0918_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1542_ _0832_ _0835_ _0782_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2591_ _0065_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2117__A1 _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I custom_settings[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2025_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\] _0900_ _0321_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1809_ _1214_ _1216_ _1217_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2614__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2574_ _0048_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2712_ _0186_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.latch_control_reg\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2643_ _0117_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1525_ _0928_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1456_ _0904_ _0721_ _0722_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1387_ _0773_ _0812_ _0775_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_22_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2008_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[1\] _0307_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1734__I _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2637__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2501__A1 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2290_ _0537_ _0538_ _0540_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1310_ _0758_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _0756_ _0759_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__1644__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2557_ _0031_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2626_ _0100_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1508_ _0953_ _0904_ _0954_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1439_ _0803_ _0751_ _0763_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2488_ _0654_ _0682_ _0684_ _0676_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2385__I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1790_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\] _1029_ _1202_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1461__A1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2411_ _0626_ _0607_ _0608_ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2342_ _0573_ _0580_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2273_ _0524_ _0525_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1988_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\] _0292_ _0293_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2609_ _0083_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1691__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1773_ _1186_ _1187_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1842_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\] _0914_ _1244_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\] _0231_ _0233_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_12_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2325_ tt_um_rejunity_sn76489.pwm.accumulator\[11\] net26 _0569_ _0570_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_40_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2256_ tt_um_rejunity_sn76489.pwm.accumulator\[0\] _0511_ _0460_ _0512_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2187_ _1131_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2506__C _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2041_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\] _0983_ _0334_ _0335_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2110_ _0289_ _0392_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1756_ _1169_ _1173_ _1174_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1825_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\] _1230_ _1203_ _1231_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2308_ tt_um_rejunity_sn76489.pwm.accumulator\[8\] _1013_ _1039_ _0556_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1894__A1 _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1687_ net9 _1085_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2670__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2239_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\] _0492_ _0499_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_23_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2071__A1 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_sn76489_34 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_41_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1637__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1610_ _1050_ _1053_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2590_ _0064_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1541_ _0985_ _0986_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1472_ _0920_ net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2543__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2024_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\] _0900_ _0320_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2693__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1808_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\] _0993_ _1217_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1739_ _1159_ _1160_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2566__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2072__B _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2283__A1 _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2711_ _0185_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1524_ _0958_ _0970_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2573_ _0047_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2642_ _0116_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1455_ _0858_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1386_ _0773_ _0833_ _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_10_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2007_ _0305_ _0306_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2514__C _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1660__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2556_ _0030_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1507_ _0953_ _0709_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2625_ _0099_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2487_ _0767_ _0683_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1438_ _0804_ _0757_ _0765_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1369_ _0812_ _0813_ _0817_ net59 _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__2495__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2334__C _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2341_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\] _0578_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
+ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2410_ tt_um_rejunity_sn76489.latch_control_reg\[2\] net10 _0627_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_2
X_2272_ tt_um_rejunity_sn76489.pwm.accumulator\[2\] _0521_ _0520_ _0525_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2486__I _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2477__A1 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2627__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1987_ _0283_ _0290_ _0292_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_15_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2608_ _0082_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2539_ _0013_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2329__C _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2345__B net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2459__A1 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1910_ _0231_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1772_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\] _0891_ _1187_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1841_ _1211_ _1243_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1370__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2324_ _0565_ _0567_ _0568_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2255_ _0787_ _0790_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_25_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2186_ _0453_ _0455_ _1132_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _0328_ _0332_ _0333_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_17_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1755_ _1172_ _1022_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1824_ _0761_ _0766_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1686_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\] _1118_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2307_ _0553_ _0554_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2238_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2169_ _0426_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_31_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1885__A2 _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_sn76489_35 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1540_ _0958_ _0970_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1471_ net57 net53 _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1663__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2023_ _0315_ _0319_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1807_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\] _0993_ _1216_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1738_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\] _0972_ _1155_ _1160_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1669_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\] _1089_ _1099_ _1106_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1316__A1 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2710_ _0184_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__1658__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1523_ _0969_ _0967_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1454_ _0882_ _0899_ _0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2572_ _0046_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2641_ _0115_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1385_ _0771_ _0767_ _0769_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2006_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\] _0789_ _0297_ _0306_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2533__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1700__A1 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2624_ _0098_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2555_ _0029_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1437_ _0760_ _0841_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1506_ _0710_ _0952_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2486_ _0681_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2556__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1299_ _0745_ _0740_ _0747_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1368_ _0814_ _0816_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2247__A2 _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2183__A1 _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2525__C _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2410__A2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2340_ _0573_ _0579_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2271_ tt_um_rejunity_sn76489.pwm.accumulator\[2\] _0521_ _0524_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2229__A2 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1986_ _0291_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2607_ _0081_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2469_ _0657_ _0668_ _0669_ _0609_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2538_ _0012_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2080__C _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\] _0914_ _1242_ _1243_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_29_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1771_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\] _0891_ _1186_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2395__A1 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2323_ tt_um_rejunity_sn76489.pwm.accumulator\[10\] _1073_ _0568_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2254_ _0842_ _0507_ _0510_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2185_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\] _0403_ _0454_ _0455_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ tt_um_rejunity_sn76489.clk_counter\[5\] tt_um_rejunity_sn76489.clk_counter\[4\]
+ tt_um_rejunity_sn76489.clk_counter\[6\] _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2310__A1 _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2129__A1 _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2617__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1823_ _1226_ _1229_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1754_ _1172_ _1022_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1685_ _1105_ _1111_ _1117_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2306_ _0550_ _1010_ _0547_ _0548_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2237_ _0497_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2099_ _0383_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2168_ _0440_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xwrapped_sn76489_36 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1470_ _0918_ _0903_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_22_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2522__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2022_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\] _0900_ _0318_ _0319_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_9_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1806_ _1211_ _1215_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_20_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1599_ _1011_ net43 _1041_ _1042_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_1737_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\] _0972_ _1159_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2513__A1 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1668_ _1104_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1713__B _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2504__A1 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _0114_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2571_ _0045_ clknet_4_5_0_wb_clk_i net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1522_ _0968_ _0941_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1453_ _0900_ _0901_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2005_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\] _0789_ _0305_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1384_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2554_ _0028_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2623_ _0097_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1436_ _0836_ _0883_ _0884_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_1367_ _0777_ _0815_ _0781_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1505_ _0713_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2485_ _0681_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1298_ _0746_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1694__A1 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2650__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1438__B _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2269__B _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2270_ _0520_ _0522_ _0523_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1685__A1 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1985_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\] tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
+ _0285_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2606_ _0080_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2537_ _0011_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2673__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1419_ _0830_ net49 _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2468_ _0626_ tt_um_rejunity_sn76489.latch_control_reg\[0\] _0669_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2399_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\] _0617_ _0615_ _0619_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1770_ _1181_ _1183_ _1184_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2546__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2322_ tt_um_rejunity_sn76489.pwm.accumulator\[10\] net25 _0567_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_2
X_2253_ _0842_ _0507_ _0460_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2184_ _0281_ _0449_ _0452_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_47_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__I _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1968_ net2 _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_28_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1899_ _1091_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__C _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2569__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1822_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\] _1051_ _1228_ _1229_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1753_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\] _1172_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1684_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\] _1112_ _1115_ _1117_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2305_ _0550_ _1010_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2167_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\] _0425_ _0437_ _0438_ _0439_
+ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_0_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2236_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\] _0355_ _0494_ _0496_ _0482_
+ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_48_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2098_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\] _0362_ _0380_ _0382_ _0377_
+ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__2711__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2359__A2 _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_sn76489_37 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1270__A2 _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2021_ _0312_ _0316_ _0317_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_15_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1805_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\] _0993_ _1214_ _1215_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1736_ _1155_ _1156_ _1158_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1356__B _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1598_ _1017_ _1038_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1667_ net6 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2219_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\] _0468_ _0480_ _0481_ _0482_
+ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_51_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_46_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2607__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2570_ _0044_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1521_ _0935_ _0939_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1452_ _0881_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1383_ _0831_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _0220_ _0304_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1719_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\] _0870_ _1137_ _1144_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2699_ _0173_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2422__A1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2553_ _0027_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1504_ _0747_ _0949_ _0950_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2622_ _0096_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1435_ _0778_ _0838_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1366_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _0815_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2484_ _0655_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1297_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _0730_ _0746_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1437__A2 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1984_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\] _0289_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
+ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2605_ _0079_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2536_ _0010_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2467_ _0622_ _1082_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1418_ _0821_ _0865_ _0866_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1349_ _0737_ _0795_ _0738_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2398_ _1102_ _0611_ _0618_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_6_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2321_ _0541_ _0566_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2183_ _0365_ _0449_ _0452_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2252_ _0456_ _0509_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1830__A2 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1898_ tt_um_rejunity_sn76489.clk_counter\[4\] _0219_ tt_um_rejunity_sn76489.clk_counter\[5\]
+ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _0232_ _0273_ _0274_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1822__B _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2640__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2519_ tt_um_rejunity_sn76489.control_noise\[0\]\[0\] _0702_ _0652_ _0704_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_3_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2065__A2 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2663__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1752_ _1141_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_29_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ _1102_ _1111_ _1116_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1821_ _1227_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2304_ _0549_ _0551_ _0552_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2166_ _1227_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2097_ _0375_ _0379_ _0381_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2235_ _0366_ _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2056__A2 _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_sn76489_38 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_39_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2536__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2686__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\] _0869_ _0317_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1804_ _1212_ _1213_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1735_ _1155_ _1156_ _1157_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1666_ _1102_ _1088_ _1103_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1597_ _1017_ _1038_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2559__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2149_ _0424_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2218_ _1098_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1520_ _0962_ _0966_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1451_ _0876_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1382_ _0771_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _0769_ _0831_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2701__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2003_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\] _0302_ _0304_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1718_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\] _0870_ _1143_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2698_ _0172_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1649_ _1087_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_16_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1791__I _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2110__A1 _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2552_ _0026_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1503_ _0947_ _0906_ _0747_ _0875_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2483_ _0627_ _0658_ _0679_ _0656_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2621_ _0095_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1434_ _0815_ _0783_ _0831_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1296_ _0732_ _0744_ _0734_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1365_ _0771_ _0780_ _0781_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_5_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1391__A2 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1735__B _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2604_ _0078_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1983_ _0288_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2398__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1417_ _0824_ _0864_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2466_ _0637_ _0661_ _0667_ _0665_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2535_ _0009_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_43_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1279_ _0725_ _0714_ _0727_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1348_ _0736_ _0738_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2397_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\] _0617_ _0615_ _0618_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_6_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2320_ tt_um_rejunity_sn76489.pwm.accumulator\[10\] net25 _0565_ _0566_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2251_ _0504_ _0508_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2182_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\] _0441_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
+ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1966_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\] _0232_ _0235_ _0274_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_50_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1897_ _0220_ _0221_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2518_ _0702_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2449_ _0604_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1820_ _1091_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ _1142_ _1170_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1682_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\] _1112_ _1115_ _1116_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1974__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2303_ _0549_ _0551_ _0539_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2234_ _0489_ _0493_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2165_ _0433_ _0436_ _0429_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2096_ _0288_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_0_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1949_ _0234_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2516__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_sn76489_39 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_34_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2507__A1 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1803_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\] _0998_ _1207_ _1213_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2630__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1596_ _1040_ net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1734_ _1126_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1665_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\] _1089_ _1099_ _1103_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2217_ _0474_ _0479_ _0475_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2148_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\] _0384_ _0422_ _0423_ _0419_
+ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2079_ _0359_ _0363_ _0366_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1879__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2503__I _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2653__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1450_ _0890_ _0894_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1381_ _0829_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_33_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2002_ _0301_ _0303_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2195__A2 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1579_ _1021_ _1023_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2526__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1717_ _1141_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2697_ _0171_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1648_ _1087_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2676__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2549__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2620_ _0094_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2551_ _0025_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1433_ _0876_ _0881_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1502_ _0947_ _0906_ _0948_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1982__I _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2482_ _1083_ net10 _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1364_ _0783_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1295_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\] _0744_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__2481__C _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _0287_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2603_ _0077_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2534_ _0008_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1416_ _0824_ _0864_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1347_ _0736_ _0795_ _0739_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2396_ _0610_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2465_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _0662_ _0667_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1278_ _0726_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2714__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2001__A1 _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2250_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\] _0507_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
+ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2181_ _0447_ _0353_ _0450_ _0451_ _1141_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_47_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1965_ _0739_ _0272_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1896_ tt_um_rejunity_sn76489.clk_counter\[4\] _0219_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2517_ _1109_ _1119_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2379_ _1075_ _0137_ _0603_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2448_ _0623_ _0644_ _0653_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2059__A1 _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__A1 _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\] _1022_ _1169_ _1170_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2470__A1 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2416__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _1098_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2302_ _0550_ _1010_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input9_I io_in_1[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2164_ _0433_ _0436_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2233_ _0489_ _0493_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_48_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2095_ _0375_ _0379_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1879_ _1097_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1948_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\] _0260_ _0261_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_sn76489_29 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_22_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2452__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2582__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2443__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1802_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\] _0998_ _1212_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1733_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\] _0972_ _1156_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1595_ _1013_ _1039_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1664_ _1101_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2216_ _0474_ _0479_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2147_ _0417_ _0421_ _0381_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1895__I _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2078_ _0365_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1380_ _0785_ _0827_ _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_10_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2001_ _0224_ _0302_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1716_ _1140_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2696_ _0170_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1578_ _1019_ _1022_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2479__C _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1647_ _1081_ _1082_ _1086_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xrebuffer20 _0841_ net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2620__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2550_ _0024_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1432_ _0860_ _0878_ _0880_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2481_ _0637_ _0672_ _0678_ _0676_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1363_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _0812_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1501_ _0947_ _0744_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1294_ _0731_ _0735_ _0740_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_2679_ _0153_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2643__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2419__I _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1981_ _0286_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2602_ _0076_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2533_ _0007_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1993__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1415_ _0830_ _0848_ _0863_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2464_ _0634_ _0661_ _0666_ _0665_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2395_ _1096_ _0611_ _0616_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1346_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\] _0795_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1277_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _0717_ _0726_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2064__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2180_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] _0448_ _0444_ _0451_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1895_ _1210_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1964_ tt_um_rejunity_sn76489.control_noise\[0\]\[2\] tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
+ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2447_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\] _0648_ _0652_ _0653_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2516_ _0283_ _1109_ _1119_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2378_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\] _0589_ _0132_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\]
+ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1329_ _0777_ _0768_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XTAP_TAPCELL_ROW_3_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2301_ tt_um_rejunity_sn76489.pwm.accumulator\[7\] _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1680_ _1096_ _1111_ _1114_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2704__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2163_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\] _0426_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
+ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2232_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\] _0492_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
+ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2094_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\] _0373_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
+ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1878_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\] _1052_ _0208_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1947_ _0237_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_22_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2452__A2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2201__B _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1732_ _1150_ _0923_ _1154_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1801_ _1210_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1663_ net5 _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_13_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1594_ _1017_ _1038_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2146_ _0417_ _0421_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2215_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\] _0478_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
+ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2077_ _0286_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\] _0299_ _0295_ _0302_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1715_ _1130_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1646_ _1083_ _1085_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2695_ _0169_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1577_ _1020_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer10 _0841_ net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer21 _0772_ net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_2129_ _0315_ _0408_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2016__B _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1394__A2 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1500_ _0732_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2480_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _0673_ _0678_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1431_ _0720_ _0879_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1362_ _0808_ _0810_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1293_ _0741_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2595__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1629_ _1043_ _1061_ _1071_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_41_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2678_ _0152_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1980_ _0285_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_15_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2601_ _0075_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xrebuffer1 _0785_ net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2532_ _0006_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2463_ _0947_ _0662_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1414_ _0855_ _0862_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1345_ _0725_ _0714_ _0792_ _0793_ _0716_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_1276_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\] _0724_ _0717_ _0725_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2394_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\] _0612_ _0615_ _0616_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2610__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_37_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1894_ _0215_ _0218_ _0219_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_28_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ _0270_ _0271_ _0235_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2515_ _0701_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2446_ _1091_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2377_ _0602_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1328_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\] _0777_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1259_ tt_um_rejunity_sn76489.chan\[2\].attenuation.in _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2656__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2300_ _0547_ _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2231_ _0478_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2093_ _0378_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2162_ _0435_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1877_ _0194_ _0207_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2529__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1946_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\] _0252_ _0259_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2679__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2429_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\] _0635_ _0638_ _0641_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1800_ _1140_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1731_ _1149_ _1153_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1662_ _1096_ _1088_ _1100_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1593_ _1024_ _1037_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2214_ _0465_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2145_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\] _0413_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
+ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2076_ _0359_ _0363_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1929_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\] _0238_ _0247_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_34_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2189__A2 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1607__I _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1576_ _1019_ _1020_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1714_ _1137_ _1138_ _1139_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1645_ net11 _1084_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_6_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2694_ _0168_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xrebuffer11 _0759_ net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2059_ _0315_ _0349_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2128_ _0402_ _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1394__A3 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1606__A1 _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1430_ _0711_ _0709_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1361_ _0751_ _0806_ _0809_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1292_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _0729_ _0741_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_53_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1628_ _1044_ _1060_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1559_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _0735_ _1005_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2677_ _0151_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2078__I _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_37_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xrebuffer2 _0569_ net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2600_ _0074_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_21_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2252__A1 _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2562__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1413_ _0856_ _0857_ _0859_ _0861_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2462_ _0632_ _0661_ _0664_ _0665_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2531_ _0005_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2393_ _0614_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1818__A1 _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1344_ _0720_ _0725_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1275_ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2491__A1 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output16_I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2585__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1512__A3 _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\] _0237_ _0271_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1893_ tt_um_rejunity_sn76489.clk_counter\[3\] _0217_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2376_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\] _1079_ _0590_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\]
+ _0581_ net25 _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2130__B _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2445_ _0620_ _0644_ _0651_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2514_ tt_um_rejunity_sn76489.latch_control_reg\[2\] _0698_ _1086_ _1228_ _0701_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1327_ _0773_ _0774_ _0775_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__2464__A1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2091__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2455__A1 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2230_ _0491_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2161_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\] _0425_ _0433_ _0434_ _0419_
+ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2092_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\] _0362_ _0375_ _0376_ _0377_
+ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_0_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2125__B _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1945_ _0257_ _0258_ _0251_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1876_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\] _1052_ _0206_ _0207_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_43_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2359_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\] _0000_ _0132_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\]
+ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_39_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2428_ _0620_ _0630_ _0640_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2623__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2428__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1592_ _1026_ _1027_ _1036_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1730_ _1150_ _0923_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1661_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\] _1089_ _1099_ _1100_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input7_I io_in_1[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2144_ _0420_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2213_ _0477_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1678__C _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2075_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\] _0358_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
+ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1859_ _1257_ _1258_ _1238_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1928_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\] _0241_ _0246_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1633__A2 _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1713_ _1137_ _1138_ _1127_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2669__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1575_ _0877_ _0727_ _0860_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2693_ _0167_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1644_ net10 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xrebuffer12 _0885_ net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2127_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\] _0406_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
+ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2058_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\] _1063_ _0348_ _0349_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_16_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1360_ _0765_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1291_ _0736_ _0737_ _0739_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2676_ _0150_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1627_ _1067_ _1069_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1558_ _0859_ _0793_ _1003_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1489_ _0813_ _0834_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2261__A2 _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer3 _1012_ net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2530_ _0004_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2707__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1412_ _0721_ _0860_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1343_ _0710_ _0723_ _0718_ _0720_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2461_ _1092_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2392_ _1097_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1274_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\] _0723_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2243__A2 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2659_ _0133_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2482__A2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ tt_um_rejunity_sn76489.clk_counter\[3\] _0217_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1961_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\] _0263_ _0270_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2513_ _0623_ _0698_ _0700_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2375_ _0601_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1326_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2444_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\] _0648_ _0646_ _0651_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_49_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2552__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2160_ _0428_ _0432_ _0429_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2391__A1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2091_ _1227_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1875_ _0201_ _0204_ _0205_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2192__I _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1944_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\] _0249_ _0258_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2427_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\] _0635_ _0638_ _0640_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2289_ _0537_ _0538_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2358_ _0591_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_39_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1309_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\] _0758_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1591_ _1034_ _1035_ _0995_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ _1098_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2143_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\] _0384_ _0417_ _0418_ _0419_
+ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2212_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\] _0468_ _0474_ _0476_ _0439_
+ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2074_ _0361_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1858_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\] _0997_ _1258_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1927_ _0244_ _0245_ _0240_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1789_ _1196_ _1032_ _1200_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_50_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1397__A2 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1712_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\] _0870_ _1138_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2692_ _0166_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1643_ net9 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1574_ _1018_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2057_ _0346_ _0347_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer13 _0919_ net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2126_ _0287_ _0389_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2613__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1290_ _0738_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2636__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1626_ _1053_ _1068_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2675_ _0149_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1557_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _0719_ _1003_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1488_ net61 _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1297__A1 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2109_ _0386_ _0390_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2460_ _0733_ _0662_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer4 _0845_ net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_23_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1342_ _0787_ _0790_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1273_ _0709_ _0714_ _0719_ _0721_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_1411_ _0710_ _0711_ _0713_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2391_ _0605_ _0611_ _0613_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1609_ _1051_ _1052_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2658_ _0132_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2589_ _0063_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1891_ _0215_ _0216_ _0217_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_28_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1960_ _0268_ _0269_ _0262_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1984__A2 _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2443_ _0637_ _0643_ _0650_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2512_ _0606_ _1085_ _0652_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2374_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\] _0596_ _0590_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\]
+ _0597_ net24 _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_1325_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _0774_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1975__A2 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2512__B _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2090_ _0370_ _0374_ _0366_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1642__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1874_ _0203_ _1026_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_31_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1943_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\] _0252_ _0257_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2426_ _0637_ _0629_ _0639_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2357_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\] _0589_ _0521_ _0585_
+ _0590_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\] _0591_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_TAPCELL_ROW_39_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2288_ _0209_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1308_ _0754_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1645__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ _0999_ _0992_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2142_ _1227_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2211_ _0470_ _0473_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2073_ _0287_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1788_ _1195_ _1199_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1857_ _1255_ _1256_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1926_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\] _0238_ _0245_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1866__A1 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2542__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2692__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2409_ tt_um_rejunity_sn76489.latch_control_reg\[1\] _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2288__I _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2565__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1711_ _1133_ _1135_ _1136_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_6_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2691_ _0165_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1642_ net7 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1573_ _0852_ _0873_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2056_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\] _1018_ _0343_ _0347_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xrebuffer14 net19 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2125_ _0402_ _0405_ _0213_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1909_ _0230_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2588__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2504__C _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ _0148_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1625_ _1050_ _1058_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1556_ _0996_ _1001_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_41_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1487_ net51 _0806_ _0934_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2039_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\] _0973_ _0333_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2246__A1 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2108_ _0386_ _0390_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_17_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1410_ _0856_ _0857_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xrebuffer5 net44 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1272_ _0720_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1341_ _0788_ _0789_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2390_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\] _0612_ _0539_ _0613_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2400__A1 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2657_ _0131_ clknet_4_15_0_wb_clk_i net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1608_ _1049_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1539_ _0983_ _0984_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2588_ _0062_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2626__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1890_ _0212_ tt_um_rejunity_sn76489.clk_counter\[1\] tt_um_rejunity_sn76489.clk_counter\[2\]
+ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2373_ _0600_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2442_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\] _0648_ _0646_ _0650_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2511_ _0620_ _0698_ _0699_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1324_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _0773_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1994__B _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2709_ _0183_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1942_ _0255_ _0256_ _0251_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1873_ _0203_ _1026_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2356_ _0574_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2425_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\] _0635_ _0638_ _0639_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2287_ tt_um_rejunity_sn76489.pwm.accumulator\[5\] net20 _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_39_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1307_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1989__B _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2210_ _0365_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1627__A2 _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_28_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2141_ _0414_ _0416_ _0381_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2072_ _0354_ _0360_ _0213_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2052__A2 _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1925_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\] _0241_ _0244_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1787_ _1196_ _1032_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1856_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\] _1028_ _1252_ _1256_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_12_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2339_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\] _0578_ _0579_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2408_ _0623_ _0612_ _0625_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2062__C _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2253__B _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1572_ _1002_ _1008_ _1016_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1710_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\] _0822_ _1136_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2690_ _0164_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1641_ net8 _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input5_I io_in_1[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2124_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\] _0403_ _0404_ _0405_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xrebuffer15 _1072_ net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2055_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\] _1018_ _0346_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1839_ _1240_ _1241_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1908_ tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
+ _0229_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2532__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2248__B _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2682__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2673_ _0147_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1624_ _1065_ _1066_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1555_ _0967_ _0969_ _1000_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2191__A1 _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1486_ _0809_ net60 net44 _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2107_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\] _0389_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
+ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2038_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\] _0973_ _0332_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1997__B _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2555__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1340_ _0743_ _0748_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xrebuffer6 _0845_ net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__A1 _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1271_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _0708_ _0720_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_46_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1987__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2656_ _0130_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1607_ _1048_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1538_ _0957_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1469_ _0917_ _0908_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2587_ _0061_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1902__A1 _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2510_ _0607_ _0698_ _0652_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2372_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\] _0596_ _0590_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\]
+ _0597_ net23 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_1323_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _0771_ _0769_ _0772_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2441_ _0634_ _0643_ _0649_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2708_ _0182_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2137__A1 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2639_ _0113_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2256__B _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2100__I _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1872_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\] _0203_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1941_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\] _0249_ _0256_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2355_ _1079_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2286_ _0536_ net56 _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1306_ tt_um_rejunity_sn76489.chan\[0\].attenuation.in _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_2424_ _0614_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2616__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2140_ _0414_ _0416_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2639__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2071_ _0355_ _0359_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1855_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\] _1028_ _1255_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1924_ _0242_ _0243_ _0240_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1786_ _1195_ _1197_ _1198_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2269_ _0520_ _0522_ _0460_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2338_ _0573_ _0577_ _0578_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2407_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\] _0617_ _0624_ _0625_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1571_ _1014_ _1015_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1640_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\] _1080_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1664__I _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer16 _0534_ net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_2123_ _0281_ _0398_ _0401_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2054_ _0343_ _0344_ _0345_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1838_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\] _0892_ _1236_ _1241_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1907_ _0228_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1574__I _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1769_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\] _0818_ _1184_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1659__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2672_ _0146_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1623_ _1047_ _1059_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1554_ _0999_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1485_ _0829_ _0912_ _0911_ _0915_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_1_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

