magic
tech gf180mcuD
magscale 1 5
timestamp 1702416648
<< obsm1 >>
rect 672 1538 114296 113385
<< metal2 >>
rect 1904 114600 1960 115000
rect 5376 114600 5432 115000
rect 8848 114600 8904 115000
rect 12320 114600 12376 115000
rect 15792 114600 15848 115000
rect 19264 114600 19320 115000
rect 22736 114600 22792 115000
rect 26208 114600 26264 115000
rect 29680 114600 29736 115000
rect 33152 114600 33208 115000
rect 36624 114600 36680 115000
rect 40096 114600 40152 115000
rect 43568 114600 43624 115000
rect 47040 114600 47096 115000
rect 50512 114600 50568 115000
rect 53984 114600 54040 115000
rect 57456 114600 57512 115000
rect 60928 114600 60984 115000
rect 64400 114600 64456 115000
rect 67872 114600 67928 115000
rect 71344 114600 71400 115000
rect 74816 114600 74872 115000
rect 78288 114600 78344 115000
rect 81760 114600 81816 115000
rect 85232 114600 85288 115000
rect 88704 114600 88760 115000
rect 92176 114600 92232 115000
rect 95648 114600 95704 115000
rect 99120 114600 99176 115000
rect 102592 114600 102648 115000
rect 106064 114600 106120 115000
rect 109536 114600 109592 115000
rect 113008 114600 113064 115000
rect 1904 0 1960 400
rect 5376 0 5432 400
rect 8848 0 8904 400
rect 12320 0 12376 400
rect 15792 0 15848 400
rect 19264 0 19320 400
rect 22736 0 22792 400
rect 26208 0 26264 400
rect 29680 0 29736 400
rect 33152 0 33208 400
rect 36624 0 36680 400
rect 40096 0 40152 400
rect 43568 0 43624 400
rect 47040 0 47096 400
rect 50512 0 50568 400
rect 53984 0 54040 400
rect 57456 0 57512 400
rect 60928 0 60984 400
rect 64400 0 64456 400
rect 67872 0 67928 400
rect 71344 0 71400 400
rect 74816 0 74872 400
rect 78288 0 78344 400
rect 81760 0 81816 400
rect 85232 0 85288 400
rect 88704 0 88760 400
rect 92176 0 92232 400
rect 95648 0 95704 400
rect 99120 0 99176 400
rect 102592 0 102648 400
rect 106064 0 106120 400
rect 109536 0 109592 400
rect 113008 0 113064 400
<< obsm2 >>
rect 406 114570 1874 114674
rect 1990 114570 5346 114674
rect 5462 114570 8818 114674
rect 8934 114570 12290 114674
rect 12406 114570 15762 114674
rect 15878 114570 19234 114674
rect 19350 114570 22706 114674
rect 22822 114570 26178 114674
rect 26294 114570 29650 114674
rect 29766 114570 33122 114674
rect 33238 114570 36594 114674
rect 36710 114570 40066 114674
rect 40182 114570 43538 114674
rect 43654 114570 47010 114674
rect 47126 114570 50482 114674
rect 50598 114570 53954 114674
rect 54070 114570 57426 114674
rect 57542 114570 60898 114674
rect 61014 114570 64370 114674
rect 64486 114570 67842 114674
rect 67958 114570 71314 114674
rect 71430 114570 74786 114674
rect 74902 114570 78258 114674
rect 78374 114570 81730 114674
rect 81846 114570 85202 114674
rect 85318 114570 88674 114674
rect 88790 114570 92146 114674
rect 92262 114570 95618 114674
rect 95734 114570 99090 114674
rect 99206 114570 102562 114674
rect 102678 114570 106034 114674
rect 106150 114570 109506 114674
rect 109622 114570 112978 114674
rect 113094 114570 114170 114674
rect 406 430 114170 114570
rect 406 121 1874 430
rect 1990 121 5346 430
rect 5462 121 8818 430
rect 8934 121 12290 430
rect 12406 121 15762 430
rect 15878 121 19234 430
rect 19350 121 22706 430
rect 22822 121 26178 430
rect 26294 121 29650 430
rect 29766 121 33122 430
rect 33238 121 36594 430
rect 36710 121 40066 430
rect 40182 121 43538 430
rect 43654 121 47010 430
rect 47126 121 50482 430
rect 50598 121 53954 430
rect 54070 121 57426 430
rect 57542 121 60898 430
rect 61014 121 64370 430
rect 64486 121 67842 430
rect 67958 121 71314 430
rect 71430 121 74786 430
rect 74902 121 78258 430
rect 78374 121 81730 430
rect 81846 121 85202 430
rect 85318 121 88674 430
rect 88790 121 92146 430
rect 92262 121 95618 430
rect 95734 121 99090 430
rect 99206 121 102562 430
rect 102678 121 106034 430
rect 106150 121 109506 430
rect 109622 121 112978 430
rect 113094 121 114170 430
<< metal3 >>
rect 0 111888 400 111944
rect 0 108864 400 108920
rect 0 105840 400 105896
rect 0 102816 400 102872
rect 0 99792 400 99848
rect 0 96768 400 96824
rect 0 93744 400 93800
rect 0 90720 400 90776
rect 0 87696 400 87752
rect 0 84672 400 84728
rect 0 81648 400 81704
rect 0 78624 400 78680
rect 0 75600 400 75656
rect 0 72576 400 72632
rect 0 69552 400 69608
rect 0 66528 400 66584
rect 0 63504 400 63560
rect 0 60480 400 60536
rect 0 57456 400 57512
rect 0 54432 400 54488
rect 0 51408 400 51464
rect 0 48384 400 48440
rect 0 45360 400 45416
rect 0 42336 400 42392
rect 0 39312 400 39368
rect 0 36288 400 36344
rect 0 33264 400 33320
rect 0 30240 400 30296
rect 0 27216 400 27272
rect 0 24192 400 24248
rect 0 21168 400 21224
rect 0 18144 400 18200
rect 0 15120 400 15176
rect 0 12096 400 12152
rect 0 9072 400 9128
rect 0 6048 400 6104
rect 0 3024 400 3080
<< obsm3 >>
rect 400 111974 114175 113610
rect 430 111858 114175 111974
rect 400 108950 114175 111858
rect 430 108834 114175 108950
rect 400 105926 114175 108834
rect 430 105810 114175 105926
rect 400 102902 114175 105810
rect 430 102786 114175 102902
rect 400 99878 114175 102786
rect 430 99762 114175 99878
rect 400 96854 114175 99762
rect 430 96738 114175 96854
rect 400 93830 114175 96738
rect 430 93714 114175 93830
rect 400 90806 114175 93714
rect 430 90690 114175 90806
rect 400 87782 114175 90690
rect 430 87666 114175 87782
rect 400 84758 114175 87666
rect 430 84642 114175 84758
rect 400 81734 114175 84642
rect 430 81618 114175 81734
rect 400 78710 114175 81618
rect 430 78594 114175 78710
rect 400 75686 114175 78594
rect 430 75570 114175 75686
rect 400 72662 114175 75570
rect 430 72546 114175 72662
rect 400 69638 114175 72546
rect 430 69522 114175 69638
rect 400 66614 114175 69522
rect 430 66498 114175 66614
rect 400 63590 114175 66498
rect 430 63474 114175 63590
rect 400 60566 114175 63474
rect 430 60450 114175 60566
rect 400 57542 114175 60450
rect 430 57426 114175 57542
rect 400 54518 114175 57426
rect 430 54402 114175 54518
rect 400 51494 114175 54402
rect 430 51378 114175 51494
rect 400 48470 114175 51378
rect 430 48354 114175 48470
rect 400 45446 114175 48354
rect 430 45330 114175 45446
rect 400 42422 114175 45330
rect 430 42306 114175 42422
rect 400 39398 114175 42306
rect 430 39282 114175 39398
rect 400 36374 114175 39282
rect 430 36258 114175 36374
rect 400 33350 114175 36258
rect 430 33234 114175 33350
rect 400 30326 114175 33234
rect 430 30210 114175 30326
rect 400 27302 114175 30210
rect 430 27186 114175 27302
rect 400 24278 114175 27186
rect 430 24162 114175 24278
rect 400 21254 114175 24162
rect 430 21138 114175 21254
rect 400 18230 114175 21138
rect 430 18114 114175 18230
rect 400 15206 114175 18114
rect 430 15090 114175 15206
rect 400 12182 114175 15090
rect 430 12066 114175 12182
rect 400 9158 114175 12066
rect 430 9042 114175 9158
rect 400 6134 114175 9042
rect 430 6018 114175 6134
rect 400 3110 114175 6018
rect 430 2994 114175 3110
rect 400 126 114175 2994
<< metal4 >>
rect 2224 1538 2384 113318
rect 9904 1538 10064 113318
rect 17584 1538 17744 113318
rect 25264 1538 25424 113318
rect 32944 1538 33104 113318
rect 40624 1538 40784 113318
rect 48304 1538 48464 113318
rect 55984 1538 56144 113318
rect 63664 1538 63824 113318
rect 71344 1538 71504 113318
rect 79024 1538 79184 113318
rect 86704 1538 86864 113318
rect 94384 1538 94544 113318
rect 102064 1538 102224 113318
rect 109744 1538 109904 113318
<< obsm4 >>
rect 966 113348 113274 113615
rect 966 1508 2194 113348
rect 2414 1508 9874 113348
rect 10094 1508 17554 113348
rect 17774 1508 25234 113348
rect 25454 1508 32914 113348
rect 33134 1508 40594 113348
rect 40814 1508 48274 113348
rect 48494 1508 55954 113348
rect 56174 1508 63634 113348
rect 63854 1508 71314 113348
rect 71534 1508 78994 113348
rect 79214 1508 86674 113348
rect 86894 1508 94354 113348
rect 94574 1508 102034 113348
rect 102254 1508 109714 113348
rect 109934 1508 113274 113348
rect 966 233 113274 1508
<< labels >>
rlabel metal3 s 0 9072 400 9128 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 12096 400 12152 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 0 15120 400 15176 6 io_in[0]
port 3 nsew signal input
rlabel metal3 s 0 45360 400 45416 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 0 48384 400 48440 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 0 51408 400 51464 6 io_in[12]
port 6 nsew signal input
rlabel metal3 s 0 54432 400 54488 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 0 57456 400 57512 6 io_in[14]
port 8 nsew signal input
rlabel metal3 s 0 60480 400 60536 6 io_in[15]
port 9 nsew signal input
rlabel metal3 s 0 63504 400 63560 6 io_in[16]
port 10 nsew signal input
rlabel metal3 s 0 66528 400 66584 6 io_in[17]
port 11 nsew signal input
rlabel metal3 s 0 69552 400 69608 6 io_in[18]
port 12 nsew signal input
rlabel metal3 s 0 72576 400 72632 6 io_in[19]
port 13 nsew signal input
rlabel metal3 s 0 18144 400 18200 6 io_in[1]
port 14 nsew signal input
rlabel metal3 s 0 75600 400 75656 6 io_in[20]
port 15 nsew signal input
rlabel metal3 s 0 78624 400 78680 6 io_in[21]
port 16 nsew signal input
rlabel metal3 s 0 81648 400 81704 6 io_in[22]
port 17 nsew signal input
rlabel metal3 s 0 84672 400 84728 6 io_in[23]
port 18 nsew signal input
rlabel metal3 s 0 87696 400 87752 6 io_in[24]
port 19 nsew signal input
rlabel metal3 s 0 90720 400 90776 6 io_in[25]
port 20 nsew signal input
rlabel metal3 s 0 93744 400 93800 6 io_in[26]
port 21 nsew signal input
rlabel metal3 s 0 96768 400 96824 6 io_in[27]
port 22 nsew signal input
rlabel metal3 s 0 99792 400 99848 6 io_in[28]
port 23 nsew signal input
rlabel metal3 s 0 102816 400 102872 6 io_in[29]
port 24 nsew signal input
rlabel metal3 s 0 21168 400 21224 6 io_in[2]
port 25 nsew signal input
rlabel metal3 s 0 105840 400 105896 6 io_in[30]
port 26 nsew signal input
rlabel metal3 s 0 108864 400 108920 6 io_in[31]
port 27 nsew signal input
rlabel metal3 s 0 111888 400 111944 6 io_in[32]
port 28 nsew signal input
rlabel metal3 s 0 24192 400 24248 6 io_in[3]
port 29 nsew signal input
rlabel metal3 s 0 27216 400 27272 6 io_in[4]
port 30 nsew signal input
rlabel metal3 s 0 30240 400 30296 6 io_in[5]
port 31 nsew signal input
rlabel metal3 s 0 33264 400 33320 6 io_in[6]
port 32 nsew signal input
rlabel metal3 s 0 36288 400 36344 6 io_in[7]
port 33 nsew signal input
rlabel metal3 s 0 39312 400 39368 6 io_in[8]
port 34 nsew signal input
rlabel metal3 s 0 42336 400 42392 6 io_in[9]
port 35 nsew signal input
rlabel metal2 s 1904 114600 1960 115000 6 io_oeb[0]
port 36 nsew signal output
rlabel metal2 s 36624 114600 36680 115000 6 io_oeb[10]
port 37 nsew signal output
rlabel metal2 s 40096 114600 40152 115000 6 io_oeb[11]
port 38 nsew signal output
rlabel metal2 s 43568 114600 43624 115000 6 io_oeb[12]
port 39 nsew signal output
rlabel metal2 s 47040 114600 47096 115000 6 io_oeb[13]
port 40 nsew signal output
rlabel metal2 s 50512 114600 50568 115000 6 io_oeb[14]
port 41 nsew signal output
rlabel metal2 s 53984 114600 54040 115000 6 io_oeb[15]
port 42 nsew signal output
rlabel metal2 s 57456 114600 57512 115000 6 io_oeb[16]
port 43 nsew signal output
rlabel metal2 s 60928 114600 60984 115000 6 io_oeb[17]
port 44 nsew signal output
rlabel metal2 s 64400 114600 64456 115000 6 io_oeb[18]
port 45 nsew signal output
rlabel metal2 s 67872 114600 67928 115000 6 io_oeb[19]
port 46 nsew signal output
rlabel metal2 s 5376 114600 5432 115000 6 io_oeb[1]
port 47 nsew signal output
rlabel metal2 s 71344 114600 71400 115000 6 io_oeb[20]
port 48 nsew signal output
rlabel metal2 s 74816 114600 74872 115000 6 io_oeb[21]
port 49 nsew signal output
rlabel metal2 s 78288 114600 78344 115000 6 io_oeb[22]
port 50 nsew signal output
rlabel metal2 s 81760 114600 81816 115000 6 io_oeb[23]
port 51 nsew signal output
rlabel metal2 s 85232 114600 85288 115000 6 io_oeb[24]
port 52 nsew signal output
rlabel metal2 s 88704 114600 88760 115000 6 io_oeb[25]
port 53 nsew signal output
rlabel metal2 s 92176 114600 92232 115000 6 io_oeb[26]
port 54 nsew signal output
rlabel metal2 s 95648 114600 95704 115000 6 io_oeb[27]
port 55 nsew signal output
rlabel metal2 s 99120 114600 99176 115000 6 io_oeb[28]
port 56 nsew signal output
rlabel metal2 s 102592 114600 102648 115000 6 io_oeb[29]
port 57 nsew signal output
rlabel metal2 s 8848 114600 8904 115000 6 io_oeb[2]
port 58 nsew signal output
rlabel metal2 s 106064 114600 106120 115000 6 io_oeb[30]
port 59 nsew signal output
rlabel metal2 s 109536 114600 109592 115000 6 io_oeb[31]
port 60 nsew signal output
rlabel metal2 s 113008 114600 113064 115000 6 io_oeb[32]
port 61 nsew signal output
rlabel metal2 s 12320 114600 12376 115000 6 io_oeb[3]
port 62 nsew signal output
rlabel metal2 s 15792 114600 15848 115000 6 io_oeb[4]
port 63 nsew signal output
rlabel metal2 s 19264 114600 19320 115000 6 io_oeb[5]
port 64 nsew signal output
rlabel metal2 s 22736 114600 22792 115000 6 io_oeb[6]
port 65 nsew signal output
rlabel metal2 s 26208 114600 26264 115000 6 io_oeb[7]
port 66 nsew signal output
rlabel metal2 s 29680 114600 29736 115000 6 io_oeb[8]
port 67 nsew signal output
rlabel metal2 s 33152 114600 33208 115000 6 io_oeb[9]
port 68 nsew signal output
rlabel metal2 s 1904 0 1960 400 6 io_out[0]
port 69 nsew signal output
rlabel metal2 s 36624 0 36680 400 6 io_out[10]
port 70 nsew signal output
rlabel metal2 s 40096 0 40152 400 6 io_out[11]
port 71 nsew signal output
rlabel metal2 s 43568 0 43624 400 6 io_out[12]
port 72 nsew signal output
rlabel metal2 s 47040 0 47096 400 6 io_out[13]
port 73 nsew signal output
rlabel metal2 s 50512 0 50568 400 6 io_out[14]
port 74 nsew signal output
rlabel metal2 s 53984 0 54040 400 6 io_out[15]
port 75 nsew signal output
rlabel metal2 s 57456 0 57512 400 6 io_out[16]
port 76 nsew signal output
rlabel metal2 s 60928 0 60984 400 6 io_out[17]
port 77 nsew signal output
rlabel metal2 s 64400 0 64456 400 6 io_out[18]
port 78 nsew signal output
rlabel metal2 s 67872 0 67928 400 6 io_out[19]
port 79 nsew signal output
rlabel metal2 s 5376 0 5432 400 6 io_out[1]
port 80 nsew signal output
rlabel metal2 s 71344 0 71400 400 6 io_out[20]
port 81 nsew signal output
rlabel metal2 s 74816 0 74872 400 6 io_out[21]
port 82 nsew signal output
rlabel metal2 s 78288 0 78344 400 6 io_out[22]
port 83 nsew signal output
rlabel metal2 s 81760 0 81816 400 6 io_out[23]
port 84 nsew signal output
rlabel metal2 s 85232 0 85288 400 6 io_out[24]
port 85 nsew signal output
rlabel metal2 s 88704 0 88760 400 6 io_out[25]
port 86 nsew signal output
rlabel metal2 s 92176 0 92232 400 6 io_out[26]
port 87 nsew signal output
rlabel metal2 s 95648 0 95704 400 6 io_out[27]
port 88 nsew signal output
rlabel metal2 s 99120 0 99176 400 6 io_out[28]
port 89 nsew signal output
rlabel metal2 s 102592 0 102648 400 6 io_out[29]
port 90 nsew signal output
rlabel metal2 s 8848 0 8904 400 6 io_out[2]
port 91 nsew signal output
rlabel metal2 s 106064 0 106120 400 6 io_out[30]
port 92 nsew signal output
rlabel metal2 s 109536 0 109592 400 6 io_out[31]
port 93 nsew signal output
rlabel metal2 s 113008 0 113064 400 6 io_out[32]
port 94 nsew signal output
rlabel metal2 s 12320 0 12376 400 6 io_out[3]
port 95 nsew signal output
rlabel metal2 s 15792 0 15848 400 6 io_out[4]
port 96 nsew signal output
rlabel metal2 s 19264 0 19320 400 6 io_out[5]
port 97 nsew signal output
rlabel metal2 s 22736 0 22792 400 6 io_out[6]
port 98 nsew signal output
rlabel metal2 s 26208 0 26264 400 6 io_out[7]
port 99 nsew signal output
rlabel metal2 s 29680 0 29736 400 6 io_out[8]
port 100 nsew signal output
rlabel metal2 s 33152 0 33208 400 6 io_out[9]
port 101 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 rst_n
port 102 nsew signal input
rlabel metal4 s 2224 1538 2384 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 113318 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 113318 6 vss
port 104 nsew ground bidirectional
rlabel metal3 s 0 3024 400 3080 6 wb_clk_i
port 105 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 115000 115000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 47561482
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_tholin_riscv/runs/23_12_12_19_33/results/signoff/wrapped_tholin_riscv.magic.gds
string GDS_START 593546
<< end >>

