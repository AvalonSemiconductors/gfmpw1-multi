magic
tech gf180mcuD
magscale 1 10
timestamp 1702299510
<< metal1 >>
rect 1344 42362 44576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 44576 42362
rect 1344 42276 44576 42310
rect 18286 42194 18338 42206
rect 18286 42130 18338 42142
rect 33518 42194 33570 42206
rect 33518 42130 33570 42142
rect 6190 42082 6242 42094
rect 6190 42018 6242 42030
rect 9998 42082 10050 42094
rect 9998 42018 10050 42030
rect 5070 41970 5122 41982
rect 5070 41906 5122 41918
rect 5854 41970 5906 41982
rect 5854 41906 5906 41918
rect 8878 41970 8930 41982
rect 8878 41906 8930 41918
rect 9662 41970 9714 41982
rect 13458 41918 13470 41970
rect 13522 41918 13534 41970
rect 17266 41918 17278 41970
rect 17330 41918 17342 41970
rect 21074 41918 21086 41970
rect 21138 41918 21150 41970
rect 24882 41918 24894 41970
rect 24946 41918 24958 41970
rect 30818 41918 30830 41970
rect 30882 41918 30894 41970
rect 32610 41918 32622 41970
rect 32674 41918 32686 41970
rect 36306 41918 36318 41970
rect 36370 41918 36382 41970
rect 40338 41918 40350 41970
rect 40402 41918 40414 41970
rect 9662 41906 9714 41918
rect 14478 41858 14530 41870
rect 14478 41794 14530 41806
rect 22094 41858 22146 41870
rect 22094 41794 22146 41806
rect 25902 41858 25954 41870
rect 25902 41794 25954 41806
rect 28926 41858 28978 41870
rect 28926 41794 28978 41806
rect 37326 41858 37378 41870
rect 37326 41794 37378 41806
rect 41134 41858 41186 41870
rect 41134 41794 41186 41806
rect 1344 41578 44576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 44576 41578
rect 1344 41492 44576 41526
rect 43586 41246 43598 41298
rect 43650 41246 43662 41298
rect 41570 41134 41582 41186
rect 41634 41134 41646 41186
rect 1344 40794 44576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 44576 40794
rect 1344 40708 44576 40742
rect 24334 40626 24386 40638
rect 24334 40562 24386 40574
rect 8766 40514 8818 40526
rect 5618 40462 5630 40514
rect 5682 40462 5694 40514
rect 8766 40450 8818 40462
rect 8318 40402 8370 40414
rect 16942 40402 16994 40414
rect 23662 40402 23714 40414
rect 4946 40350 4958 40402
rect 5010 40350 5022 40402
rect 9762 40350 9774 40402
rect 9826 40350 9838 40402
rect 13346 40350 13358 40402
rect 13410 40350 13422 40402
rect 17602 40350 17614 40402
rect 17666 40350 17678 40402
rect 8318 40338 8370 40350
rect 16942 40338 16994 40350
rect 23662 40338 23714 40350
rect 24110 40402 24162 40414
rect 31166 40402 31218 40414
rect 36430 40402 36482 40414
rect 27794 40350 27806 40402
rect 27858 40350 27870 40402
rect 28466 40350 28478 40402
rect 28530 40350 28542 40402
rect 33170 40350 33182 40402
rect 33234 40350 33246 40402
rect 24110 40338 24162 40350
rect 31166 40338 31218 40350
rect 36430 40338 36482 40350
rect 40462 40402 40514 40414
rect 41010 40350 41022 40402
rect 41074 40350 41086 40402
rect 40462 40338 40514 40350
rect 24222 40290 24274 40302
rect 7746 40238 7758 40290
rect 7810 40238 7822 40290
rect 10546 40238 10558 40290
rect 10610 40238 10622 40290
rect 12674 40238 12686 40290
rect 12738 40238 12750 40290
rect 14018 40238 14030 40290
rect 14082 40238 14094 40290
rect 16146 40238 16158 40290
rect 16210 40238 16222 40290
rect 18386 40238 18398 40290
rect 18450 40238 18462 40290
rect 20514 40238 20526 40290
rect 20578 40238 20590 40290
rect 24222 40226 24274 40238
rect 25454 40290 25506 40302
rect 30594 40238 30606 40290
rect 30658 40238 30670 40290
rect 33842 40238 33854 40290
rect 33906 40238 33918 40290
rect 35970 40238 35982 40290
rect 36034 40238 36046 40290
rect 41794 40238 41806 40290
rect 41858 40238 41870 40290
rect 43922 40238 43934 40290
rect 43986 40238 43998 40290
rect 25454 40226 25506 40238
rect 1344 40010 44576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 44576 40010
rect 1344 39924 44576 39958
rect 5742 39730 5794 39742
rect 4722 39678 4734 39730
rect 4786 39678 4798 39730
rect 5742 39666 5794 39678
rect 8766 39730 8818 39742
rect 18958 39730 19010 39742
rect 18386 39678 18398 39730
rect 18450 39678 18462 39730
rect 8766 39666 8818 39678
rect 18958 39666 19010 39678
rect 20190 39730 20242 39742
rect 33070 39730 33122 39742
rect 23538 39678 23550 39730
rect 23602 39678 23614 39730
rect 25666 39678 25678 39730
rect 25730 39678 25742 39730
rect 32610 39678 32622 39730
rect 32674 39678 32686 39730
rect 39218 39678 39230 39730
rect 39282 39678 39294 39730
rect 20190 39666 20242 39678
rect 33070 39666 33122 39678
rect 17950 39618 18002 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 17950 39554 18002 39566
rect 19518 39618 19570 39630
rect 26910 39618 26962 39630
rect 26450 39566 26462 39618
rect 26514 39566 26526 39618
rect 29810 39566 29822 39618
rect 29874 39566 29886 39618
rect 42018 39566 42030 39618
rect 42082 39566 42094 39618
rect 19518 39554 19570 39566
rect 26910 39554 26962 39566
rect 14590 39506 14642 39518
rect 2594 39454 2606 39506
rect 2658 39454 2670 39506
rect 14590 39442 14642 39454
rect 14926 39506 14978 39518
rect 14926 39442 14978 39454
rect 18510 39506 18562 39518
rect 18510 39442 18562 39454
rect 19070 39506 19122 39518
rect 19070 39442 19122 39454
rect 19854 39506 19906 39518
rect 30482 39454 30494 39506
rect 30546 39454 30558 39506
rect 41346 39454 41358 39506
rect 41410 39454 41422 39506
rect 19854 39442 19906 39454
rect 8878 39394 8930 39406
rect 8878 39330 8930 39342
rect 12910 39394 12962 39406
rect 12910 39330 12962 39342
rect 16382 39394 16434 39406
rect 16382 39330 16434 39342
rect 18286 39394 18338 39406
rect 18286 39330 18338 39342
rect 18846 39394 18898 39406
rect 18846 39330 18898 39342
rect 20078 39394 20130 39406
rect 20078 39330 20130 39342
rect 20302 39394 20354 39406
rect 20302 39330 20354 39342
rect 38894 39394 38946 39406
rect 38894 39330 38946 39342
rect 1344 39226 44576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 44576 39226
rect 1344 39140 44576 39174
rect 20302 39058 20354 39070
rect 20302 38994 20354 39006
rect 24782 39058 24834 39070
rect 24782 38994 24834 39006
rect 25790 39058 25842 39070
rect 38334 39058 38386 39070
rect 26450 39006 26462 39058
rect 26514 39006 26526 39058
rect 25790 38994 25842 39006
rect 38334 38994 38386 39006
rect 41358 39058 41410 39070
rect 41358 38994 41410 39006
rect 41470 39058 41522 39070
rect 41470 38994 41522 39006
rect 41694 39058 41746 39070
rect 41694 38994 41746 39006
rect 20526 38946 20578 38958
rect 20526 38882 20578 38894
rect 24110 38946 24162 38958
rect 24110 38882 24162 38894
rect 24446 38946 24498 38958
rect 24446 38882 24498 38894
rect 24558 38946 24610 38958
rect 24558 38882 24610 38894
rect 27134 38946 27186 38958
rect 27134 38882 27186 38894
rect 39902 38946 39954 38958
rect 39902 38882 39954 38894
rect 20190 38834 20242 38846
rect 20190 38770 20242 38782
rect 25566 38834 25618 38846
rect 25566 38770 25618 38782
rect 25790 38834 25842 38846
rect 25790 38770 25842 38782
rect 26126 38834 26178 38846
rect 27246 38834 27298 38846
rect 37774 38834 37826 38846
rect 39790 38834 39842 38846
rect 26674 38782 26686 38834
rect 26738 38782 26750 38834
rect 37538 38782 37550 38834
rect 37602 38782 37614 38834
rect 38098 38782 38110 38834
rect 38162 38782 38174 38834
rect 26126 38770 26178 38782
rect 27246 38770 27298 38782
rect 37774 38770 37826 38782
rect 39790 38770 39842 38782
rect 40126 38834 40178 38846
rect 40126 38770 40178 38782
rect 40798 38834 40850 38846
rect 41122 38782 41134 38834
rect 41186 38782 41198 38834
rect 41906 38782 41918 38834
rect 41970 38782 41982 38834
rect 42130 38782 42142 38834
rect 42194 38782 42206 38834
rect 40798 38770 40850 38782
rect 23886 38722 23938 38734
rect 38782 38722 38834 38734
rect 34626 38670 34638 38722
rect 34690 38670 34702 38722
rect 36754 38670 36766 38722
rect 36818 38670 36830 38722
rect 41794 38670 41806 38722
rect 41858 38670 41870 38722
rect 23886 38658 23938 38670
rect 38782 38658 38834 38670
rect 23550 38610 23602 38622
rect 23550 38546 23602 38558
rect 37998 38610 38050 38622
rect 37998 38546 38050 38558
rect 1344 38442 44576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 44576 38442
rect 1344 38356 44576 38390
rect 20414 38274 20466 38286
rect 20414 38210 20466 38222
rect 24446 38274 24498 38286
rect 25554 38222 25566 38274
rect 25618 38222 25630 38274
rect 24446 38210 24498 38222
rect 5742 38162 5794 38174
rect 23550 38162 23602 38174
rect 5058 38110 5070 38162
rect 5122 38110 5134 38162
rect 7746 38110 7758 38162
rect 7810 38110 7822 38162
rect 16594 38110 16606 38162
rect 16658 38110 16670 38162
rect 18722 38110 18734 38162
rect 18786 38110 18798 38162
rect 25778 38110 25790 38162
rect 25842 38110 25854 38162
rect 5742 38098 5794 38110
rect 23550 38098 23602 38110
rect 11118 38050 11170 38062
rect 24110 38050 24162 38062
rect 2258 37998 2270 38050
rect 2322 37998 2334 38050
rect 10546 37998 10558 38050
rect 10610 37998 10622 38050
rect 15810 37998 15822 38050
rect 15874 37998 15886 38050
rect 11118 37986 11170 37998
rect 24110 37986 24162 37998
rect 24222 38050 24274 38062
rect 24222 37986 24274 37998
rect 37438 38050 37490 38062
rect 37438 37986 37490 37998
rect 40574 38050 40626 38062
rect 40574 37986 40626 37998
rect 20078 37938 20130 37950
rect 2930 37886 2942 37938
rect 2994 37886 3006 37938
rect 9874 37886 9886 37938
rect 9938 37886 9950 37938
rect 19730 37886 19742 37938
rect 19794 37886 19806 37938
rect 20078 37874 20130 37886
rect 20526 37938 20578 37950
rect 20526 37874 20578 37886
rect 23662 37938 23714 37950
rect 37102 37938 37154 37950
rect 26002 37886 26014 37938
rect 26066 37886 26078 37938
rect 23662 37874 23714 37886
rect 37102 37874 37154 37886
rect 37214 37938 37266 37950
rect 37214 37874 37266 37886
rect 40238 37938 40290 37950
rect 40238 37874 40290 37886
rect 40350 37938 40402 37950
rect 40350 37874 40402 37886
rect 41022 37938 41074 37950
rect 41022 37874 41074 37886
rect 41134 37938 41186 37950
rect 41134 37874 41186 37886
rect 41358 37938 41410 37950
rect 41358 37874 41410 37886
rect 19182 37826 19234 37838
rect 19182 37762 19234 37774
rect 23438 37826 23490 37838
rect 23438 37762 23490 37774
rect 26574 37826 26626 37838
rect 26574 37762 26626 37774
rect 1344 37658 44576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 44576 37658
rect 1344 37572 44576 37606
rect 4622 37490 4674 37502
rect 4622 37426 4674 37438
rect 5070 37490 5122 37502
rect 5070 37426 5122 37438
rect 14254 37490 14306 37502
rect 14254 37426 14306 37438
rect 20414 37490 20466 37502
rect 20414 37426 20466 37438
rect 24110 37490 24162 37502
rect 41358 37490 41410 37502
rect 25218 37438 25230 37490
rect 25282 37438 25294 37490
rect 24110 37426 24162 37438
rect 41358 37426 41410 37438
rect 41134 37378 41186 37390
rect 41134 37314 41186 37326
rect 5630 37266 5682 37278
rect 20750 37266 20802 37278
rect 4386 37214 4398 37266
rect 4450 37214 4462 37266
rect 10994 37214 11006 37266
rect 11058 37214 11070 37266
rect 5630 37202 5682 37214
rect 20750 37202 20802 37214
rect 41022 37266 41074 37278
rect 41022 37202 41074 37214
rect 5182 37154 5234 37166
rect 25790 37154 25842 37166
rect 11666 37102 11678 37154
rect 11730 37102 11742 37154
rect 13794 37102 13806 37154
rect 13858 37102 13870 37154
rect 5182 37090 5234 37102
rect 25790 37090 25842 37102
rect 4734 37042 4786 37054
rect 4734 36978 4786 36990
rect 25566 37042 25618 37054
rect 25566 36978 25618 36990
rect 1344 36874 44576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 44576 36874
rect 1344 36788 44576 36822
rect 7422 36706 7474 36718
rect 40798 36706 40850 36718
rect 21298 36654 21310 36706
rect 21362 36654 21374 36706
rect 7422 36642 7474 36654
rect 40798 36642 40850 36654
rect 6974 36594 7026 36606
rect 6974 36530 7026 36542
rect 7758 36482 7810 36494
rect 7758 36418 7810 36430
rect 19742 36482 19794 36494
rect 21646 36482 21698 36494
rect 20178 36430 20190 36482
rect 20242 36430 20254 36482
rect 19742 36418 19794 36430
rect 21646 36418 21698 36430
rect 21870 36482 21922 36494
rect 21870 36418 21922 36430
rect 37662 36482 37714 36494
rect 37662 36418 37714 36430
rect 37102 36370 37154 36382
rect 7970 36318 7982 36370
rect 8034 36318 8046 36370
rect 8530 36318 8542 36370
rect 8594 36318 8606 36370
rect 37102 36306 37154 36318
rect 37774 36370 37826 36382
rect 37774 36306 37826 36318
rect 40686 36370 40738 36382
rect 40686 36306 40738 36318
rect 37214 36258 37266 36270
rect 20402 36206 20414 36258
rect 20466 36206 20478 36258
rect 37214 36194 37266 36206
rect 37438 36258 37490 36270
rect 37438 36194 37490 36206
rect 37998 36258 38050 36270
rect 37998 36194 38050 36206
rect 40798 36258 40850 36270
rect 40798 36194 40850 36206
rect 1344 36090 44576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 44576 36090
rect 1344 36004 44576 36038
rect 24546 35870 24558 35922
rect 24610 35870 24622 35922
rect 19854 35810 19906 35822
rect 19854 35746 19906 35758
rect 20078 35810 20130 35822
rect 37438 35810 37490 35822
rect 23650 35758 23662 35810
rect 23714 35758 23726 35810
rect 29698 35758 29710 35810
rect 29762 35758 29774 35810
rect 20078 35746 20130 35758
rect 37438 35746 37490 35758
rect 40014 35810 40066 35822
rect 40014 35746 40066 35758
rect 30942 35698 30994 35710
rect 37102 35698 37154 35710
rect 23538 35646 23550 35698
rect 23602 35646 23614 35698
rect 24658 35646 24670 35698
rect 24722 35646 24734 35698
rect 30482 35646 30494 35698
rect 30546 35646 30558 35698
rect 36754 35646 36766 35698
rect 36818 35646 36830 35698
rect 30942 35634 30994 35646
rect 37102 35634 37154 35646
rect 37550 35698 37602 35710
rect 37550 35634 37602 35646
rect 38110 35698 38162 35710
rect 38110 35634 38162 35646
rect 39454 35698 39506 35710
rect 39454 35634 39506 35646
rect 39790 35698 39842 35710
rect 39790 35634 39842 35646
rect 40462 35698 40514 35710
rect 40898 35646 40910 35698
rect 40962 35646 40974 35698
rect 40462 35634 40514 35646
rect 9886 35586 9938 35598
rect 37214 35586 37266 35598
rect 27570 35534 27582 35586
rect 27634 35534 27646 35586
rect 33842 35534 33854 35586
rect 33906 35534 33918 35586
rect 35970 35534 35982 35586
rect 36034 35534 36046 35586
rect 9886 35522 9938 35534
rect 37214 35522 37266 35534
rect 40238 35586 40290 35598
rect 41682 35534 41694 35586
rect 41746 35534 41758 35586
rect 43810 35534 43822 35586
rect 43874 35534 43886 35586
rect 40238 35522 40290 35534
rect 20190 35474 20242 35486
rect 20190 35410 20242 35422
rect 1344 35306 44576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 44576 35306
rect 1344 35220 44576 35254
rect 21422 35138 21474 35150
rect 21422 35074 21474 35086
rect 37102 35138 37154 35150
rect 37102 35074 37154 35086
rect 5742 35026 5794 35038
rect 5058 34974 5070 35026
rect 5122 34974 5134 35026
rect 5742 34962 5794 34974
rect 6974 35026 7026 35038
rect 11006 35026 11058 35038
rect 20638 35026 20690 35038
rect 8530 34974 8542 35026
rect 8594 34974 8606 35026
rect 13794 34974 13806 35026
rect 13858 34974 13870 35026
rect 27122 34974 27134 35026
rect 27186 34974 27198 35026
rect 33394 34974 33406 35026
rect 33458 34974 33470 35026
rect 6974 34962 7026 34974
rect 11006 34962 11058 34974
rect 20638 34962 20690 34974
rect 7310 34914 7362 34926
rect 9774 34914 9826 34926
rect 20190 34914 20242 34926
rect 2258 34862 2270 34914
rect 2322 34862 2334 34914
rect 7634 34862 7646 34914
rect 7698 34862 7710 34914
rect 8418 34862 8430 34914
rect 8482 34862 8494 34914
rect 9314 34862 9326 34914
rect 9378 34862 9390 34914
rect 9538 34862 9550 34914
rect 9602 34862 9614 34914
rect 16594 34862 16606 34914
rect 16658 34862 16670 34914
rect 7310 34850 7362 34862
rect 9774 34850 9826 34862
rect 20190 34850 20242 34862
rect 20414 34914 20466 34926
rect 20414 34850 20466 34862
rect 21310 34914 21362 34926
rect 24434 34862 24446 34914
rect 24498 34862 24510 34914
rect 25218 34862 25230 34914
rect 25282 34862 25294 34914
rect 26674 34862 26686 34914
rect 26738 34862 26750 34914
rect 27010 34862 27022 34914
rect 27074 34862 27086 34914
rect 30594 34862 30606 34914
rect 30658 34862 30670 34914
rect 21310 34850 21362 34862
rect 10110 34802 10162 34814
rect 20750 34802 20802 34814
rect 37102 34802 37154 34814
rect 2930 34750 2942 34802
rect 2994 34750 3006 34802
rect 15922 34750 15934 34802
rect 15986 34750 15998 34802
rect 28018 34750 28030 34802
rect 28082 34750 28094 34802
rect 31266 34750 31278 34802
rect 31330 34750 31342 34802
rect 10110 34738 10162 34750
rect 20750 34738 20802 34750
rect 37102 34738 37154 34750
rect 37214 34802 37266 34814
rect 37214 34738 37266 34750
rect 40686 34802 40738 34814
rect 40686 34738 40738 34750
rect 9998 34690 10050 34702
rect 9998 34626 10050 34638
rect 10670 34690 10722 34702
rect 10670 34626 10722 34638
rect 17166 34690 17218 34702
rect 17166 34626 17218 34638
rect 21422 34690 21474 34702
rect 33854 34690 33906 34702
rect 24210 34638 24222 34690
rect 24274 34638 24286 34690
rect 21422 34626 21474 34638
rect 33854 34626 33906 34638
rect 40350 34690 40402 34702
rect 40350 34626 40402 34638
rect 40574 34690 40626 34702
rect 40574 34626 40626 34638
rect 1344 34522 44576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 44576 34522
rect 1344 34436 44576 34470
rect 8542 34354 8594 34366
rect 8542 34290 8594 34302
rect 8766 34354 8818 34366
rect 8766 34290 8818 34302
rect 10894 34354 10946 34366
rect 10894 34290 10946 34302
rect 11678 34354 11730 34366
rect 11678 34290 11730 34302
rect 15598 34354 15650 34366
rect 15598 34290 15650 34302
rect 32062 34354 32114 34366
rect 32062 34290 32114 34302
rect 9998 34242 10050 34254
rect 23326 34242 23378 34254
rect 12002 34190 12014 34242
rect 12066 34190 12078 34242
rect 9998 34178 10050 34190
rect 23326 34178 23378 34190
rect 23438 34242 23490 34254
rect 23438 34178 23490 34190
rect 25230 34242 25282 34254
rect 25230 34178 25282 34190
rect 31838 34242 31890 34254
rect 31838 34178 31890 34190
rect 8878 34130 8930 34142
rect 10558 34130 10610 34142
rect 10210 34078 10222 34130
rect 10274 34078 10286 34130
rect 8878 34066 8930 34078
rect 10558 34066 10610 34078
rect 10670 34130 10722 34142
rect 10670 34066 10722 34078
rect 11006 34130 11058 34142
rect 11006 34066 11058 34078
rect 11342 34130 11394 34142
rect 11342 34066 11394 34078
rect 15374 34130 15426 34142
rect 15374 34066 15426 34078
rect 15710 34130 15762 34142
rect 15710 34066 15762 34078
rect 15934 34130 15986 34142
rect 15934 34066 15986 34078
rect 20638 34130 20690 34142
rect 22206 34130 22258 34142
rect 21074 34078 21086 34130
rect 21138 34078 21150 34130
rect 20638 34066 20690 34078
rect 22206 34066 22258 34078
rect 22766 34130 22818 34142
rect 22766 34066 22818 34078
rect 25342 34130 25394 34142
rect 30830 34130 30882 34142
rect 25778 34078 25790 34130
rect 25842 34078 25854 34130
rect 25342 34066 25394 34078
rect 30830 34066 30882 34078
rect 30942 34130 30994 34142
rect 30942 34066 30994 34078
rect 31166 34130 31218 34142
rect 31726 34130 31778 34142
rect 31378 34078 31390 34130
rect 31442 34078 31454 34130
rect 31166 34066 31218 34078
rect 31726 34066 31778 34078
rect 9662 34018 9714 34030
rect 9662 33954 9714 33966
rect 12462 34018 12514 34030
rect 12462 33954 12514 33966
rect 16382 34018 16434 34030
rect 16382 33954 16434 33966
rect 23886 34018 23938 34030
rect 23886 33954 23938 33966
rect 29710 34018 29762 34030
rect 29710 33954 29762 33966
rect 30158 34018 30210 34030
rect 32398 34018 32450 34030
rect 31266 33966 31278 34018
rect 31330 33966 31342 34018
rect 30158 33954 30210 33966
rect 32398 33954 32450 33966
rect 10334 33906 10386 33918
rect 10334 33842 10386 33854
rect 23102 33906 23154 33918
rect 23102 33842 23154 33854
rect 23662 33906 23714 33918
rect 23662 33842 23714 33854
rect 25566 33906 25618 33918
rect 25566 33842 25618 33854
rect 1344 33738 44576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 44576 33738
rect 1344 33652 44576 33686
rect 11902 33458 11954 33470
rect 6962 33406 6974 33458
rect 7026 33406 7038 33458
rect 11902 33394 11954 33406
rect 12798 33458 12850 33470
rect 34638 33458 34690 33470
rect 15362 33406 15374 33458
rect 15426 33406 15438 33458
rect 43810 33406 43822 33458
rect 43874 33406 43886 33458
rect 12798 33394 12850 33406
rect 34638 33394 34690 33406
rect 8206 33346 8258 33358
rect 8206 33282 8258 33294
rect 12350 33346 12402 33358
rect 40014 33346 40066 33358
rect 25890 33294 25902 33346
rect 25954 33294 25966 33346
rect 26562 33294 26574 33346
rect 26626 33294 26638 33346
rect 12350 33282 12402 33294
rect 40014 33282 40066 33294
rect 40350 33346 40402 33358
rect 40898 33294 40910 33346
rect 40962 33294 40974 33346
rect 40350 33282 40402 33294
rect 7422 33234 7474 33246
rect 7298 33182 7310 33234
rect 7362 33182 7374 33234
rect 7422 33170 7474 33182
rect 11790 33234 11842 33246
rect 11790 33170 11842 33182
rect 12126 33234 12178 33246
rect 12126 33170 12178 33182
rect 15038 33234 15090 33246
rect 15038 33170 15090 33182
rect 15486 33234 15538 33246
rect 40462 33234 40514 33246
rect 25554 33182 25566 33234
rect 25618 33182 25630 33234
rect 41682 33182 41694 33234
rect 41746 33182 41758 33234
rect 15486 33170 15538 33182
rect 40462 33170 40514 33182
rect 7534 33122 7586 33134
rect 7534 33058 7586 33070
rect 7758 33122 7810 33134
rect 7758 33058 7810 33070
rect 10670 33122 10722 33134
rect 10670 33058 10722 33070
rect 14702 33122 14754 33134
rect 14702 33058 14754 33070
rect 15262 33122 15314 33134
rect 15262 33058 15314 33070
rect 17054 33122 17106 33134
rect 35758 33122 35810 33134
rect 26450 33070 26462 33122
rect 26514 33070 26526 33122
rect 17054 33058 17106 33070
rect 35758 33058 35810 33070
rect 35982 33122 36034 33134
rect 40686 33122 40738 33134
rect 36306 33070 36318 33122
rect 36370 33070 36382 33122
rect 35982 33058 36034 33070
rect 40686 33058 40738 33070
rect 1344 32954 44576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 44576 32954
rect 1344 32868 44576 32902
rect 5630 32786 5682 32798
rect 5630 32722 5682 32734
rect 6638 32786 6690 32798
rect 6638 32722 6690 32734
rect 7870 32786 7922 32798
rect 7870 32722 7922 32734
rect 8542 32786 8594 32798
rect 8542 32722 8594 32734
rect 11790 32786 11842 32798
rect 11790 32722 11842 32734
rect 12126 32786 12178 32798
rect 13918 32786 13970 32798
rect 13010 32734 13022 32786
rect 13074 32734 13086 32786
rect 12126 32722 12178 32734
rect 13918 32722 13970 32734
rect 15486 32786 15538 32798
rect 15486 32722 15538 32734
rect 17614 32786 17666 32798
rect 17614 32722 17666 32734
rect 20302 32786 20354 32798
rect 20302 32722 20354 32734
rect 21758 32786 21810 32798
rect 21758 32722 21810 32734
rect 33742 32786 33794 32798
rect 33742 32722 33794 32734
rect 41694 32786 41746 32798
rect 41694 32722 41746 32734
rect 41806 32786 41858 32798
rect 41806 32722 41858 32734
rect 6862 32674 6914 32686
rect 6862 32610 6914 32622
rect 7758 32674 7810 32686
rect 7758 32610 7810 32622
rect 11902 32674 11954 32686
rect 15822 32674 15874 32686
rect 13570 32622 13582 32674
rect 13634 32622 13646 32674
rect 11902 32610 11954 32622
rect 15822 32610 15874 32622
rect 17838 32674 17890 32686
rect 17838 32610 17890 32622
rect 25790 32674 25842 32686
rect 40786 32622 40798 32674
rect 40850 32671 40862 32674
rect 41010 32671 41022 32674
rect 40850 32625 41022 32671
rect 40850 32622 40862 32625
rect 41010 32622 41022 32625
rect 41074 32622 41086 32674
rect 25790 32610 25842 32622
rect 12462 32562 12514 32574
rect 2258 32510 2270 32562
rect 2322 32510 2334 32562
rect 7074 32510 7086 32562
rect 7138 32510 7150 32562
rect 7298 32510 7310 32562
rect 7362 32510 7374 32562
rect 12462 32498 12514 32510
rect 12686 32562 12738 32574
rect 12686 32498 12738 32510
rect 16046 32562 16098 32574
rect 16046 32498 16098 32510
rect 16494 32562 16546 32574
rect 16494 32498 16546 32510
rect 17278 32562 17330 32574
rect 17278 32498 17330 32510
rect 22206 32562 22258 32574
rect 22206 32498 22258 32510
rect 22430 32562 22482 32574
rect 41134 32562 41186 32574
rect 34178 32510 34190 32562
rect 34242 32510 34254 32562
rect 34962 32510 34974 32562
rect 35026 32510 35038 32562
rect 41458 32510 41470 32562
rect 41522 32510 41534 32562
rect 22430 32498 22482 32510
rect 41134 32498 41186 32510
rect 15038 32450 15090 32462
rect 3042 32398 3054 32450
rect 3106 32398 3118 32450
rect 5170 32398 5182 32450
rect 5234 32398 5246 32450
rect 6962 32398 6974 32450
rect 7026 32398 7038 32450
rect 15038 32386 15090 32398
rect 19406 32450 19458 32462
rect 19406 32386 19458 32398
rect 22654 32450 22706 32462
rect 30494 32450 30546 32462
rect 25666 32398 25678 32450
rect 25730 32398 25742 32450
rect 22654 32386 22706 32398
rect 30494 32386 30546 32398
rect 34638 32450 34690 32462
rect 35746 32398 35758 32450
rect 35810 32398 35822 32450
rect 37874 32398 37886 32450
rect 37938 32398 37950 32450
rect 34638 32386 34690 32398
rect 16270 32338 16322 32350
rect 16270 32274 16322 32286
rect 16942 32338 16994 32350
rect 16942 32274 16994 32286
rect 17950 32338 18002 32350
rect 17950 32274 18002 32286
rect 19630 32338 19682 32350
rect 19630 32274 19682 32286
rect 19854 32338 19906 32350
rect 19854 32274 19906 32286
rect 26014 32338 26066 32350
rect 26014 32274 26066 32286
rect 1344 32170 44576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 44576 32170
rect 1344 32084 44576 32118
rect 25678 32002 25730 32014
rect 25678 31938 25730 31950
rect 41694 32002 41746 32014
rect 41694 31938 41746 31950
rect 6190 31890 6242 31902
rect 6190 31826 6242 31838
rect 8542 31890 8594 31902
rect 8542 31826 8594 31838
rect 12686 31890 12738 31902
rect 20078 31890 20130 31902
rect 20638 31890 20690 31902
rect 26350 31890 26402 31902
rect 18274 31838 18286 31890
rect 18338 31838 18350 31890
rect 20402 31838 20414 31890
rect 20466 31838 20478 31890
rect 24882 31838 24894 31890
rect 24946 31838 24958 31890
rect 12686 31826 12738 31838
rect 20078 31826 20130 31838
rect 20638 31826 20690 31838
rect 26350 31826 26402 31838
rect 8766 31778 8818 31790
rect 8766 31714 8818 31726
rect 8990 31778 9042 31790
rect 19854 31778 19906 31790
rect 15586 31726 15598 31778
rect 15650 31726 15662 31778
rect 8990 31714 9042 31726
rect 19854 31714 19906 31726
rect 25230 31778 25282 31790
rect 25230 31714 25282 31726
rect 25454 31778 25506 31790
rect 25454 31714 25506 31726
rect 26126 31778 26178 31790
rect 26126 31714 26178 31726
rect 26574 31778 26626 31790
rect 30370 31726 30382 31778
rect 30434 31726 30446 31778
rect 30706 31726 30718 31778
rect 30770 31726 30782 31778
rect 26574 31714 26626 31726
rect 6078 31666 6130 31678
rect 6078 31602 6130 31614
rect 20414 31666 20466 31678
rect 37214 31666 37266 31678
rect 34066 31614 34078 31666
rect 34130 31614 34142 31666
rect 20414 31602 20466 31614
rect 37214 31602 37266 31614
rect 41582 31666 41634 31678
rect 41582 31602 41634 31614
rect 9438 31554 9490 31566
rect 9438 31490 9490 31502
rect 11118 31554 11170 31566
rect 29822 31554 29874 31566
rect 11442 31502 11454 31554
rect 11506 31502 11518 31554
rect 11118 31490 11170 31502
rect 29822 31490 29874 31502
rect 29934 31554 29986 31566
rect 29934 31490 29986 31502
rect 30046 31554 30098 31566
rect 30046 31490 30098 31502
rect 36878 31554 36930 31566
rect 36878 31490 36930 31502
rect 37102 31554 37154 31566
rect 37102 31490 37154 31502
rect 41694 31554 41746 31566
rect 41694 31490 41746 31502
rect 1344 31386 44576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 44576 31386
rect 1344 31300 44576 31334
rect 6638 31218 6690 31230
rect 6638 31154 6690 31166
rect 10222 31218 10274 31230
rect 25902 31218 25954 31230
rect 18946 31166 18958 31218
rect 19010 31166 19022 31218
rect 10222 31154 10274 31166
rect 25902 31154 25954 31166
rect 26686 31218 26738 31230
rect 26686 31154 26738 31166
rect 34750 31218 34802 31230
rect 34750 31154 34802 31166
rect 35534 31218 35586 31230
rect 39330 31166 39342 31218
rect 39394 31166 39406 31218
rect 40338 31166 40350 31218
rect 40402 31166 40414 31218
rect 35534 31154 35586 31166
rect 29038 31106 29090 31118
rect 12002 31054 12014 31106
rect 12066 31054 12078 31106
rect 29038 31042 29090 31054
rect 35086 31106 35138 31118
rect 35086 31042 35138 31054
rect 10110 30994 10162 31006
rect 25566 30994 25618 31006
rect 15810 30942 15822 30994
rect 15874 30942 15886 30994
rect 19058 30942 19070 30994
rect 19122 30942 19134 30994
rect 19282 30942 19294 30994
rect 19346 30942 19358 30994
rect 19506 30942 19518 30994
rect 19570 30942 19582 30994
rect 10110 30930 10162 30942
rect 25566 30930 25618 30942
rect 26014 30994 26066 31006
rect 26014 30930 26066 30942
rect 26238 30994 26290 31006
rect 34862 30994 34914 31006
rect 26898 30942 26910 30994
rect 26962 30942 26974 30994
rect 29810 30942 29822 30994
rect 29874 30942 29886 30994
rect 30818 30942 30830 30994
rect 30882 30942 30894 30994
rect 26238 30930 26290 30942
rect 34862 30930 34914 30942
rect 35198 30994 35250 31006
rect 36094 30994 36146 31006
rect 35746 30942 35758 30994
rect 35810 30942 35822 30994
rect 35198 30930 35250 30942
rect 36094 30930 36146 30942
rect 39006 30994 39058 31006
rect 39006 30930 39058 30942
rect 40014 30994 40066 31006
rect 40014 30930 40066 30942
rect 9886 30882 9938 30894
rect 9886 30818 9938 30830
rect 16382 30882 16434 30894
rect 16382 30818 16434 30830
rect 20638 30882 20690 30894
rect 20638 30818 20690 30830
rect 26574 30882 26626 30894
rect 35870 30882 35922 30894
rect 31266 30830 31278 30882
rect 31330 30830 31342 30882
rect 26574 30818 26626 30830
rect 35870 30818 35922 30830
rect 38670 30882 38722 30894
rect 38670 30818 38722 30830
rect 10222 30770 10274 30782
rect 10222 30706 10274 30718
rect 1344 30602 44576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 44576 30602
rect 1344 30516 44576 30550
rect 19182 30434 19234 30446
rect 19182 30370 19234 30382
rect 19406 30434 19458 30446
rect 19406 30370 19458 30382
rect 19966 30322 20018 30334
rect 5842 30270 5854 30322
rect 5906 30270 5918 30322
rect 14914 30270 14926 30322
rect 14978 30270 14990 30322
rect 19966 30258 20018 30270
rect 6638 30210 6690 30222
rect 6066 30158 6078 30210
rect 6130 30158 6142 30210
rect 6638 30146 6690 30158
rect 6974 30210 7026 30222
rect 8878 30210 8930 30222
rect 13806 30210 13858 30222
rect 7410 30158 7422 30210
rect 7474 30158 7486 30210
rect 9202 30158 9214 30210
rect 9266 30158 9278 30210
rect 11218 30158 11230 30210
rect 11282 30158 11294 30210
rect 6974 30146 7026 30158
rect 8878 30146 8930 30158
rect 13806 30146 13858 30158
rect 14590 30210 14642 30222
rect 14590 30146 14642 30158
rect 16046 30210 16098 30222
rect 18734 30210 18786 30222
rect 16258 30158 16270 30210
rect 16322 30158 16334 30210
rect 16046 30146 16098 30158
rect 18734 30146 18786 30158
rect 19630 30210 19682 30222
rect 19630 30146 19682 30158
rect 19742 30210 19794 30222
rect 19742 30146 19794 30158
rect 25566 30210 25618 30222
rect 30382 30210 30434 30222
rect 26226 30158 26238 30210
rect 26290 30158 26302 30210
rect 27346 30158 27358 30210
rect 27410 30158 27422 30210
rect 25566 30146 25618 30158
rect 30382 30146 30434 30158
rect 30606 30210 30658 30222
rect 31726 30210 31778 30222
rect 31266 30158 31278 30210
rect 31330 30158 31342 30210
rect 30606 30146 30658 30158
rect 31726 30146 31778 30158
rect 36990 30210 37042 30222
rect 36990 30146 37042 30158
rect 7086 30098 7138 30110
rect 12126 30098 12178 30110
rect 11554 30046 11566 30098
rect 11618 30046 11630 30098
rect 7086 30034 7138 30046
rect 12126 30034 12178 30046
rect 15262 30098 15314 30110
rect 15262 30034 15314 30046
rect 15598 30098 15650 30110
rect 15598 30034 15650 30046
rect 25902 30098 25954 30110
rect 31950 30098 32002 30110
rect 27234 30046 27246 30098
rect 27298 30046 27310 30098
rect 25902 30034 25954 30046
rect 31950 30034 32002 30046
rect 32062 30098 32114 30110
rect 32062 30034 32114 30046
rect 37102 30098 37154 30110
rect 39554 30046 39566 30098
rect 39618 30046 39630 30098
rect 37102 30034 37154 30046
rect 11678 29986 11730 29998
rect 11678 29922 11730 29934
rect 13918 29986 13970 29998
rect 13918 29922 13970 29934
rect 15038 29986 15090 29998
rect 15038 29922 15090 29934
rect 15822 29986 15874 29998
rect 15822 29922 15874 29934
rect 15934 29986 15986 29998
rect 20414 29986 20466 29998
rect 18386 29934 18398 29986
rect 18450 29934 18462 29986
rect 15934 29922 15986 29934
rect 20414 29922 20466 29934
rect 25790 29986 25842 29998
rect 37326 29986 37378 29998
rect 26338 29934 26350 29986
rect 26402 29934 26414 29986
rect 25790 29922 25842 29934
rect 37326 29922 37378 29934
rect 38894 29986 38946 29998
rect 38894 29922 38946 29934
rect 39230 29986 39282 29998
rect 39230 29922 39282 29934
rect 1344 29818 44576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 44576 29818
rect 1344 29732 44576 29766
rect 5182 29650 5234 29662
rect 5182 29586 5234 29598
rect 9998 29650 10050 29662
rect 9998 29586 10050 29598
rect 14702 29650 14754 29662
rect 32386 29598 32398 29650
rect 32450 29598 32462 29650
rect 14702 29586 14754 29598
rect 10446 29538 10498 29550
rect 10446 29474 10498 29486
rect 11118 29538 11170 29550
rect 11118 29474 11170 29486
rect 14254 29538 14306 29550
rect 14254 29474 14306 29486
rect 14590 29538 14642 29550
rect 26014 29538 26066 29550
rect 33630 29538 33682 29550
rect 16258 29486 16270 29538
rect 16322 29486 16334 29538
rect 25554 29486 25566 29538
rect 25618 29486 25630 29538
rect 31714 29486 31726 29538
rect 31778 29486 31790 29538
rect 14590 29474 14642 29486
rect 26014 29474 26066 29486
rect 33630 29474 33682 29486
rect 5966 29426 6018 29438
rect 10222 29426 10274 29438
rect 1810 29374 1822 29426
rect 1874 29374 1886 29426
rect 9762 29374 9774 29426
rect 9826 29374 9838 29426
rect 5966 29362 6018 29374
rect 10222 29362 10274 29374
rect 11230 29426 11282 29438
rect 11230 29362 11282 29374
rect 11678 29426 11730 29438
rect 16494 29426 16546 29438
rect 15250 29374 15262 29426
rect 15314 29374 15326 29426
rect 15922 29374 15934 29426
rect 15986 29374 15998 29426
rect 11678 29362 11730 29374
rect 16494 29362 16546 29374
rect 25230 29426 25282 29438
rect 26910 29426 26962 29438
rect 26450 29374 26462 29426
rect 26514 29374 26526 29426
rect 25230 29362 25282 29374
rect 26910 29362 26962 29374
rect 31054 29426 31106 29438
rect 32062 29426 32114 29438
rect 31490 29374 31502 29426
rect 31554 29374 31566 29426
rect 31054 29362 31106 29374
rect 32062 29362 32114 29374
rect 33294 29426 33346 29438
rect 40350 29426 40402 29438
rect 33954 29374 33966 29426
rect 34018 29374 34030 29426
rect 40898 29374 40910 29426
rect 40962 29374 40974 29426
rect 33294 29362 33346 29374
rect 40350 29362 40402 29374
rect 24670 29314 24722 29326
rect 2594 29262 2606 29314
rect 2658 29262 2670 29314
rect 4722 29262 4734 29314
rect 4786 29262 4798 29314
rect 6402 29262 6414 29314
rect 6466 29262 6478 29314
rect 9986 29262 9998 29314
rect 10050 29262 10062 29314
rect 38546 29262 38558 29314
rect 38610 29262 38622 29314
rect 41682 29262 41694 29314
rect 41746 29262 41758 29314
rect 43810 29262 43822 29314
rect 43874 29262 43886 29314
rect 24670 29250 24722 29262
rect 11118 29202 11170 29214
rect 15698 29150 15710 29202
rect 15762 29150 15774 29202
rect 11118 29138 11170 29150
rect 1344 29034 44576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 44576 29034
rect 1344 28948 44576 28982
rect 6750 28866 6802 28878
rect 6750 28802 6802 28814
rect 9438 28866 9490 28878
rect 9438 28802 9490 28814
rect 15486 28866 15538 28878
rect 15486 28802 15538 28814
rect 16606 28866 16658 28878
rect 16606 28802 16658 28814
rect 42478 28866 42530 28878
rect 42478 28802 42530 28814
rect 6638 28754 6690 28766
rect 6638 28690 6690 28702
rect 9326 28754 9378 28766
rect 16718 28754 16770 28766
rect 10322 28702 10334 28754
rect 10386 28702 10398 28754
rect 9326 28690 9378 28702
rect 16718 28690 16770 28702
rect 17166 28754 17218 28766
rect 17166 28690 17218 28702
rect 19406 28754 19458 28766
rect 19406 28690 19458 28702
rect 33070 28754 33122 28766
rect 33070 28690 33122 28702
rect 33630 28754 33682 28766
rect 33630 28690 33682 28702
rect 41918 28754 41970 28766
rect 41918 28690 41970 28702
rect 10782 28642 10834 28654
rect 10098 28590 10110 28642
rect 10162 28590 10174 28642
rect 10782 28578 10834 28590
rect 15262 28642 15314 28654
rect 37326 28642 37378 28654
rect 15474 28590 15486 28642
rect 15538 28590 15550 28642
rect 15262 28578 15314 28590
rect 37326 28578 37378 28590
rect 37550 28642 37602 28654
rect 37550 28578 37602 28590
rect 37774 28642 37826 28654
rect 37774 28578 37826 28590
rect 41470 28642 41522 28654
rect 41470 28578 41522 28590
rect 42142 28642 42194 28654
rect 42142 28578 42194 28590
rect 15822 28530 15874 28542
rect 15822 28466 15874 28478
rect 16270 28530 16322 28542
rect 16270 28466 16322 28478
rect 36990 28530 37042 28542
rect 36990 28466 37042 28478
rect 38110 28530 38162 28542
rect 38110 28466 38162 28478
rect 41694 28530 41746 28542
rect 41694 28466 41746 28478
rect 42366 28530 42418 28542
rect 42366 28466 42418 28478
rect 42478 28530 42530 28542
rect 42478 28466 42530 28478
rect 16158 28418 16210 28430
rect 16158 28354 16210 28366
rect 37102 28418 37154 28430
rect 37102 28354 37154 28366
rect 37998 28418 38050 28430
rect 37998 28354 38050 28366
rect 1344 28250 44576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 44576 28250
rect 1344 28164 44576 28198
rect 15822 28082 15874 28094
rect 15822 28018 15874 28030
rect 16046 28082 16098 28094
rect 16046 28018 16098 28030
rect 38222 28082 38274 28094
rect 38994 28030 39006 28082
rect 39058 28030 39070 28082
rect 38222 28018 38274 28030
rect 13682 27918 13694 27970
rect 13746 27918 13758 27970
rect 25218 27918 25230 27970
rect 25282 27918 25294 27970
rect 36978 27918 36990 27970
rect 37042 27918 37054 27970
rect 15710 27858 15762 27870
rect 13570 27806 13582 27858
rect 13634 27806 13646 27858
rect 14018 27806 14030 27858
rect 14082 27806 14094 27858
rect 14914 27806 14926 27858
rect 14978 27806 14990 27858
rect 15710 27794 15762 27806
rect 16158 27858 16210 27870
rect 16158 27794 16210 27806
rect 18734 27858 18786 27870
rect 18734 27794 18786 27806
rect 19070 27858 19122 27870
rect 19070 27794 19122 27806
rect 19294 27858 19346 27870
rect 26014 27858 26066 27870
rect 39342 27858 39394 27870
rect 19730 27806 19742 27858
rect 19794 27806 19806 27858
rect 25442 27806 25454 27858
rect 25506 27806 25518 27858
rect 37762 27806 37774 27858
rect 37826 27806 37838 27858
rect 19294 27794 19346 27806
rect 26014 27794 26066 27806
rect 39342 27794 39394 27806
rect 13246 27746 13298 27758
rect 13246 27682 13298 27694
rect 15934 27746 15986 27758
rect 15934 27682 15986 27694
rect 18958 27746 19010 27758
rect 38670 27746 38722 27758
rect 20514 27694 20526 27746
rect 20578 27694 20590 27746
rect 22642 27694 22654 27746
rect 22706 27694 22718 27746
rect 34850 27694 34862 27746
rect 34914 27694 34926 27746
rect 18958 27682 19010 27694
rect 38670 27682 38722 27694
rect 15038 27634 15090 27646
rect 15038 27570 15090 27582
rect 1344 27466 44576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 44576 27466
rect 1344 27380 44576 27414
rect 30382 27298 30434 27310
rect 30382 27234 30434 27246
rect 30718 27298 30770 27310
rect 30718 27234 30770 27246
rect 15374 27186 15426 27198
rect 13794 27134 13806 27186
rect 13858 27134 13870 27186
rect 15374 27122 15426 27134
rect 19742 27186 19794 27198
rect 19742 27122 19794 27134
rect 21310 27186 21362 27198
rect 31266 27134 31278 27186
rect 31330 27134 31342 27186
rect 21310 27122 21362 27134
rect 12910 27074 12962 27086
rect 12910 27010 12962 27022
rect 13918 27074 13970 27086
rect 21422 27074 21474 27086
rect 35758 27074 35810 27086
rect 14354 27022 14366 27074
rect 14418 27022 14430 27074
rect 21746 27022 21758 27074
rect 21810 27022 21822 27074
rect 31826 27022 31838 27074
rect 31890 27022 31902 27074
rect 13918 27010 13970 27022
rect 21422 27010 21474 27022
rect 35758 27010 35810 27022
rect 13806 26962 13858 26974
rect 13806 26898 13858 26910
rect 25566 26962 25618 26974
rect 30046 26962 30098 26974
rect 25890 26910 25902 26962
rect 25954 26910 25966 26962
rect 25566 26898 25618 26910
rect 30046 26898 30098 26910
rect 30942 26962 30994 26974
rect 31714 26910 31726 26962
rect 31778 26910 31790 26962
rect 36082 26910 36094 26962
rect 36146 26910 36158 26962
rect 30942 26898 30994 26910
rect 7310 26850 7362 26862
rect 7310 26786 7362 26798
rect 12574 26850 12626 26862
rect 12574 26786 12626 26798
rect 14142 26850 14194 26862
rect 14142 26786 14194 26798
rect 1344 26682 44576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 44576 26682
rect 1344 26596 44576 26630
rect 5182 26514 5234 26526
rect 5182 26450 5234 26462
rect 7086 26514 7138 26526
rect 7086 26450 7138 26462
rect 11006 26514 11058 26526
rect 11006 26450 11058 26462
rect 11790 26514 11842 26526
rect 11790 26450 11842 26462
rect 12126 26514 12178 26526
rect 12126 26450 12178 26462
rect 12350 26514 12402 26526
rect 12350 26450 12402 26462
rect 15374 26514 15426 26526
rect 15374 26450 15426 26462
rect 17390 26514 17442 26526
rect 17390 26450 17442 26462
rect 23214 26514 23266 26526
rect 35634 26462 35646 26514
rect 35698 26462 35710 26514
rect 23214 26450 23266 26462
rect 6974 26402 7026 26414
rect 6974 26338 7026 26350
rect 11230 26402 11282 26414
rect 11230 26338 11282 26350
rect 12014 26402 12066 26414
rect 16830 26402 16882 26414
rect 12674 26350 12686 26402
rect 12738 26350 12750 26402
rect 12014 26338 12066 26350
rect 16830 26338 16882 26350
rect 17950 26402 18002 26414
rect 17950 26338 18002 26350
rect 18734 26402 18786 26414
rect 18734 26338 18786 26350
rect 19630 26402 19682 26414
rect 31602 26350 31614 26402
rect 31666 26350 31678 26402
rect 19630 26338 19682 26350
rect 10670 26290 10722 26302
rect 15486 26290 15538 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 6514 26238 6526 26290
rect 6578 26238 6590 26290
rect 6738 26238 6750 26290
rect 6802 26238 6814 26290
rect 7746 26238 7758 26290
rect 7810 26238 7822 26290
rect 11554 26238 11566 26290
rect 11618 26238 11630 26290
rect 10670 26226 10722 26238
rect 15486 26226 15538 26238
rect 16270 26290 16322 26302
rect 19294 26290 19346 26302
rect 30046 26290 30098 26302
rect 16594 26238 16606 26290
rect 16658 26238 16670 26290
rect 18946 26238 18958 26290
rect 19010 26238 19022 26290
rect 27010 26238 27022 26290
rect 27074 26238 27086 26290
rect 16270 26226 16322 26238
rect 19294 26226 19346 26238
rect 30046 26226 30098 26238
rect 30494 26290 30546 26302
rect 30494 26226 30546 26238
rect 30718 26290 30770 26302
rect 30718 26226 30770 26238
rect 31278 26290 31330 26302
rect 31278 26226 31330 26238
rect 31950 26290 32002 26302
rect 35410 26238 35422 26290
rect 35474 26238 35486 26290
rect 31950 26226 32002 26238
rect 7310 26178 7362 26190
rect 10894 26178 10946 26190
rect 2594 26126 2606 26178
rect 2658 26126 2670 26178
rect 4722 26126 4734 26178
rect 4786 26126 4798 26178
rect 8194 26126 8206 26178
rect 8258 26126 8270 26178
rect 7310 26114 7362 26126
rect 10894 26114 10946 26126
rect 13134 26178 13186 26190
rect 13134 26114 13186 26126
rect 16494 26178 16546 26190
rect 16494 26114 16546 26126
rect 17502 26178 17554 26190
rect 17502 26114 17554 26126
rect 19070 26178 19122 26190
rect 19070 26114 19122 26126
rect 23774 26178 23826 26190
rect 30270 26178 30322 26190
rect 27682 26126 27694 26178
rect 27746 26126 27758 26178
rect 29810 26126 29822 26178
rect 29874 26126 29886 26178
rect 32386 26126 32398 26178
rect 32450 26126 32462 26178
rect 23774 26114 23826 26126
rect 30270 26114 30322 26126
rect 1344 25898 44576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 44576 25898
rect 1344 25812 44576 25846
rect 4062 25730 4114 25742
rect 4062 25666 4114 25678
rect 7422 25730 7474 25742
rect 11330 25678 11342 25730
rect 11394 25727 11406 25730
rect 11554 25727 11566 25730
rect 11394 25681 11566 25727
rect 11394 25678 11406 25681
rect 11554 25678 11566 25681
rect 11618 25678 11630 25730
rect 7422 25666 7474 25678
rect 4398 25618 4450 25630
rect 40238 25618 40290 25630
rect 5842 25566 5854 25618
rect 5906 25566 5918 25618
rect 37874 25566 37886 25618
rect 37938 25566 37950 25618
rect 44034 25566 44046 25618
rect 44098 25566 44110 25618
rect 4398 25554 4450 25566
rect 40238 25554 40290 25566
rect 6750 25506 6802 25518
rect 40574 25506 40626 25518
rect 7074 25454 7086 25506
rect 7138 25454 7150 25506
rect 30818 25454 30830 25506
rect 30882 25454 30894 25506
rect 37426 25454 37438 25506
rect 37490 25454 37502 25506
rect 41122 25454 41134 25506
rect 41186 25454 41198 25506
rect 6750 25442 6802 25454
rect 40574 25442 40626 25454
rect 5854 25394 5906 25406
rect 5854 25330 5906 25342
rect 6302 25394 6354 25406
rect 29598 25394 29650 25406
rect 36990 25394 37042 25406
rect 17266 25342 17278 25394
rect 17330 25342 17342 25394
rect 29922 25342 29934 25394
rect 29986 25342 29998 25394
rect 30706 25342 30718 25394
rect 30770 25342 30782 25394
rect 6302 25330 6354 25342
rect 29598 25330 29650 25342
rect 36990 25330 37042 25342
rect 40686 25394 40738 25406
rect 41906 25342 41918 25394
rect 41970 25342 41982 25394
rect 40686 25330 40738 25342
rect 4174 25282 4226 25294
rect 4174 25218 4226 25230
rect 4846 25282 4898 25294
rect 4846 25218 4898 25230
rect 5742 25282 5794 25294
rect 5742 25218 5794 25230
rect 6078 25282 6130 25294
rect 6078 25218 6130 25230
rect 7310 25282 7362 25294
rect 7310 25218 7362 25230
rect 7758 25282 7810 25294
rect 7758 25218 7810 25230
rect 11454 25282 11506 25294
rect 11454 25218 11506 25230
rect 17614 25282 17666 25294
rect 17614 25218 17666 25230
rect 31278 25282 31330 25294
rect 31278 25218 31330 25230
rect 40910 25282 40962 25294
rect 40910 25218 40962 25230
rect 1344 25114 44576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 44576 25114
rect 1344 25028 44576 25062
rect 8654 24946 8706 24958
rect 8654 24882 8706 24894
rect 25230 24946 25282 24958
rect 25230 24882 25282 24894
rect 29262 24946 29314 24958
rect 29262 24882 29314 24894
rect 35646 24946 35698 24958
rect 35646 24882 35698 24894
rect 36542 24946 36594 24958
rect 36542 24882 36594 24894
rect 41806 24946 41858 24958
rect 41806 24882 41858 24894
rect 5518 24834 5570 24846
rect 5518 24770 5570 24782
rect 6638 24834 6690 24846
rect 6638 24770 6690 24782
rect 8878 24834 8930 24846
rect 8878 24770 8930 24782
rect 28702 24834 28754 24846
rect 28702 24770 28754 24782
rect 29934 24834 29986 24846
rect 35870 24834 35922 24846
rect 31378 24782 31390 24834
rect 31442 24782 31454 24834
rect 29934 24770 29986 24782
rect 35870 24770 35922 24782
rect 35982 24834 36034 24846
rect 35982 24770 36034 24782
rect 36654 24834 36706 24846
rect 36654 24770 36706 24782
rect 39230 24834 39282 24846
rect 40002 24782 40014 24834
rect 40066 24782 40078 24834
rect 39230 24770 39282 24782
rect 6078 24722 6130 24734
rect 6078 24658 6130 24670
rect 6190 24722 6242 24734
rect 6190 24658 6242 24670
rect 6414 24722 6466 24734
rect 6414 24658 6466 24670
rect 8990 24722 9042 24734
rect 28590 24722 28642 24734
rect 15586 24670 15598 24722
rect 15650 24670 15662 24722
rect 16034 24670 16046 24722
rect 16098 24670 16110 24722
rect 8990 24658 9042 24670
rect 28590 24658 28642 24670
rect 28926 24722 28978 24734
rect 28926 24658 28978 24670
rect 29150 24722 29202 24734
rect 36206 24722 36258 24734
rect 29474 24670 29486 24722
rect 29538 24670 29550 24722
rect 31602 24670 31614 24722
rect 31666 24670 31678 24722
rect 29150 24658 29202 24670
rect 36206 24658 36258 24670
rect 39118 24722 39170 24734
rect 41470 24722 41522 24734
rect 39778 24670 39790 24722
rect 39842 24670 39854 24722
rect 39118 24658 39170 24670
rect 41470 24658 41522 24670
rect 41918 24722 41970 24734
rect 41918 24658 41970 24670
rect 42030 24722 42082 24734
rect 42030 24658 42082 24670
rect 6302 24610 6354 24622
rect 6302 24546 6354 24558
rect 16270 24610 16322 24622
rect 16270 24546 16322 24558
rect 25790 24610 25842 24622
rect 25790 24546 25842 24558
rect 38782 24610 38834 24622
rect 38782 24546 38834 24558
rect 5630 24498 5682 24510
rect 5630 24434 5682 24446
rect 36542 24498 36594 24510
rect 36542 24434 36594 24446
rect 39230 24498 39282 24510
rect 39230 24434 39282 24446
rect 1344 24330 44576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 44576 24330
rect 1344 24244 44576 24278
rect 3726 24162 3778 24174
rect 3726 24098 3778 24110
rect 4062 24162 4114 24174
rect 4062 24098 4114 24110
rect 13806 24162 13858 24174
rect 13806 24098 13858 24110
rect 9214 24050 9266 24062
rect 9214 23986 9266 23998
rect 11454 24050 11506 24062
rect 11454 23986 11506 23998
rect 14254 24050 14306 24062
rect 38670 24050 38722 24062
rect 16258 23998 16270 24050
rect 16322 23998 16334 24050
rect 21410 23998 21422 24050
rect 21474 23998 21486 24050
rect 41794 23998 41806 24050
rect 41858 23998 41870 24050
rect 14254 23986 14306 23998
rect 38670 23986 38722 23998
rect 9438 23938 9490 23950
rect 16718 23938 16770 23950
rect 9090 23886 9102 23938
rect 9154 23886 9166 23938
rect 10770 23886 10782 23938
rect 10834 23886 10846 23938
rect 11218 23886 11230 23938
rect 11282 23886 11294 23938
rect 9438 23874 9490 23886
rect 16718 23874 16770 23886
rect 16942 23938 16994 23950
rect 16942 23874 16994 23886
rect 17166 23938 17218 23950
rect 17166 23874 17218 23886
rect 17278 23938 17330 23950
rect 17278 23874 17330 23886
rect 20750 23938 20802 23950
rect 42030 23938 42082 23950
rect 24210 23886 24222 23938
rect 24274 23886 24286 23938
rect 38882 23886 38894 23938
rect 38946 23886 38958 23938
rect 20750 23874 20802 23886
rect 42030 23874 42082 23886
rect 42366 23938 42418 23950
rect 42366 23874 42418 23886
rect 13582 23826 13634 23838
rect 20402 23774 20414 23826
rect 20466 23774 20478 23826
rect 23538 23774 23550 23826
rect 23602 23774 23614 23826
rect 39666 23774 39678 23826
rect 39730 23774 39742 23826
rect 13582 23762 13634 23774
rect 3838 23714 3890 23726
rect 3838 23650 3890 23662
rect 8878 23714 8930 23726
rect 8878 23650 8930 23662
rect 13694 23714 13746 23726
rect 13694 23650 13746 23662
rect 17726 23714 17778 23726
rect 17726 23650 17778 23662
rect 24782 23714 24834 23726
rect 24782 23650 24834 23662
rect 42254 23714 42306 23726
rect 42254 23650 42306 23662
rect 1344 23546 44576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 44576 23546
rect 1344 23460 44576 23494
rect 11230 23378 11282 23390
rect 8194 23326 8206 23378
rect 8258 23326 8270 23378
rect 11230 23314 11282 23326
rect 11454 23378 11506 23390
rect 12350 23378 12402 23390
rect 12002 23326 12014 23378
rect 12066 23326 12078 23378
rect 11454 23314 11506 23326
rect 12350 23314 12402 23326
rect 17390 23378 17442 23390
rect 17390 23314 17442 23326
rect 39566 23378 39618 23390
rect 39566 23314 39618 23326
rect 6302 23266 6354 23278
rect 6302 23202 6354 23214
rect 17502 23266 17554 23278
rect 17502 23202 17554 23214
rect 35310 23266 35362 23278
rect 35310 23202 35362 23214
rect 36094 23266 36146 23278
rect 36094 23202 36146 23214
rect 36206 23266 36258 23278
rect 36206 23202 36258 23214
rect 39902 23266 39954 23278
rect 39902 23202 39954 23214
rect 6190 23154 6242 23166
rect 11118 23154 11170 23166
rect 5842 23102 5854 23154
rect 5906 23102 5918 23154
rect 7970 23102 7982 23154
rect 8034 23102 8046 23154
rect 10210 23102 10222 23154
rect 10274 23102 10286 23154
rect 6190 23090 6242 23102
rect 11118 23090 11170 23102
rect 11566 23154 11618 23166
rect 28478 23154 28530 23166
rect 36430 23154 36482 23166
rect 17714 23102 17726 23154
rect 17778 23102 17790 23154
rect 17938 23102 17950 23154
rect 18002 23102 18014 23154
rect 19170 23102 19182 23154
rect 19234 23102 19246 23154
rect 28242 23102 28254 23154
rect 28306 23102 28318 23154
rect 31378 23102 31390 23154
rect 31442 23102 31454 23154
rect 35634 23102 35646 23154
rect 35698 23102 35710 23154
rect 11566 23090 11618 23102
rect 28478 23090 28530 23102
rect 36430 23090 36482 23102
rect 39230 23154 39282 23166
rect 39230 23090 39282 23102
rect 39678 23154 39730 23166
rect 39678 23090 39730 23102
rect 11342 23042 11394 23054
rect 27582 23042 27634 23054
rect 9874 22990 9886 23042
rect 9938 22990 9950 23042
rect 18834 22990 18846 23042
rect 18898 22990 18910 23042
rect 11342 22978 11394 22990
rect 27582 22978 27634 22990
rect 30830 23042 30882 23054
rect 32286 23042 32338 23054
rect 31714 22990 31726 23042
rect 31778 22990 31790 23042
rect 36082 22990 36094 23042
rect 36146 22990 36158 23042
rect 30830 22978 30882 22990
rect 32286 22978 32338 22990
rect 10210 22878 10222 22930
rect 10274 22878 10286 22930
rect 19282 22878 19294 22930
rect 19346 22878 19358 22930
rect 1344 22762 44576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 44576 22762
rect 1344 22676 44576 22710
rect 21758 22594 21810 22606
rect 21758 22530 21810 22542
rect 4174 22482 4226 22494
rect 21422 22482 21474 22494
rect 5730 22430 5742 22482
rect 5794 22430 5806 22482
rect 8418 22430 8430 22482
rect 8482 22430 8494 22482
rect 19842 22430 19854 22482
rect 19906 22430 19918 22482
rect 26674 22430 26686 22482
rect 26738 22430 26750 22482
rect 36418 22430 36430 22482
rect 36482 22430 36494 22482
rect 4174 22418 4226 22430
rect 21422 22418 21474 22430
rect 6078 22370 6130 22382
rect 17950 22370 18002 22382
rect 3826 22318 3838 22370
rect 3890 22318 3902 22370
rect 5618 22318 5630 22370
rect 5682 22318 5694 22370
rect 9762 22318 9774 22370
rect 9826 22318 9838 22370
rect 11218 22318 11230 22370
rect 11282 22318 11294 22370
rect 6078 22306 6130 22318
rect 17950 22306 18002 22318
rect 18286 22370 18338 22382
rect 18286 22306 18338 22318
rect 18622 22370 18674 22382
rect 19742 22370 19794 22382
rect 37102 22370 37154 22382
rect 19282 22318 19294 22370
rect 19346 22318 19358 22370
rect 22194 22318 22206 22370
rect 22258 22318 22270 22370
rect 33618 22318 33630 22370
rect 33682 22318 33694 22370
rect 18622 22306 18674 22318
rect 19742 22306 19794 22318
rect 37102 22306 37154 22318
rect 6302 22258 6354 22270
rect 18398 22258 18450 22270
rect 9874 22206 9886 22258
rect 9938 22206 9950 22258
rect 10882 22206 10894 22258
rect 10946 22206 10958 22258
rect 34290 22206 34302 22258
rect 34354 22206 34366 22258
rect 6302 22194 6354 22206
rect 18398 22194 18450 22206
rect 4062 22146 4114 22158
rect 4062 22082 4114 22094
rect 5854 22146 5906 22158
rect 19518 22146 19570 22158
rect 17602 22094 17614 22146
rect 17666 22094 17678 22146
rect 5854 22082 5906 22094
rect 19518 22082 19570 22094
rect 19854 22146 19906 22158
rect 19854 22082 19906 22094
rect 21646 22146 21698 22158
rect 21646 22082 21698 22094
rect 1344 21978 44576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 44576 21978
rect 1344 21892 44576 21926
rect 15486 21810 15538 21822
rect 4834 21758 4846 21810
rect 4898 21758 4910 21810
rect 15486 21746 15538 21758
rect 21982 21810 22034 21822
rect 21982 21746 22034 21758
rect 35310 21810 35362 21822
rect 35310 21746 35362 21758
rect 15934 21698 15986 21710
rect 2594 21646 2606 21698
rect 2658 21646 2670 21698
rect 15934 21634 15986 21646
rect 35422 21698 35474 21710
rect 35422 21634 35474 21646
rect 15710 21586 15762 21598
rect 1922 21534 1934 21586
rect 1986 21534 1998 21586
rect 15250 21534 15262 21586
rect 15314 21534 15326 21586
rect 25442 21534 25454 21586
rect 25506 21534 25518 21586
rect 29586 21534 29598 21586
rect 29650 21534 29662 21586
rect 15710 21522 15762 21534
rect 5518 21474 5570 21486
rect 5518 21410 5570 21422
rect 15598 21474 15650 21486
rect 28702 21474 28754 21486
rect 33182 21474 33234 21486
rect 26114 21422 26126 21474
rect 26178 21422 26190 21474
rect 28242 21422 28254 21474
rect 28306 21422 28318 21474
rect 30258 21422 30270 21474
rect 30322 21422 30334 21474
rect 32386 21422 32398 21474
rect 32450 21422 32462 21474
rect 15598 21410 15650 21422
rect 28702 21410 28754 21422
rect 33182 21410 33234 21422
rect 1344 21194 44576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 44576 21194
rect 1344 21108 44576 21142
rect 10894 21026 10946 21038
rect 10894 20962 10946 20974
rect 14702 21026 14754 21038
rect 14702 20962 14754 20974
rect 27022 21026 27074 21038
rect 27022 20962 27074 20974
rect 27358 21026 27410 21038
rect 27358 20962 27410 20974
rect 30494 21026 30546 21038
rect 30494 20962 30546 20974
rect 41806 21026 41858 21038
rect 41806 20962 41858 20974
rect 19630 20914 19682 20926
rect 10546 20862 10558 20914
rect 10610 20862 10622 20914
rect 14354 20862 14366 20914
rect 14418 20862 14430 20914
rect 19630 20850 19682 20862
rect 23774 20914 23826 20926
rect 23774 20850 23826 20862
rect 24110 20914 24162 20926
rect 36318 20914 36370 20926
rect 30258 20862 30270 20914
rect 30322 20862 30334 20914
rect 36194 20862 36206 20914
rect 36258 20862 36270 20914
rect 24110 20850 24162 20862
rect 36318 20850 36370 20862
rect 18846 20802 18898 20814
rect 18846 20738 18898 20750
rect 26686 20802 26738 20814
rect 29822 20802 29874 20814
rect 41918 20802 41970 20814
rect 27010 20750 27022 20802
rect 27074 20750 27086 20802
rect 30146 20750 30158 20802
rect 30210 20750 30222 20802
rect 32386 20750 32398 20802
rect 32450 20750 32462 20802
rect 35970 20750 35982 20802
rect 36034 20750 36046 20802
rect 26686 20738 26738 20750
rect 29822 20738 29874 20750
rect 41918 20738 41970 20750
rect 19170 20638 19182 20690
rect 19234 20638 19246 20690
rect 24434 20638 24446 20690
rect 24498 20638 24510 20690
rect 32162 20638 32174 20690
rect 32226 20638 32238 20690
rect 10670 20578 10722 20590
rect 10670 20514 10722 20526
rect 13582 20578 13634 20590
rect 13582 20514 13634 20526
rect 14478 20578 14530 20590
rect 14478 20514 14530 20526
rect 24782 20578 24834 20590
rect 24782 20514 24834 20526
rect 25118 20578 25170 20590
rect 31950 20578 32002 20590
rect 25442 20526 25454 20578
rect 25506 20526 25518 20578
rect 25118 20514 25170 20526
rect 31950 20514 32002 20526
rect 41806 20578 41858 20590
rect 41806 20514 41858 20526
rect 1344 20410 44576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 44576 20410
rect 1344 20324 44576 20358
rect 19630 20242 19682 20254
rect 19630 20178 19682 20190
rect 23998 20242 24050 20254
rect 23998 20178 24050 20190
rect 24558 20242 24610 20254
rect 24558 20178 24610 20190
rect 18846 20130 18898 20142
rect 10546 20078 10558 20130
rect 10610 20078 10622 20130
rect 14354 20078 14366 20130
rect 14418 20078 14430 20130
rect 18846 20066 18898 20078
rect 19182 20130 19234 20142
rect 39118 20130 39170 20142
rect 23650 20078 23662 20130
rect 23714 20078 23726 20130
rect 19182 20066 19234 20078
rect 39118 20066 39170 20078
rect 39454 20130 39506 20142
rect 39778 20078 39790 20130
rect 39842 20078 39854 20130
rect 39454 20066 39506 20078
rect 17614 20018 17666 20030
rect 9874 19966 9886 20018
rect 9938 19966 9950 20018
rect 13682 19966 13694 20018
rect 13746 19966 13758 20018
rect 17614 19954 17666 19966
rect 17950 20018 18002 20030
rect 19406 20018 19458 20030
rect 18274 19966 18286 20018
rect 18338 19966 18350 20018
rect 17950 19954 18002 19966
rect 19406 19954 19458 19966
rect 19742 20018 19794 20030
rect 20962 19966 20974 20018
rect 21026 19966 21038 20018
rect 41122 19966 41134 20018
rect 41186 19966 41198 20018
rect 19742 19954 19794 19966
rect 12686 19906 12738 19918
rect 20638 19906 20690 19918
rect 16482 19854 16494 19906
rect 16546 19854 16558 19906
rect 19618 19854 19630 19906
rect 19682 19854 19694 19906
rect 12686 19842 12738 19854
rect 20638 19842 20690 19854
rect 40350 19906 40402 19918
rect 41906 19854 41918 19906
rect 41970 19854 41982 19906
rect 44034 19854 44046 19906
rect 44098 19854 44110 19906
rect 40350 19842 40402 19854
rect 20974 19794 21026 19806
rect 20974 19730 21026 19742
rect 1344 19626 44576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 44576 19626
rect 1344 19540 44576 19574
rect 6414 19346 6466 19358
rect 6066 19294 6078 19346
rect 6130 19294 6142 19346
rect 6414 19282 6466 19294
rect 18958 19346 19010 19358
rect 18958 19282 19010 19294
rect 41806 19346 41858 19358
rect 41806 19282 41858 19294
rect 36206 19234 36258 19246
rect 11218 19182 11230 19234
rect 11282 19182 11294 19234
rect 36206 19170 36258 19182
rect 42478 19234 42530 19246
rect 42478 19170 42530 19182
rect 6190 19122 6242 19134
rect 38894 19122 38946 19134
rect 11442 19070 11454 19122
rect 11506 19070 11518 19122
rect 13794 19070 13806 19122
rect 13858 19070 13870 19122
rect 6190 19058 6242 19070
rect 38894 19058 38946 19070
rect 39230 19122 39282 19134
rect 41358 19122 41410 19134
rect 39554 19070 39566 19122
rect 39618 19070 39630 19122
rect 39230 19058 39282 19070
rect 41358 19058 41410 19070
rect 41582 19122 41634 19134
rect 41582 19058 41634 19070
rect 41918 19122 41970 19134
rect 41918 19058 41970 19070
rect 42142 19122 42194 19134
rect 42142 19058 42194 19070
rect 42366 19122 42418 19134
rect 42366 19058 42418 19070
rect 6862 19010 6914 19022
rect 6862 18946 6914 18958
rect 14142 19010 14194 19022
rect 14142 18946 14194 18958
rect 14590 19010 14642 19022
rect 14590 18946 14642 18958
rect 35646 19010 35698 19022
rect 35646 18946 35698 18958
rect 35870 19010 35922 19022
rect 35870 18946 35922 18958
rect 36094 19010 36146 19022
rect 36094 18946 36146 18958
rect 1344 18842 44576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 44576 18842
rect 1344 18756 44576 18790
rect 5630 18674 5682 18686
rect 5630 18610 5682 18622
rect 6974 18674 7026 18686
rect 34862 18674 34914 18686
rect 20178 18622 20190 18674
rect 20242 18622 20254 18674
rect 6974 18610 7026 18622
rect 34862 18610 34914 18622
rect 35198 18674 35250 18686
rect 35198 18610 35250 18622
rect 41246 18674 41298 18686
rect 41246 18610 41298 18622
rect 40910 18562 40962 18574
rect 9538 18510 9550 18562
rect 9602 18510 9614 18562
rect 14802 18510 14814 18562
rect 14866 18510 14878 18562
rect 40910 18498 40962 18510
rect 41022 18562 41074 18574
rect 41022 18498 41074 18510
rect 41582 18562 41634 18574
rect 41582 18498 41634 18510
rect 41694 18562 41746 18574
rect 41694 18498 41746 18510
rect 5854 18450 5906 18462
rect 6750 18450 6802 18462
rect 4946 18398 4958 18450
rect 5010 18398 5022 18450
rect 6178 18398 6190 18450
rect 6242 18398 6254 18450
rect 6514 18398 6526 18450
rect 6578 18398 6590 18450
rect 5854 18386 5906 18398
rect 6750 18386 6802 18398
rect 6862 18450 6914 18462
rect 9886 18450 9938 18462
rect 7186 18398 7198 18450
rect 7250 18398 7262 18450
rect 7522 18398 7534 18450
rect 7586 18398 7598 18450
rect 6862 18386 6914 18398
rect 9886 18386 9938 18398
rect 11678 18450 11730 18462
rect 11678 18386 11730 18398
rect 11902 18450 11954 18462
rect 11902 18386 11954 18398
rect 12350 18450 12402 18462
rect 35310 18450 35362 18462
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 22418 18398 22430 18450
rect 22482 18398 22494 18450
rect 23202 18398 23214 18450
rect 23266 18398 23278 18450
rect 29810 18398 29822 18450
rect 29874 18398 29886 18450
rect 12350 18386 12402 18398
rect 35310 18386 35362 18398
rect 35646 18450 35698 18462
rect 37214 18450 37266 18462
rect 36082 18398 36094 18450
rect 36146 18398 36158 18450
rect 35646 18386 35698 18398
rect 37214 18386 37266 18398
rect 5742 18338 5794 18350
rect 5742 18274 5794 18286
rect 23662 18338 23714 18350
rect 23662 18274 23714 18286
rect 30046 18338 30098 18350
rect 36418 18286 36430 18338
rect 36482 18286 36494 18338
rect 30046 18274 30098 18286
rect 4958 18226 5010 18238
rect 4958 18162 5010 18174
rect 5294 18226 5346 18238
rect 5294 18162 5346 18174
rect 7758 18226 7810 18238
rect 7758 18162 7810 18174
rect 7982 18226 8034 18238
rect 7982 18162 8034 18174
rect 8094 18226 8146 18238
rect 30158 18226 30210 18238
rect 11330 18174 11342 18226
rect 11394 18174 11406 18226
rect 8094 18162 8146 18174
rect 30158 18162 30210 18174
rect 35198 18226 35250 18238
rect 35198 18162 35250 18174
rect 41582 18226 41634 18238
rect 41582 18162 41634 18174
rect 1344 18058 44576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 44576 18058
rect 1344 17972 44576 18006
rect 19182 17778 19234 17790
rect 34862 17778 34914 17790
rect 36430 17778 36482 17790
rect 2594 17726 2606 17778
rect 2658 17726 2670 17778
rect 4722 17726 4734 17778
rect 4786 17726 4798 17778
rect 27346 17726 27358 17778
rect 27410 17726 27422 17778
rect 33170 17726 33182 17778
rect 33234 17726 33246 17778
rect 35186 17726 35198 17778
rect 35250 17726 35262 17778
rect 19182 17714 19234 17726
rect 34862 17714 34914 17726
rect 36430 17714 36482 17726
rect 6414 17666 6466 17678
rect 1922 17614 1934 17666
rect 1986 17614 1998 17666
rect 5730 17614 5742 17666
rect 5794 17614 5806 17666
rect 6414 17602 6466 17614
rect 6974 17666 7026 17678
rect 6974 17602 7026 17614
rect 7310 17666 7362 17678
rect 7310 17602 7362 17614
rect 18062 17666 18114 17678
rect 40350 17666 40402 17678
rect 18610 17614 18622 17666
rect 18674 17614 18686 17666
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 24546 17614 24558 17666
rect 24610 17614 24622 17666
rect 30146 17614 30158 17666
rect 30210 17614 30222 17666
rect 35298 17614 35310 17666
rect 35362 17614 35374 17666
rect 35522 17614 35534 17666
rect 35586 17614 35598 17666
rect 18062 17602 18114 17614
rect 40350 17602 40402 17614
rect 41582 17666 41634 17678
rect 41582 17602 41634 17614
rect 6526 17554 6578 17566
rect 5954 17502 5966 17554
rect 6018 17502 6030 17554
rect 6526 17490 6578 17502
rect 18174 17554 18226 17566
rect 18174 17490 18226 17502
rect 18286 17554 18338 17566
rect 18286 17490 18338 17502
rect 23998 17554 24050 17566
rect 23998 17490 24050 17502
rect 24110 17554 24162 17566
rect 35758 17554 35810 17566
rect 25218 17502 25230 17554
rect 25282 17502 25294 17554
rect 24110 17490 24162 17502
rect 35758 17490 35810 17502
rect 35982 17554 36034 17566
rect 35982 17490 36034 17502
rect 36990 17554 37042 17566
rect 36990 17490 37042 17502
rect 37326 17554 37378 17566
rect 40910 17554 40962 17566
rect 37426 17502 37438 17554
rect 37490 17502 37502 17554
rect 37326 17490 37378 17502
rect 40910 17490 40962 17502
rect 41134 17554 41186 17566
rect 41134 17490 41186 17502
rect 6750 17442 6802 17454
rect 6750 17378 6802 17390
rect 7086 17442 7138 17454
rect 7086 17378 7138 17390
rect 17950 17442 18002 17454
rect 17950 17378 18002 17390
rect 27806 17442 27858 17454
rect 27806 17378 27858 17390
rect 28590 17442 28642 17454
rect 28590 17378 28642 17390
rect 34750 17442 34802 17454
rect 34750 17378 34802 17390
rect 37102 17442 37154 17454
rect 37102 17378 37154 17390
rect 37214 17442 37266 17454
rect 37214 17378 37266 17390
rect 40462 17442 40514 17454
rect 40462 17378 40514 17390
rect 40686 17442 40738 17454
rect 40686 17378 40738 17390
rect 41246 17442 41298 17454
rect 41246 17378 41298 17390
rect 1344 17274 44576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 44576 17274
rect 1344 17188 44576 17222
rect 4958 17106 5010 17118
rect 4958 17042 5010 17054
rect 17950 17106 18002 17118
rect 17950 17042 18002 17054
rect 20638 17106 20690 17118
rect 20638 17042 20690 17054
rect 17502 16994 17554 17006
rect 27694 16994 27746 17006
rect 32510 16994 32562 17006
rect 13570 16942 13582 16994
rect 13634 16942 13646 16994
rect 22530 16942 22542 16994
rect 22594 16942 22606 16994
rect 31266 16942 31278 16994
rect 31330 16942 31342 16994
rect 36754 16942 36766 16994
rect 36818 16942 36830 16994
rect 17502 16930 17554 16942
rect 27694 16930 27746 16942
rect 32510 16930 32562 16942
rect 16606 16882 16658 16894
rect 11666 16830 11678 16882
rect 11730 16830 11742 16882
rect 16606 16818 16658 16830
rect 17838 16882 17890 16894
rect 20974 16882 21026 16894
rect 22990 16882 23042 16894
rect 19730 16830 19742 16882
rect 19794 16830 19806 16882
rect 22306 16830 22318 16882
rect 22370 16830 22382 16882
rect 28354 16830 28366 16882
rect 28418 16830 28430 16882
rect 32050 16830 32062 16882
rect 32114 16830 32126 16882
rect 33282 16830 33294 16882
rect 33346 16830 33358 16882
rect 17838 16818 17890 16830
rect 20974 16818 21026 16830
rect 22990 16818 23042 16830
rect 20078 16770 20130 16782
rect 28578 16718 28590 16770
rect 28642 16718 28654 16770
rect 29138 16718 29150 16770
rect 29202 16718 29214 16770
rect 20078 16706 20130 16718
rect 17390 16658 17442 16670
rect 17390 16594 17442 16606
rect 17950 16658 18002 16670
rect 17950 16594 18002 16606
rect 19742 16658 19794 16670
rect 19742 16594 19794 16606
rect 1344 16490 44576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 44576 16490
rect 1344 16404 44576 16438
rect 24770 16270 24782 16322
rect 24834 16270 24846 16322
rect 9102 16210 9154 16222
rect 9102 16146 9154 16158
rect 12350 16210 12402 16222
rect 21422 16210 21474 16222
rect 37102 16210 37154 16222
rect 18498 16158 18510 16210
rect 18562 16158 18574 16210
rect 34290 16158 34302 16210
rect 34354 16158 34366 16210
rect 36418 16158 36430 16210
rect 36482 16158 36494 16210
rect 41234 16158 41246 16210
rect 41298 16158 41310 16210
rect 43362 16158 43374 16210
rect 43426 16158 43438 16210
rect 12350 16146 12402 16158
rect 21422 16146 21474 16158
rect 37102 16146 37154 16158
rect 7422 16098 7474 16110
rect 7422 16034 7474 16046
rect 7758 16098 7810 16110
rect 7758 16034 7810 16046
rect 7870 16098 7922 16110
rect 10782 16098 10834 16110
rect 8194 16046 8206 16098
rect 8258 16046 8270 16098
rect 7870 16034 7922 16046
rect 10782 16034 10834 16046
rect 12686 16098 12738 16110
rect 12686 16034 12738 16046
rect 13022 16098 13074 16110
rect 26910 16098 26962 16110
rect 15474 16046 15486 16098
rect 15538 16046 15550 16098
rect 25554 16046 25566 16098
rect 25618 16046 25630 16098
rect 29138 16046 29150 16098
rect 29202 16046 29214 16098
rect 32946 16046 32958 16098
rect 33010 16046 33022 16098
rect 33618 16046 33630 16098
rect 33682 16046 33694 16098
rect 40450 16046 40462 16098
rect 40514 16046 40526 16098
rect 13022 16034 13074 16046
rect 26910 16034 26962 16046
rect 8542 15986 8594 15998
rect 8542 15922 8594 15934
rect 8654 15986 8706 15998
rect 8654 15922 8706 15934
rect 25230 15986 25282 15998
rect 25230 15922 25282 15934
rect 25342 15986 25394 15998
rect 32286 15986 32338 15998
rect 26114 15934 26126 15986
rect 26178 15934 26190 15986
rect 26786 15934 26798 15986
rect 26850 15934 26862 15986
rect 29250 15934 29262 15986
rect 29314 15934 29326 15986
rect 25342 15922 25394 15934
rect 32286 15922 32338 15934
rect 7534 15874 7586 15886
rect 12798 15874 12850 15886
rect 40126 15874 40178 15886
rect 10434 15822 10446 15874
rect 10498 15822 10510 15874
rect 26562 15822 26574 15874
rect 26626 15822 26638 15874
rect 29362 15822 29374 15874
rect 29426 15822 29438 15874
rect 7534 15810 7586 15822
rect 12798 15810 12850 15822
rect 40126 15810 40178 15822
rect 1344 15706 44576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 44576 15706
rect 1344 15620 44576 15654
rect 9662 15538 9714 15550
rect 8866 15486 8878 15538
rect 8930 15486 8942 15538
rect 9662 15474 9714 15486
rect 14366 15538 14418 15550
rect 14366 15474 14418 15486
rect 21870 15538 21922 15550
rect 21870 15474 21922 15486
rect 30270 15538 30322 15550
rect 30270 15474 30322 15486
rect 30606 15538 30658 15550
rect 30606 15474 30658 15486
rect 33294 15538 33346 15550
rect 33294 15474 33346 15486
rect 5742 15426 5794 15438
rect 2706 15374 2718 15426
rect 2770 15374 2782 15426
rect 5742 15362 5794 15374
rect 7758 15426 7810 15438
rect 7758 15362 7810 15374
rect 9886 15426 9938 15438
rect 30158 15426 30210 15438
rect 14018 15374 14030 15426
rect 14082 15374 14094 15426
rect 9886 15362 9938 15374
rect 30158 15362 30210 15374
rect 37438 15426 37490 15438
rect 37438 15362 37490 15374
rect 6862 15314 6914 15326
rect 1922 15262 1934 15314
rect 1986 15262 1998 15314
rect 6862 15250 6914 15262
rect 7310 15314 7362 15326
rect 7310 15250 7362 15262
rect 9550 15314 9602 15326
rect 9550 15250 9602 15262
rect 9998 15314 10050 15326
rect 9998 15250 10050 15262
rect 13694 15314 13746 15326
rect 13694 15250 13746 15262
rect 30382 15314 30434 15326
rect 30382 15250 30434 15262
rect 13134 15202 13186 15214
rect 4834 15150 4846 15202
rect 4898 15150 4910 15202
rect 13134 15138 13186 15150
rect 14814 15202 14866 15214
rect 29598 15202 29650 15214
rect 21746 15150 21758 15202
rect 21810 15150 21822 15202
rect 14814 15138 14866 15150
rect 29598 15138 29650 15150
rect 29822 15202 29874 15214
rect 29822 15138 29874 15150
rect 22094 15090 22146 15102
rect 37550 15090 37602 15102
rect 29250 15038 29262 15090
rect 29314 15038 29326 15090
rect 22094 15026 22146 15038
rect 37550 15026 37602 15038
rect 1344 14922 44576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 44576 14922
rect 1344 14836 44576 14870
rect 9998 14754 10050 14766
rect 29474 14702 29486 14754
rect 29538 14751 29550 14754
rect 29922 14751 29934 14754
rect 29538 14705 29934 14751
rect 29538 14702 29550 14705
rect 29922 14702 29934 14705
rect 29986 14702 29998 14754
rect 9998 14690 10050 14702
rect 18510 14642 18562 14654
rect 15922 14590 15934 14642
rect 15986 14590 15998 14642
rect 18050 14590 18062 14642
rect 18114 14590 18126 14642
rect 18510 14578 18562 14590
rect 25790 14642 25842 14654
rect 25790 14578 25842 14590
rect 29934 14642 29986 14654
rect 38098 14590 38110 14642
rect 38162 14590 38174 14642
rect 40226 14590 40238 14642
rect 40290 14590 40302 14642
rect 29934 14578 29986 14590
rect 9986 14478 9998 14530
rect 10050 14478 10062 14530
rect 15250 14478 15262 14530
rect 15314 14478 15326 14530
rect 37314 14478 37326 14530
rect 37378 14478 37390 14530
rect 9662 14418 9714 14430
rect 9662 14354 9714 14366
rect 5070 14306 5122 14318
rect 5070 14242 5122 14254
rect 13470 14306 13522 14318
rect 14254 14306 14306 14318
rect 13794 14254 13806 14306
rect 13858 14254 13870 14306
rect 13470 14242 13522 14254
rect 14254 14242 14306 14254
rect 36430 14306 36482 14318
rect 36430 14242 36482 14254
rect 1344 14138 44576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 44576 14138
rect 1344 14052 44576 14086
rect 8094 13970 8146 13982
rect 7746 13918 7758 13970
rect 7810 13918 7822 13970
rect 8094 13906 8146 13918
rect 19518 13970 19570 13982
rect 19518 13906 19570 13918
rect 34414 13970 34466 13982
rect 34414 13906 34466 13918
rect 20626 13806 20638 13858
rect 20690 13806 20702 13858
rect 26114 13806 26126 13858
rect 26178 13806 26190 13858
rect 19842 13694 19854 13746
rect 19906 13694 19918 13746
rect 24658 13694 24670 13746
rect 24722 13694 24734 13746
rect 26338 13694 26350 13746
rect 26402 13694 26414 13746
rect 24334 13634 24386 13646
rect 22754 13582 22766 13634
rect 22818 13582 22830 13634
rect 24334 13570 24386 13582
rect 24670 13522 24722 13534
rect 24670 13458 24722 13470
rect 25230 13522 25282 13534
rect 25230 13458 25282 13470
rect 25342 13522 25394 13534
rect 25342 13458 25394 13470
rect 25566 13522 25618 13534
rect 25566 13458 25618 13470
rect 25678 13522 25730 13534
rect 25678 13458 25730 13470
rect 1344 13354 44576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 44576 13354
rect 1344 13268 44576 13302
rect 29486 13186 29538 13198
rect 29486 13122 29538 13134
rect 22866 13022 22878 13074
rect 22930 13022 22942 13074
rect 24994 13022 25006 13074
rect 25058 13022 25070 13074
rect 35186 13022 35198 13074
rect 35250 13022 35262 13074
rect 7982 12962 8034 12974
rect 7746 12910 7758 12962
rect 7810 12910 7822 12962
rect 7982 12898 8034 12910
rect 8094 12962 8146 12974
rect 29710 12962 29762 12974
rect 30382 12962 30434 12974
rect 25778 12910 25790 12962
rect 25842 12910 25854 12962
rect 29922 12910 29934 12962
rect 29986 12910 29998 12962
rect 8094 12898 8146 12910
rect 29710 12898 29762 12910
rect 30382 12898 30434 12910
rect 30830 12962 30882 12974
rect 30830 12898 30882 12910
rect 33294 12962 33346 12974
rect 34750 12962 34802 12974
rect 33954 12910 33966 12962
rect 34018 12910 34030 12962
rect 33294 12898 33346 12910
rect 34750 12898 34802 12910
rect 29374 12850 29426 12862
rect 29374 12786 29426 12798
rect 30270 12850 30322 12862
rect 30270 12786 30322 12798
rect 30606 12850 30658 12862
rect 30606 12786 30658 12798
rect 32846 12850 32898 12862
rect 32846 12786 32898 12798
rect 33182 12850 33234 12862
rect 33182 12786 33234 12798
rect 26238 12738 26290 12750
rect 8530 12686 8542 12738
rect 8594 12686 8606 12738
rect 26238 12674 26290 12686
rect 33070 12738 33122 12750
rect 33070 12674 33122 12686
rect 33742 12738 33794 12750
rect 33742 12674 33794 12686
rect 1344 12570 44576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 44576 12570
rect 1344 12484 44576 12518
rect 6302 12402 6354 12414
rect 6302 12338 6354 12350
rect 9662 12402 9714 12414
rect 9662 12338 9714 12350
rect 16046 12402 16098 12414
rect 16046 12338 16098 12350
rect 16830 12402 16882 12414
rect 16830 12338 16882 12350
rect 7646 12290 7698 12302
rect 2594 12238 2606 12290
rect 2658 12238 2670 12290
rect 7646 12226 7698 12238
rect 8766 12290 8818 12302
rect 8766 12226 8818 12238
rect 12238 12290 12290 12302
rect 12238 12226 12290 12238
rect 12798 12290 12850 12302
rect 28802 12238 28814 12290
rect 28866 12238 28878 12290
rect 35186 12238 35198 12290
rect 35250 12238 35262 12290
rect 12798 12226 12850 12238
rect 7534 12178 7586 12190
rect 1922 12126 1934 12178
rect 1986 12126 1998 12178
rect 6066 12126 6078 12178
rect 6130 12126 6142 12178
rect 7534 12114 7586 12126
rect 7870 12178 7922 12190
rect 8654 12178 8706 12190
rect 8306 12126 8318 12178
rect 8370 12126 8382 12178
rect 7870 12114 7922 12126
rect 8654 12114 8706 12126
rect 11566 12178 11618 12190
rect 11566 12114 11618 12126
rect 11902 12178 11954 12190
rect 11902 12114 11954 12126
rect 15934 12178 15986 12190
rect 25230 12178 25282 12190
rect 20514 12126 20526 12178
rect 20578 12126 20590 12178
rect 15934 12114 15986 12126
rect 25230 12114 25282 12126
rect 25454 12178 25506 12190
rect 31390 12178 31442 12190
rect 28130 12126 28142 12178
rect 28194 12126 28206 12178
rect 35858 12126 35870 12178
rect 35922 12126 35934 12178
rect 25454 12114 25506 12126
rect 31390 12114 31442 12126
rect 5182 12066 5234 12078
rect 4722 12014 4734 12066
rect 4786 12014 4798 12066
rect 5182 12002 5234 12014
rect 11790 12066 11842 12078
rect 11790 12002 11842 12014
rect 14814 12066 14866 12078
rect 36430 12066 36482 12078
rect 17714 12014 17726 12066
rect 17778 12014 17790 12066
rect 19842 12014 19854 12066
rect 19906 12014 19918 12066
rect 30930 12014 30942 12066
rect 30994 12014 31006 12066
rect 33058 12014 33070 12066
rect 33122 12014 33134 12066
rect 14814 12002 14866 12014
rect 36430 12002 36482 12014
rect 15038 11954 15090 11966
rect 8082 11902 8094 11954
rect 8146 11902 8158 11954
rect 15038 11890 15090 11902
rect 15262 11954 15314 11966
rect 15262 11890 15314 11902
rect 15710 11954 15762 11966
rect 15710 11890 15762 11902
rect 16046 11954 16098 11966
rect 25778 11902 25790 11954
rect 25842 11902 25854 11954
rect 16046 11890 16098 11902
rect 1344 11786 44576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 44576 11786
rect 1344 11700 44576 11734
rect 13806 11618 13858 11630
rect 29922 11566 29934 11618
rect 29986 11566 29998 11618
rect 13806 11554 13858 11566
rect 9326 11506 9378 11518
rect 8418 11454 8430 11506
rect 8482 11454 8494 11506
rect 9326 11442 9378 11454
rect 17838 11506 17890 11518
rect 17838 11442 17890 11454
rect 17950 11506 18002 11518
rect 17950 11442 18002 11454
rect 32958 11506 33010 11518
rect 32958 11442 33010 11454
rect 6638 11394 6690 11406
rect 6638 11330 6690 11342
rect 6974 11394 7026 11406
rect 6974 11330 7026 11342
rect 7422 11394 7474 11406
rect 12238 11394 12290 11406
rect 7858 11342 7870 11394
rect 7922 11342 7934 11394
rect 8866 11342 8878 11394
rect 8930 11342 8942 11394
rect 7422 11330 7474 11342
rect 12238 11330 12290 11342
rect 16830 11394 16882 11406
rect 16830 11330 16882 11342
rect 17054 11394 17106 11406
rect 17614 11394 17666 11406
rect 17378 11342 17390 11394
rect 17442 11342 17454 11394
rect 17054 11330 17106 11342
rect 17614 11330 17666 11342
rect 18062 11394 18114 11406
rect 18062 11330 18114 11342
rect 18286 11394 18338 11406
rect 32510 11394 32562 11406
rect 30706 11342 30718 11394
rect 30770 11342 30782 11394
rect 18286 11330 18338 11342
rect 32510 11330 32562 11342
rect 32846 11394 32898 11406
rect 32846 11330 32898 11342
rect 33518 11394 33570 11406
rect 33518 11330 33570 11342
rect 7198 11282 7250 11294
rect 7198 11218 7250 11230
rect 8430 11282 8482 11294
rect 8430 11218 8482 11230
rect 12350 11282 12402 11294
rect 12350 11218 12402 11230
rect 13694 11282 13746 11294
rect 13694 11218 13746 11230
rect 16718 11282 16770 11294
rect 16718 11218 16770 11230
rect 18622 11282 18674 11294
rect 18622 11218 18674 11230
rect 30382 11282 30434 11294
rect 30382 11218 30434 11230
rect 30494 11282 30546 11294
rect 30494 11218 30546 11230
rect 33070 11282 33122 11294
rect 33070 11218 33122 11230
rect 6750 11170 6802 11182
rect 6750 11106 6802 11118
rect 7534 11170 7586 11182
rect 7534 11106 7586 11118
rect 7646 11170 7698 11182
rect 7646 11106 7698 11118
rect 8318 11170 8370 11182
rect 8318 11106 8370 11118
rect 8654 11170 8706 11182
rect 8654 11106 8706 11118
rect 12574 11170 12626 11182
rect 12574 11106 12626 11118
rect 13806 11170 13858 11182
rect 13806 11106 13858 11118
rect 18846 11170 18898 11182
rect 18846 11106 18898 11118
rect 18958 11170 19010 11182
rect 18958 11106 19010 11118
rect 1344 11002 44576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 44576 11002
rect 1344 10916 44576 10950
rect 8318 10834 8370 10846
rect 8318 10770 8370 10782
rect 8542 10834 8594 10846
rect 8542 10770 8594 10782
rect 8654 10834 8706 10846
rect 8654 10770 8706 10782
rect 9102 10834 9154 10846
rect 9102 10770 9154 10782
rect 10222 10722 10274 10734
rect 10222 10658 10274 10670
rect 11790 10722 11842 10734
rect 15934 10722 15986 10734
rect 15138 10670 15150 10722
rect 15202 10670 15214 10722
rect 30370 10670 30382 10722
rect 30434 10670 30446 10722
rect 11790 10658 11842 10670
rect 15934 10658 15986 10670
rect 7198 10610 7250 10622
rect 7198 10546 7250 10558
rect 7422 10610 7474 10622
rect 7422 10546 7474 10558
rect 7870 10610 7922 10622
rect 10446 10610 10498 10622
rect 8082 10558 8094 10610
rect 8146 10558 8158 10610
rect 7870 10546 7922 10558
rect 10446 10546 10498 10558
rect 11230 10610 11282 10622
rect 11230 10546 11282 10558
rect 11342 10610 11394 10622
rect 11342 10546 11394 10558
rect 11566 10610 11618 10622
rect 11566 10546 11618 10558
rect 12574 10610 12626 10622
rect 12574 10546 12626 10558
rect 12686 10610 12738 10622
rect 12686 10546 12738 10558
rect 13806 10610 13858 10622
rect 15710 10610 15762 10622
rect 14354 10558 14366 10610
rect 14418 10558 14430 10610
rect 15250 10558 15262 10610
rect 15314 10558 15326 10610
rect 13806 10546 13858 10558
rect 15710 10546 15762 10558
rect 16382 10610 16434 10622
rect 16382 10546 16434 10558
rect 30046 10610 30098 10622
rect 30046 10546 30098 10558
rect 7310 10498 7362 10510
rect 7310 10434 7362 10446
rect 11454 10498 11506 10510
rect 11454 10434 11506 10446
rect 15822 10498 15874 10510
rect 15822 10434 15874 10446
rect 10782 10386 10834 10398
rect 10782 10322 10834 10334
rect 12910 10386 12962 10398
rect 12910 10322 12962 10334
rect 13022 10386 13074 10398
rect 13022 10322 13074 10334
rect 15374 10386 15426 10398
rect 15374 10322 15426 10334
rect 1344 10218 44576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 44576 10218
rect 1344 10132 44576 10166
rect 6750 10050 6802 10062
rect 6750 9986 6802 9998
rect 29598 10050 29650 10062
rect 29598 9986 29650 9998
rect 29822 10050 29874 10062
rect 29822 9986 29874 9998
rect 16270 9938 16322 9950
rect 16270 9874 16322 9886
rect 23550 9938 23602 9950
rect 23550 9874 23602 9886
rect 24110 9938 24162 9950
rect 24110 9874 24162 9886
rect 12126 9826 12178 9838
rect 7298 9774 7310 9826
rect 7362 9774 7374 9826
rect 12126 9762 12178 9774
rect 12462 9826 12514 9838
rect 12462 9762 12514 9774
rect 12798 9826 12850 9838
rect 16606 9826 16658 9838
rect 13682 9774 13694 9826
rect 13746 9774 13758 9826
rect 14466 9774 14478 9826
rect 14530 9774 14542 9826
rect 12798 9762 12850 9774
rect 16606 9762 16658 9774
rect 19070 9826 19122 9838
rect 19070 9762 19122 9774
rect 19182 9826 19234 9838
rect 19394 9774 19406 9826
rect 19458 9774 19470 9826
rect 29362 9774 29374 9826
rect 29426 9774 29438 9826
rect 19182 9762 19234 9774
rect 6526 9714 6578 9726
rect 6526 9650 6578 9662
rect 7086 9714 7138 9726
rect 23214 9714 23266 9726
rect 13458 9662 13470 9714
rect 13522 9662 13534 9714
rect 14578 9662 14590 9714
rect 14642 9662 14654 9714
rect 18162 9662 18174 9714
rect 18226 9662 18238 9714
rect 7086 9650 7138 9662
rect 23214 9650 23266 9662
rect 29934 9714 29986 9726
rect 29934 9650 29986 9662
rect 6638 9602 6690 9614
rect 6638 9538 6690 9550
rect 7982 9602 8034 9614
rect 7982 9538 8034 9550
rect 12350 9602 12402 9614
rect 19854 9602 19906 9614
rect 18610 9550 18622 9602
rect 18674 9550 18686 9602
rect 12350 9538 12402 9550
rect 19854 9538 19906 9550
rect 23438 9602 23490 9614
rect 23438 9538 23490 9550
rect 23662 9602 23714 9614
rect 23662 9538 23714 9550
rect 1344 9434 44576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 44576 9434
rect 1344 9348 44576 9382
rect 16382 9266 16434 9278
rect 14242 9214 14254 9266
rect 14306 9214 14318 9266
rect 16382 9202 16434 9214
rect 21422 9266 21474 9278
rect 21422 9202 21474 9214
rect 27470 9266 27522 9278
rect 28914 9214 28926 9266
rect 28978 9214 28990 9266
rect 27470 9202 27522 9214
rect 16494 9154 16546 9166
rect 27582 9154 27634 9166
rect 4498 9102 4510 9154
rect 4562 9102 4574 9154
rect 25330 9102 25342 9154
rect 25394 9102 25406 9154
rect 16494 9090 16546 9102
rect 27582 9090 27634 9102
rect 28366 9154 28418 9166
rect 28366 9090 28418 9102
rect 7086 9042 7138 9054
rect 3826 8990 3838 9042
rect 3890 8990 3902 9042
rect 7086 8978 7138 8990
rect 14590 9042 14642 9054
rect 25678 9042 25730 9054
rect 21858 8990 21870 9042
rect 21922 8990 21934 9042
rect 14590 8978 14642 8990
rect 25678 8978 25730 8990
rect 27134 9042 27186 9054
rect 27134 8978 27186 8990
rect 27806 9042 27858 9054
rect 27806 8978 27858 8990
rect 28254 9042 28306 9054
rect 28254 8978 28306 8990
rect 28478 9042 28530 9054
rect 28478 8978 28530 8990
rect 6626 8878 6638 8930
rect 6690 8878 6702 8930
rect 22530 8878 22542 8930
rect 22594 8878 22606 8930
rect 24658 8878 24670 8930
rect 24722 8878 24734 8930
rect 1344 8650 44576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 44576 8650
rect 1344 8564 44576 8598
rect 12350 8482 12402 8494
rect 12350 8418 12402 8430
rect 11118 8370 11170 8382
rect 10770 8318 10782 8370
rect 10834 8318 10846 8370
rect 11118 8306 11170 8318
rect 11566 8370 11618 8382
rect 23102 8370 23154 8382
rect 12674 8318 12686 8370
rect 12738 8318 12750 8370
rect 29474 8318 29486 8370
rect 29538 8318 29550 8370
rect 31602 8318 31614 8370
rect 31666 8318 31678 8370
rect 11566 8306 11618 8318
rect 23102 8306 23154 8318
rect 22654 8258 22706 8270
rect 18274 8206 18286 8258
rect 18338 8206 18350 8258
rect 22654 8194 22706 8206
rect 22990 8258 23042 8270
rect 22990 8194 23042 8206
rect 23326 8258 23378 8270
rect 23326 8194 23378 8206
rect 23550 8258 23602 8270
rect 32958 8258 33010 8270
rect 27794 8206 27806 8258
rect 27858 8206 27870 8258
rect 32386 8206 32398 8258
rect 32450 8206 32462 8258
rect 23550 8194 23602 8206
rect 32958 8194 33010 8206
rect 10894 8146 10946 8158
rect 10894 8082 10946 8094
rect 12574 8146 12626 8158
rect 27570 8094 27582 8146
rect 27634 8094 27646 8146
rect 12574 8082 12626 8094
rect 13582 8034 13634 8046
rect 13582 7970 13634 7982
rect 18510 8034 18562 8046
rect 18510 7970 18562 7982
rect 22430 8034 22482 8046
rect 22430 7970 22482 7982
rect 22542 8034 22594 8046
rect 22542 7970 22594 7982
rect 1344 7866 44576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 44576 7866
rect 1344 7780 44576 7814
rect 22990 7698 23042 7710
rect 22990 7634 23042 7646
rect 27582 7698 27634 7710
rect 27582 7634 27634 7646
rect 26686 7586 26738 7598
rect 19506 7534 19518 7586
rect 19570 7534 19582 7586
rect 26686 7522 26738 7534
rect 28702 7586 28754 7598
rect 28702 7522 28754 7534
rect 27694 7474 27746 7486
rect 20290 7422 20302 7474
rect 20354 7422 20366 7474
rect 28242 7422 28254 7474
rect 28306 7422 28318 7474
rect 27694 7410 27746 7422
rect 20750 7362 20802 7374
rect 17378 7310 17390 7362
rect 17442 7310 17454 7362
rect 20750 7298 20802 7310
rect 1344 7082 44576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 44576 7082
rect 1344 6996 44576 7030
rect 26798 6914 26850 6926
rect 26798 6850 26850 6862
rect 10658 6750 10670 6802
rect 10722 6750 10734 6802
rect 12786 6750 12798 6802
rect 12850 6750 12862 6802
rect 13582 6690 13634 6702
rect 9986 6638 9998 6690
rect 10050 6638 10062 6690
rect 13582 6626 13634 6638
rect 25902 6690 25954 6702
rect 27470 6690 27522 6702
rect 26786 6638 26798 6690
rect 26850 6638 26862 6690
rect 25902 6626 25954 6638
rect 27470 6626 27522 6638
rect 26238 6578 26290 6590
rect 26238 6514 26290 6526
rect 26350 6578 26402 6590
rect 26350 6514 26402 6526
rect 27134 6578 27186 6590
rect 27134 6514 27186 6526
rect 27806 6578 27858 6590
rect 27806 6514 27858 6526
rect 26574 6466 26626 6478
rect 26574 6402 26626 6414
rect 27582 6466 27634 6478
rect 27582 6402 27634 6414
rect 1344 6298 44576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 44576 6298
rect 1344 6212 44576 6246
rect 15374 6130 15426 6142
rect 15374 6066 15426 6078
rect 25902 6130 25954 6142
rect 25902 6066 25954 6078
rect 26462 6018 26514 6030
rect 12786 5966 12798 6018
rect 12850 5966 12862 6018
rect 26462 5954 26514 5966
rect 27134 6018 27186 6030
rect 27134 5954 27186 5966
rect 27358 6018 27410 6030
rect 27358 5954 27410 5966
rect 28030 6018 28082 6030
rect 28030 5954 28082 5966
rect 23102 5906 23154 5918
rect 12114 5854 12126 5906
rect 12178 5854 12190 5906
rect 23102 5842 23154 5854
rect 25678 5906 25730 5918
rect 25678 5842 25730 5854
rect 26014 5906 26066 5918
rect 26014 5842 26066 5854
rect 23326 5794 23378 5806
rect 14914 5742 14926 5794
rect 14978 5742 14990 5794
rect 27458 5742 27470 5794
rect 27522 5742 27534 5794
rect 23326 5730 23378 5742
rect 26350 5682 26402 5694
rect 22754 5630 22766 5682
rect 22818 5630 22830 5682
rect 26350 5618 26402 5630
rect 27806 5682 27858 5694
rect 27806 5618 27858 5630
rect 28142 5682 28194 5694
rect 28142 5618 28194 5630
rect 1344 5514 44576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 44576 5514
rect 1344 5428 44576 5462
rect 24546 5182 24558 5234
rect 24610 5182 24622 5234
rect 20862 5122 20914 5134
rect 21634 5070 21646 5122
rect 21698 5070 21710 5122
rect 20862 5058 20914 5070
rect 22418 4958 22430 5010
rect 22482 4958 22494 5010
rect 1344 4730 44576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 44576 4730
rect 1344 4644 44576 4678
rect 22430 4562 22482 4574
rect 22430 4498 22482 4510
rect 30270 4562 30322 4574
rect 30270 4498 30322 4510
rect 22766 4450 22818 4462
rect 27682 4398 27694 4450
rect 27746 4398 27758 4450
rect 22766 4386 22818 4398
rect 27010 4286 27022 4338
rect 27074 4286 27086 4338
rect 29810 4174 29822 4226
rect 29874 4174 29886 4226
rect 1344 3946 44576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 44576 3946
rect 1344 3860 44576 3894
rect 1344 3162 44576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 44576 3162
rect 1344 3076 44576 3110
<< via1 >>
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 18286 42142 18338 42194
rect 33518 42142 33570 42194
rect 6190 42030 6242 42082
rect 9998 42030 10050 42082
rect 5070 41918 5122 41970
rect 5854 41918 5906 41970
rect 8878 41918 8930 41970
rect 9662 41918 9714 41970
rect 13470 41918 13522 41970
rect 17278 41918 17330 41970
rect 21086 41918 21138 41970
rect 24894 41918 24946 41970
rect 30830 41918 30882 41970
rect 32622 41918 32674 41970
rect 36318 41918 36370 41970
rect 40350 41918 40402 41970
rect 14478 41806 14530 41858
rect 22094 41806 22146 41858
rect 25902 41806 25954 41858
rect 28926 41806 28978 41858
rect 37326 41806 37378 41858
rect 41134 41806 41186 41858
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 43598 41246 43650 41298
rect 41582 41134 41634 41186
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 24334 40574 24386 40626
rect 5630 40462 5682 40514
rect 8766 40462 8818 40514
rect 4958 40350 5010 40402
rect 8318 40350 8370 40402
rect 9774 40350 9826 40402
rect 13358 40350 13410 40402
rect 16942 40350 16994 40402
rect 17614 40350 17666 40402
rect 23662 40350 23714 40402
rect 24110 40350 24162 40402
rect 27806 40350 27858 40402
rect 28478 40350 28530 40402
rect 31166 40350 31218 40402
rect 33182 40350 33234 40402
rect 36430 40350 36482 40402
rect 40462 40350 40514 40402
rect 41022 40350 41074 40402
rect 7758 40238 7810 40290
rect 10558 40238 10610 40290
rect 12686 40238 12738 40290
rect 14030 40238 14082 40290
rect 16158 40238 16210 40290
rect 18398 40238 18450 40290
rect 20526 40238 20578 40290
rect 24222 40238 24274 40290
rect 25454 40238 25506 40290
rect 30606 40238 30658 40290
rect 33854 40238 33906 40290
rect 35982 40238 36034 40290
rect 41806 40238 41858 40290
rect 43934 40238 43986 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 4734 39678 4786 39730
rect 5742 39678 5794 39730
rect 8766 39678 8818 39730
rect 18398 39678 18450 39730
rect 18958 39678 19010 39730
rect 20190 39678 20242 39730
rect 23550 39678 23602 39730
rect 25678 39678 25730 39730
rect 32622 39678 32674 39730
rect 33070 39678 33122 39730
rect 39230 39678 39282 39730
rect 1822 39566 1874 39618
rect 17950 39566 18002 39618
rect 19518 39566 19570 39618
rect 26462 39566 26514 39618
rect 26910 39566 26962 39618
rect 29822 39566 29874 39618
rect 42030 39566 42082 39618
rect 2606 39454 2658 39506
rect 14590 39454 14642 39506
rect 14926 39454 14978 39506
rect 18510 39454 18562 39506
rect 19070 39454 19122 39506
rect 19854 39454 19906 39506
rect 30494 39454 30546 39506
rect 41358 39454 41410 39506
rect 8878 39342 8930 39394
rect 12910 39342 12962 39394
rect 16382 39342 16434 39394
rect 18286 39342 18338 39394
rect 18846 39342 18898 39394
rect 20078 39342 20130 39394
rect 20302 39342 20354 39394
rect 38894 39342 38946 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 20302 39006 20354 39058
rect 24782 39006 24834 39058
rect 25790 39006 25842 39058
rect 26462 39006 26514 39058
rect 38334 39006 38386 39058
rect 41358 39006 41410 39058
rect 41470 39006 41522 39058
rect 41694 39006 41746 39058
rect 20526 38894 20578 38946
rect 24110 38894 24162 38946
rect 24446 38894 24498 38946
rect 24558 38894 24610 38946
rect 27134 38894 27186 38946
rect 39902 38894 39954 38946
rect 20190 38782 20242 38834
rect 25566 38782 25618 38834
rect 25790 38782 25842 38834
rect 26126 38782 26178 38834
rect 26686 38782 26738 38834
rect 27246 38782 27298 38834
rect 37550 38782 37602 38834
rect 37774 38782 37826 38834
rect 38110 38782 38162 38834
rect 39790 38782 39842 38834
rect 40126 38782 40178 38834
rect 40798 38782 40850 38834
rect 41134 38782 41186 38834
rect 41918 38782 41970 38834
rect 42142 38782 42194 38834
rect 23886 38670 23938 38722
rect 34638 38670 34690 38722
rect 36766 38670 36818 38722
rect 38782 38670 38834 38722
rect 41806 38670 41858 38722
rect 23550 38558 23602 38610
rect 37998 38558 38050 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 20414 38222 20466 38274
rect 24446 38222 24498 38274
rect 25566 38222 25618 38274
rect 5070 38110 5122 38162
rect 5742 38110 5794 38162
rect 7758 38110 7810 38162
rect 16606 38110 16658 38162
rect 18734 38110 18786 38162
rect 23550 38110 23602 38162
rect 25790 38110 25842 38162
rect 2270 37998 2322 38050
rect 10558 37998 10610 38050
rect 11118 37998 11170 38050
rect 15822 37998 15874 38050
rect 24110 37998 24162 38050
rect 24222 37998 24274 38050
rect 37438 37998 37490 38050
rect 40574 37998 40626 38050
rect 2942 37886 2994 37938
rect 9886 37886 9938 37938
rect 19742 37886 19794 37938
rect 20078 37886 20130 37938
rect 20526 37886 20578 37938
rect 23662 37886 23714 37938
rect 26014 37886 26066 37938
rect 37102 37886 37154 37938
rect 37214 37886 37266 37938
rect 40238 37886 40290 37938
rect 40350 37886 40402 37938
rect 41022 37886 41074 37938
rect 41134 37886 41186 37938
rect 41358 37886 41410 37938
rect 19182 37774 19234 37826
rect 23438 37774 23490 37826
rect 26574 37774 26626 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 4622 37438 4674 37490
rect 5070 37438 5122 37490
rect 14254 37438 14306 37490
rect 20414 37438 20466 37490
rect 24110 37438 24162 37490
rect 25230 37438 25282 37490
rect 41358 37438 41410 37490
rect 41134 37326 41186 37378
rect 4398 37214 4450 37266
rect 5630 37214 5682 37266
rect 11006 37214 11058 37266
rect 20750 37214 20802 37266
rect 41022 37214 41074 37266
rect 5182 37102 5234 37154
rect 11678 37102 11730 37154
rect 13806 37102 13858 37154
rect 25790 37102 25842 37154
rect 4734 36990 4786 37042
rect 25566 36990 25618 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 7422 36654 7474 36706
rect 21310 36654 21362 36706
rect 40798 36654 40850 36706
rect 6974 36542 7026 36594
rect 7758 36430 7810 36482
rect 19742 36430 19794 36482
rect 20190 36430 20242 36482
rect 21646 36430 21698 36482
rect 21870 36430 21922 36482
rect 37662 36430 37714 36482
rect 7982 36318 8034 36370
rect 8542 36318 8594 36370
rect 37102 36318 37154 36370
rect 37774 36318 37826 36370
rect 40686 36318 40738 36370
rect 20414 36206 20466 36258
rect 37214 36206 37266 36258
rect 37438 36206 37490 36258
rect 37998 36206 38050 36258
rect 40798 36206 40850 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 24558 35870 24610 35922
rect 19854 35758 19906 35810
rect 20078 35758 20130 35810
rect 23662 35758 23714 35810
rect 29710 35758 29762 35810
rect 37438 35758 37490 35810
rect 40014 35758 40066 35810
rect 23550 35646 23602 35698
rect 24670 35646 24722 35698
rect 30494 35646 30546 35698
rect 30942 35646 30994 35698
rect 36766 35646 36818 35698
rect 37102 35646 37154 35698
rect 37550 35646 37602 35698
rect 38110 35646 38162 35698
rect 39454 35646 39506 35698
rect 39790 35646 39842 35698
rect 40462 35646 40514 35698
rect 40910 35646 40962 35698
rect 9886 35534 9938 35586
rect 27582 35534 27634 35586
rect 33854 35534 33906 35586
rect 35982 35534 36034 35586
rect 37214 35534 37266 35586
rect 40238 35534 40290 35586
rect 41694 35534 41746 35586
rect 43822 35534 43874 35586
rect 20190 35422 20242 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 21422 35086 21474 35138
rect 37102 35086 37154 35138
rect 5070 34974 5122 35026
rect 5742 34974 5794 35026
rect 6974 34974 7026 35026
rect 8542 34974 8594 35026
rect 11006 34974 11058 35026
rect 13806 34974 13858 35026
rect 20638 34974 20690 35026
rect 27134 34974 27186 35026
rect 33406 34974 33458 35026
rect 2270 34862 2322 34914
rect 7310 34862 7362 34914
rect 7646 34862 7698 34914
rect 8430 34862 8482 34914
rect 9326 34862 9378 34914
rect 9550 34862 9602 34914
rect 9774 34862 9826 34914
rect 16606 34862 16658 34914
rect 20190 34862 20242 34914
rect 20414 34862 20466 34914
rect 21310 34862 21362 34914
rect 24446 34862 24498 34914
rect 25230 34862 25282 34914
rect 26686 34862 26738 34914
rect 27022 34862 27074 34914
rect 30606 34862 30658 34914
rect 2942 34750 2994 34802
rect 10110 34750 10162 34802
rect 15934 34750 15986 34802
rect 20750 34750 20802 34802
rect 28030 34750 28082 34802
rect 31278 34750 31330 34802
rect 37102 34750 37154 34802
rect 37214 34750 37266 34802
rect 40686 34750 40738 34802
rect 9998 34638 10050 34690
rect 10670 34638 10722 34690
rect 17166 34638 17218 34690
rect 21422 34638 21474 34690
rect 24222 34638 24274 34690
rect 33854 34638 33906 34690
rect 40350 34638 40402 34690
rect 40574 34638 40626 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 8542 34302 8594 34354
rect 8766 34302 8818 34354
rect 10894 34302 10946 34354
rect 11678 34302 11730 34354
rect 15598 34302 15650 34354
rect 32062 34302 32114 34354
rect 9998 34190 10050 34242
rect 12014 34190 12066 34242
rect 23326 34190 23378 34242
rect 23438 34190 23490 34242
rect 25230 34190 25282 34242
rect 31838 34190 31890 34242
rect 8878 34078 8930 34130
rect 10222 34078 10274 34130
rect 10558 34078 10610 34130
rect 10670 34078 10722 34130
rect 11006 34078 11058 34130
rect 11342 34078 11394 34130
rect 15374 34078 15426 34130
rect 15710 34078 15762 34130
rect 15934 34078 15986 34130
rect 20638 34078 20690 34130
rect 21086 34078 21138 34130
rect 22206 34078 22258 34130
rect 22766 34078 22818 34130
rect 25342 34078 25394 34130
rect 25790 34078 25842 34130
rect 30830 34078 30882 34130
rect 30942 34078 30994 34130
rect 31166 34078 31218 34130
rect 31390 34078 31442 34130
rect 31726 34078 31778 34130
rect 9662 33966 9714 34018
rect 12462 33966 12514 34018
rect 16382 33966 16434 34018
rect 23886 33966 23938 34018
rect 29710 33966 29762 34018
rect 30158 33966 30210 34018
rect 31278 33966 31330 34018
rect 32398 33966 32450 34018
rect 10334 33854 10386 33906
rect 23102 33854 23154 33906
rect 23662 33854 23714 33906
rect 25566 33854 25618 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 6974 33406 7026 33458
rect 11902 33406 11954 33458
rect 12798 33406 12850 33458
rect 15374 33406 15426 33458
rect 34638 33406 34690 33458
rect 43822 33406 43874 33458
rect 8206 33294 8258 33346
rect 12350 33294 12402 33346
rect 25902 33294 25954 33346
rect 26574 33294 26626 33346
rect 40014 33294 40066 33346
rect 40350 33294 40402 33346
rect 40910 33294 40962 33346
rect 7310 33182 7362 33234
rect 7422 33182 7474 33234
rect 11790 33182 11842 33234
rect 12126 33182 12178 33234
rect 15038 33182 15090 33234
rect 15486 33182 15538 33234
rect 25566 33182 25618 33234
rect 40462 33182 40514 33234
rect 41694 33182 41746 33234
rect 7534 33070 7586 33122
rect 7758 33070 7810 33122
rect 10670 33070 10722 33122
rect 14702 33070 14754 33122
rect 15262 33070 15314 33122
rect 17054 33070 17106 33122
rect 26462 33070 26514 33122
rect 35758 33070 35810 33122
rect 35982 33070 36034 33122
rect 36318 33070 36370 33122
rect 40686 33070 40738 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 5630 32734 5682 32786
rect 6638 32734 6690 32786
rect 7870 32734 7922 32786
rect 8542 32734 8594 32786
rect 11790 32734 11842 32786
rect 12126 32734 12178 32786
rect 13022 32734 13074 32786
rect 13918 32734 13970 32786
rect 15486 32734 15538 32786
rect 17614 32734 17666 32786
rect 20302 32734 20354 32786
rect 21758 32734 21810 32786
rect 33742 32734 33794 32786
rect 41694 32734 41746 32786
rect 41806 32734 41858 32786
rect 6862 32622 6914 32674
rect 7758 32622 7810 32674
rect 11902 32622 11954 32674
rect 13582 32622 13634 32674
rect 15822 32622 15874 32674
rect 17838 32622 17890 32674
rect 25790 32622 25842 32674
rect 40798 32622 40850 32674
rect 41022 32622 41074 32674
rect 2270 32510 2322 32562
rect 7086 32510 7138 32562
rect 7310 32510 7362 32562
rect 12462 32510 12514 32562
rect 12686 32510 12738 32562
rect 16046 32510 16098 32562
rect 16494 32510 16546 32562
rect 17278 32510 17330 32562
rect 22206 32510 22258 32562
rect 22430 32510 22482 32562
rect 34190 32510 34242 32562
rect 34974 32510 35026 32562
rect 41134 32510 41186 32562
rect 41470 32510 41522 32562
rect 3054 32398 3106 32450
rect 5182 32398 5234 32450
rect 6974 32398 7026 32450
rect 15038 32398 15090 32450
rect 19406 32398 19458 32450
rect 22654 32398 22706 32450
rect 25678 32398 25730 32450
rect 30494 32398 30546 32450
rect 34638 32398 34690 32450
rect 35758 32398 35810 32450
rect 37886 32398 37938 32450
rect 16270 32286 16322 32338
rect 16942 32286 16994 32338
rect 17950 32286 18002 32338
rect 19630 32286 19682 32338
rect 19854 32286 19906 32338
rect 26014 32286 26066 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 25678 31950 25730 32002
rect 41694 31950 41746 32002
rect 6190 31838 6242 31890
rect 8542 31838 8594 31890
rect 12686 31838 12738 31890
rect 18286 31838 18338 31890
rect 20078 31838 20130 31890
rect 20414 31838 20466 31890
rect 20638 31838 20690 31890
rect 24894 31838 24946 31890
rect 26350 31838 26402 31890
rect 8766 31726 8818 31778
rect 8990 31726 9042 31778
rect 15598 31726 15650 31778
rect 19854 31726 19906 31778
rect 25230 31726 25282 31778
rect 25454 31726 25506 31778
rect 26126 31726 26178 31778
rect 26574 31726 26626 31778
rect 30382 31726 30434 31778
rect 30718 31726 30770 31778
rect 6078 31614 6130 31666
rect 20414 31614 20466 31666
rect 34078 31614 34130 31666
rect 37214 31614 37266 31666
rect 41582 31614 41634 31666
rect 9438 31502 9490 31554
rect 11118 31502 11170 31554
rect 11454 31502 11506 31554
rect 29822 31502 29874 31554
rect 29934 31502 29986 31554
rect 30046 31502 30098 31554
rect 36878 31502 36930 31554
rect 37102 31502 37154 31554
rect 41694 31502 41746 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 6638 31166 6690 31218
rect 10222 31166 10274 31218
rect 18958 31166 19010 31218
rect 25902 31166 25954 31218
rect 26686 31166 26738 31218
rect 34750 31166 34802 31218
rect 35534 31166 35586 31218
rect 39342 31166 39394 31218
rect 40350 31166 40402 31218
rect 12014 31054 12066 31106
rect 29038 31054 29090 31106
rect 35086 31054 35138 31106
rect 10110 30942 10162 30994
rect 15822 30942 15874 30994
rect 19070 30942 19122 30994
rect 19294 30942 19346 30994
rect 19518 30942 19570 30994
rect 25566 30942 25618 30994
rect 26014 30942 26066 30994
rect 26238 30942 26290 30994
rect 26910 30942 26962 30994
rect 29822 30942 29874 30994
rect 30830 30942 30882 30994
rect 34862 30942 34914 30994
rect 35198 30942 35250 30994
rect 35758 30942 35810 30994
rect 36094 30942 36146 30994
rect 39006 30942 39058 30994
rect 40014 30942 40066 30994
rect 9886 30830 9938 30882
rect 16382 30830 16434 30882
rect 20638 30830 20690 30882
rect 26574 30830 26626 30882
rect 31278 30830 31330 30882
rect 35870 30830 35922 30882
rect 38670 30830 38722 30882
rect 10222 30718 10274 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19182 30382 19234 30434
rect 19406 30382 19458 30434
rect 5854 30270 5906 30322
rect 14926 30270 14978 30322
rect 19966 30270 20018 30322
rect 6078 30158 6130 30210
rect 6638 30158 6690 30210
rect 6974 30158 7026 30210
rect 7422 30158 7474 30210
rect 8878 30158 8930 30210
rect 9214 30158 9266 30210
rect 11230 30158 11282 30210
rect 13806 30158 13858 30210
rect 14590 30158 14642 30210
rect 16046 30158 16098 30210
rect 16270 30158 16322 30210
rect 18734 30158 18786 30210
rect 19630 30158 19682 30210
rect 19742 30158 19794 30210
rect 25566 30158 25618 30210
rect 26238 30158 26290 30210
rect 27358 30158 27410 30210
rect 30382 30158 30434 30210
rect 30606 30158 30658 30210
rect 31278 30158 31330 30210
rect 31726 30158 31778 30210
rect 36990 30158 37042 30210
rect 7086 30046 7138 30098
rect 11566 30046 11618 30098
rect 12126 30046 12178 30098
rect 15262 30046 15314 30098
rect 15598 30046 15650 30098
rect 25902 30046 25954 30098
rect 27246 30046 27298 30098
rect 31950 30046 32002 30098
rect 32062 30046 32114 30098
rect 37102 30046 37154 30098
rect 39566 30046 39618 30098
rect 11678 29934 11730 29986
rect 13918 29934 13970 29986
rect 15038 29934 15090 29986
rect 15822 29934 15874 29986
rect 15934 29934 15986 29986
rect 18398 29934 18450 29986
rect 20414 29934 20466 29986
rect 25790 29934 25842 29986
rect 26350 29934 26402 29986
rect 37326 29934 37378 29986
rect 38894 29934 38946 29986
rect 39230 29934 39282 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 5182 29598 5234 29650
rect 9998 29598 10050 29650
rect 14702 29598 14754 29650
rect 32398 29598 32450 29650
rect 10446 29486 10498 29538
rect 11118 29486 11170 29538
rect 14254 29486 14306 29538
rect 14590 29486 14642 29538
rect 16270 29486 16322 29538
rect 25566 29486 25618 29538
rect 26014 29486 26066 29538
rect 31726 29486 31778 29538
rect 33630 29486 33682 29538
rect 1822 29374 1874 29426
rect 5966 29374 6018 29426
rect 9774 29374 9826 29426
rect 10222 29374 10274 29426
rect 11230 29374 11282 29426
rect 11678 29374 11730 29426
rect 15262 29374 15314 29426
rect 15934 29374 15986 29426
rect 16494 29374 16546 29426
rect 25230 29374 25282 29426
rect 26462 29374 26514 29426
rect 26910 29374 26962 29426
rect 31054 29374 31106 29426
rect 31502 29374 31554 29426
rect 32062 29374 32114 29426
rect 33294 29374 33346 29426
rect 33966 29374 34018 29426
rect 40350 29374 40402 29426
rect 40910 29374 40962 29426
rect 2606 29262 2658 29314
rect 4734 29262 4786 29314
rect 6414 29262 6466 29314
rect 9998 29262 10050 29314
rect 24670 29262 24722 29314
rect 38558 29262 38610 29314
rect 41694 29262 41746 29314
rect 43822 29262 43874 29314
rect 11118 29150 11170 29202
rect 15710 29150 15762 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 6750 28814 6802 28866
rect 9438 28814 9490 28866
rect 15486 28814 15538 28866
rect 16606 28814 16658 28866
rect 42478 28814 42530 28866
rect 6638 28702 6690 28754
rect 9326 28702 9378 28754
rect 10334 28702 10386 28754
rect 16718 28702 16770 28754
rect 17166 28702 17218 28754
rect 19406 28702 19458 28754
rect 33070 28702 33122 28754
rect 33630 28702 33682 28754
rect 41918 28702 41970 28754
rect 10110 28590 10162 28642
rect 10782 28590 10834 28642
rect 15262 28590 15314 28642
rect 15486 28590 15538 28642
rect 37326 28590 37378 28642
rect 37550 28590 37602 28642
rect 37774 28590 37826 28642
rect 41470 28590 41522 28642
rect 42142 28590 42194 28642
rect 15822 28478 15874 28530
rect 16270 28478 16322 28530
rect 36990 28478 37042 28530
rect 38110 28478 38162 28530
rect 41694 28478 41746 28530
rect 42366 28478 42418 28530
rect 42478 28478 42530 28530
rect 16158 28366 16210 28418
rect 37102 28366 37154 28418
rect 37998 28366 38050 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 15822 28030 15874 28082
rect 16046 28030 16098 28082
rect 38222 28030 38274 28082
rect 39006 28030 39058 28082
rect 13694 27918 13746 27970
rect 25230 27918 25282 27970
rect 36990 27918 37042 27970
rect 13582 27806 13634 27858
rect 14030 27806 14082 27858
rect 14926 27806 14978 27858
rect 15710 27806 15762 27858
rect 16158 27806 16210 27858
rect 18734 27806 18786 27858
rect 19070 27806 19122 27858
rect 19294 27806 19346 27858
rect 19742 27806 19794 27858
rect 25454 27806 25506 27858
rect 26014 27806 26066 27858
rect 37774 27806 37826 27858
rect 39342 27806 39394 27858
rect 13246 27694 13298 27746
rect 15934 27694 15986 27746
rect 18958 27694 19010 27746
rect 20526 27694 20578 27746
rect 22654 27694 22706 27746
rect 34862 27694 34914 27746
rect 38670 27694 38722 27746
rect 15038 27582 15090 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 30382 27246 30434 27298
rect 30718 27246 30770 27298
rect 13806 27134 13858 27186
rect 15374 27134 15426 27186
rect 19742 27134 19794 27186
rect 21310 27134 21362 27186
rect 31278 27134 31330 27186
rect 12910 27022 12962 27074
rect 13918 27022 13970 27074
rect 14366 27022 14418 27074
rect 21422 27022 21474 27074
rect 21758 27022 21810 27074
rect 31838 27022 31890 27074
rect 35758 27022 35810 27074
rect 13806 26910 13858 26962
rect 25566 26910 25618 26962
rect 25902 26910 25954 26962
rect 30046 26910 30098 26962
rect 30942 26910 30994 26962
rect 31726 26910 31778 26962
rect 36094 26910 36146 26962
rect 7310 26798 7362 26850
rect 12574 26798 12626 26850
rect 14142 26798 14194 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 5182 26462 5234 26514
rect 7086 26462 7138 26514
rect 11006 26462 11058 26514
rect 11790 26462 11842 26514
rect 12126 26462 12178 26514
rect 12350 26462 12402 26514
rect 15374 26462 15426 26514
rect 17390 26462 17442 26514
rect 23214 26462 23266 26514
rect 35646 26462 35698 26514
rect 6974 26350 7026 26402
rect 11230 26350 11282 26402
rect 12014 26350 12066 26402
rect 12686 26350 12738 26402
rect 16830 26350 16882 26402
rect 17950 26350 18002 26402
rect 18734 26350 18786 26402
rect 19630 26350 19682 26402
rect 31614 26350 31666 26402
rect 1822 26238 1874 26290
rect 6526 26238 6578 26290
rect 6750 26238 6802 26290
rect 7758 26238 7810 26290
rect 10670 26238 10722 26290
rect 11566 26238 11618 26290
rect 15486 26238 15538 26290
rect 16270 26238 16322 26290
rect 16606 26238 16658 26290
rect 18958 26238 19010 26290
rect 19294 26238 19346 26290
rect 27022 26238 27074 26290
rect 30046 26238 30098 26290
rect 30494 26238 30546 26290
rect 30718 26238 30770 26290
rect 31278 26238 31330 26290
rect 31950 26238 32002 26290
rect 35422 26238 35474 26290
rect 2606 26126 2658 26178
rect 4734 26126 4786 26178
rect 7310 26126 7362 26178
rect 8206 26126 8258 26178
rect 10894 26126 10946 26178
rect 13134 26126 13186 26178
rect 16494 26126 16546 26178
rect 17502 26126 17554 26178
rect 19070 26126 19122 26178
rect 23774 26126 23826 26178
rect 27694 26126 27746 26178
rect 29822 26126 29874 26178
rect 30270 26126 30322 26178
rect 32398 26126 32450 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 4062 25678 4114 25730
rect 7422 25678 7474 25730
rect 11342 25678 11394 25730
rect 11566 25678 11618 25730
rect 4398 25566 4450 25618
rect 5854 25566 5906 25618
rect 37886 25566 37938 25618
rect 40238 25566 40290 25618
rect 44046 25566 44098 25618
rect 6750 25454 6802 25506
rect 7086 25454 7138 25506
rect 30830 25454 30882 25506
rect 37438 25454 37490 25506
rect 40574 25454 40626 25506
rect 41134 25454 41186 25506
rect 5854 25342 5906 25394
rect 6302 25342 6354 25394
rect 17278 25342 17330 25394
rect 29598 25342 29650 25394
rect 29934 25342 29986 25394
rect 30718 25342 30770 25394
rect 36990 25342 37042 25394
rect 40686 25342 40738 25394
rect 41918 25342 41970 25394
rect 4174 25230 4226 25282
rect 4846 25230 4898 25282
rect 5742 25230 5794 25282
rect 6078 25230 6130 25282
rect 7310 25230 7362 25282
rect 7758 25230 7810 25282
rect 11454 25230 11506 25282
rect 17614 25230 17666 25282
rect 31278 25230 31330 25282
rect 40910 25230 40962 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 8654 24894 8706 24946
rect 25230 24894 25282 24946
rect 29262 24894 29314 24946
rect 35646 24894 35698 24946
rect 36542 24894 36594 24946
rect 41806 24894 41858 24946
rect 5518 24782 5570 24834
rect 6638 24782 6690 24834
rect 8878 24782 8930 24834
rect 28702 24782 28754 24834
rect 29934 24782 29986 24834
rect 31390 24782 31442 24834
rect 35870 24782 35922 24834
rect 35982 24782 36034 24834
rect 36654 24782 36706 24834
rect 39230 24782 39282 24834
rect 40014 24782 40066 24834
rect 6078 24670 6130 24722
rect 6190 24670 6242 24722
rect 6414 24670 6466 24722
rect 8990 24670 9042 24722
rect 15598 24670 15650 24722
rect 16046 24670 16098 24722
rect 28590 24670 28642 24722
rect 28926 24670 28978 24722
rect 29150 24670 29202 24722
rect 29486 24670 29538 24722
rect 31614 24670 31666 24722
rect 36206 24670 36258 24722
rect 39118 24670 39170 24722
rect 39790 24670 39842 24722
rect 41470 24670 41522 24722
rect 41918 24670 41970 24722
rect 42030 24670 42082 24722
rect 6302 24558 6354 24610
rect 16270 24558 16322 24610
rect 25790 24558 25842 24610
rect 38782 24558 38834 24610
rect 5630 24446 5682 24498
rect 36542 24446 36594 24498
rect 39230 24446 39282 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3726 24110 3778 24162
rect 4062 24110 4114 24162
rect 13806 24110 13858 24162
rect 9214 23998 9266 24050
rect 11454 23998 11506 24050
rect 14254 23998 14306 24050
rect 16270 23998 16322 24050
rect 21422 23998 21474 24050
rect 38670 23998 38722 24050
rect 41806 23998 41858 24050
rect 9102 23886 9154 23938
rect 9438 23886 9490 23938
rect 10782 23886 10834 23938
rect 11230 23886 11282 23938
rect 16718 23886 16770 23938
rect 16942 23886 16994 23938
rect 17166 23886 17218 23938
rect 17278 23886 17330 23938
rect 20750 23886 20802 23938
rect 24222 23886 24274 23938
rect 38894 23886 38946 23938
rect 42030 23886 42082 23938
rect 42366 23886 42418 23938
rect 13582 23774 13634 23826
rect 20414 23774 20466 23826
rect 23550 23774 23602 23826
rect 39678 23774 39730 23826
rect 3838 23662 3890 23714
rect 8878 23662 8930 23714
rect 13694 23662 13746 23714
rect 17726 23662 17778 23714
rect 24782 23662 24834 23714
rect 42254 23662 42306 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 8206 23326 8258 23378
rect 11230 23326 11282 23378
rect 11454 23326 11506 23378
rect 12014 23326 12066 23378
rect 12350 23326 12402 23378
rect 17390 23326 17442 23378
rect 39566 23326 39618 23378
rect 6302 23214 6354 23266
rect 17502 23214 17554 23266
rect 35310 23214 35362 23266
rect 36094 23214 36146 23266
rect 36206 23214 36258 23266
rect 39902 23214 39954 23266
rect 5854 23102 5906 23154
rect 6190 23102 6242 23154
rect 7982 23102 8034 23154
rect 10222 23102 10274 23154
rect 11118 23102 11170 23154
rect 11566 23102 11618 23154
rect 17726 23102 17778 23154
rect 17950 23102 18002 23154
rect 19182 23102 19234 23154
rect 28254 23102 28306 23154
rect 28478 23102 28530 23154
rect 31390 23102 31442 23154
rect 35646 23102 35698 23154
rect 36430 23102 36482 23154
rect 39230 23102 39282 23154
rect 39678 23102 39730 23154
rect 9886 22990 9938 23042
rect 11342 22990 11394 23042
rect 18846 22990 18898 23042
rect 27582 22990 27634 23042
rect 30830 22990 30882 23042
rect 31726 22990 31778 23042
rect 32286 22990 32338 23042
rect 36094 22990 36146 23042
rect 10222 22878 10274 22930
rect 19294 22878 19346 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 21758 22542 21810 22594
rect 4174 22430 4226 22482
rect 5742 22430 5794 22482
rect 8430 22430 8482 22482
rect 19854 22430 19906 22482
rect 21422 22430 21474 22482
rect 26686 22430 26738 22482
rect 36430 22430 36482 22482
rect 3838 22318 3890 22370
rect 5630 22318 5682 22370
rect 6078 22318 6130 22370
rect 9774 22318 9826 22370
rect 11230 22318 11282 22370
rect 17950 22318 18002 22370
rect 18286 22318 18338 22370
rect 18622 22318 18674 22370
rect 19294 22318 19346 22370
rect 19742 22318 19794 22370
rect 22206 22318 22258 22370
rect 33630 22318 33682 22370
rect 37102 22318 37154 22370
rect 6302 22206 6354 22258
rect 9886 22206 9938 22258
rect 10894 22206 10946 22258
rect 18398 22206 18450 22258
rect 34302 22206 34354 22258
rect 4062 22094 4114 22146
rect 5854 22094 5906 22146
rect 17614 22094 17666 22146
rect 19518 22094 19570 22146
rect 19854 22094 19906 22146
rect 21646 22094 21698 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 4846 21758 4898 21810
rect 15486 21758 15538 21810
rect 21982 21758 22034 21810
rect 35310 21758 35362 21810
rect 2606 21646 2658 21698
rect 15934 21646 15986 21698
rect 35422 21646 35474 21698
rect 1934 21534 1986 21586
rect 15262 21534 15314 21586
rect 15710 21534 15762 21586
rect 25454 21534 25506 21586
rect 29598 21534 29650 21586
rect 5518 21422 5570 21474
rect 15598 21422 15650 21474
rect 26126 21422 26178 21474
rect 28254 21422 28306 21474
rect 28702 21422 28754 21474
rect 30270 21422 30322 21474
rect 32398 21422 32450 21474
rect 33182 21422 33234 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 10894 20974 10946 21026
rect 14702 20974 14754 21026
rect 27022 20974 27074 21026
rect 27358 20974 27410 21026
rect 30494 20974 30546 21026
rect 41806 20974 41858 21026
rect 10558 20862 10610 20914
rect 14366 20862 14418 20914
rect 19630 20862 19682 20914
rect 23774 20862 23826 20914
rect 24110 20862 24162 20914
rect 30270 20862 30322 20914
rect 36206 20862 36258 20914
rect 36318 20862 36370 20914
rect 18846 20750 18898 20802
rect 26686 20750 26738 20802
rect 27022 20750 27074 20802
rect 29822 20750 29874 20802
rect 30158 20750 30210 20802
rect 32398 20750 32450 20802
rect 35982 20750 36034 20802
rect 41918 20750 41970 20802
rect 19182 20638 19234 20690
rect 24446 20638 24498 20690
rect 32174 20638 32226 20690
rect 10670 20526 10722 20578
rect 13582 20526 13634 20578
rect 14478 20526 14530 20578
rect 24782 20526 24834 20578
rect 25118 20526 25170 20578
rect 25454 20526 25506 20578
rect 31950 20526 32002 20578
rect 41806 20526 41858 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 19630 20190 19682 20242
rect 23998 20190 24050 20242
rect 24558 20190 24610 20242
rect 10558 20078 10610 20130
rect 14366 20078 14418 20130
rect 18846 20078 18898 20130
rect 19182 20078 19234 20130
rect 23662 20078 23714 20130
rect 39118 20078 39170 20130
rect 39454 20078 39506 20130
rect 39790 20078 39842 20130
rect 9886 19966 9938 20018
rect 13694 19966 13746 20018
rect 17614 19966 17666 20018
rect 17950 19966 18002 20018
rect 18286 19966 18338 20018
rect 19406 19966 19458 20018
rect 19742 19966 19794 20018
rect 20974 19966 21026 20018
rect 41134 19966 41186 20018
rect 12686 19854 12738 19906
rect 16494 19854 16546 19906
rect 19630 19854 19682 19906
rect 20638 19854 20690 19906
rect 40350 19854 40402 19906
rect 41918 19854 41970 19906
rect 44046 19854 44098 19906
rect 20974 19742 21026 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 6078 19294 6130 19346
rect 6414 19294 6466 19346
rect 18958 19294 19010 19346
rect 41806 19294 41858 19346
rect 11230 19182 11282 19234
rect 36206 19182 36258 19234
rect 42478 19182 42530 19234
rect 6190 19070 6242 19122
rect 11454 19070 11506 19122
rect 13806 19070 13858 19122
rect 38894 19070 38946 19122
rect 39230 19070 39282 19122
rect 39566 19070 39618 19122
rect 41358 19070 41410 19122
rect 41582 19070 41634 19122
rect 41918 19070 41970 19122
rect 42142 19070 42194 19122
rect 42366 19070 42418 19122
rect 6862 18958 6914 19010
rect 14142 18958 14194 19010
rect 14590 18958 14642 19010
rect 35646 18958 35698 19010
rect 35870 18958 35922 19010
rect 36094 18958 36146 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 5630 18622 5682 18674
rect 6974 18622 7026 18674
rect 20190 18622 20242 18674
rect 34862 18622 34914 18674
rect 35198 18622 35250 18674
rect 41246 18622 41298 18674
rect 9550 18510 9602 18562
rect 14814 18510 14866 18562
rect 40910 18510 40962 18562
rect 41022 18510 41074 18562
rect 41582 18510 41634 18562
rect 41694 18510 41746 18562
rect 4958 18398 5010 18450
rect 5854 18398 5906 18450
rect 6190 18398 6242 18450
rect 6526 18398 6578 18450
rect 6750 18398 6802 18450
rect 6862 18398 6914 18450
rect 7198 18398 7250 18450
rect 7534 18398 7586 18450
rect 9886 18398 9938 18450
rect 11678 18398 11730 18450
rect 11902 18398 11954 18450
rect 12350 18398 12402 18450
rect 14590 18398 14642 18450
rect 22430 18398 22482 18450
rect 23214 18398 23266 18450
rect 29822 18398 29874 18450
rect 35310 18398 35362 18450
rect 35646 18398 35698 18450
rect 36094 18398 36146 18450
rect 37214 18398 37266 18450
rect 5742 18286 5794 18338
rect 23662 18286 23714 18338
rect 30046 18286 30098 18338
rect 36430 18286 36482 18338
rect 4958 18174 5010 18226
rect 5294 18174 5346 18226
rect 7758 18174 7810 18226
rect 7982 18174 8034 18226
rect 8094 18174 8146 18226
rect 11342 18174 11394 18226
rect 30158 18174 30210 18226
rect 35198 18174 35250 18226
rect 41582 18174 41634 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 2606 17726 2658 17778
rect 4734 17726 4786 17778
rect 19182 17726 19234 17778
rect 27358 17726 27410 17778
rect 33182 17726 33234 17778
rect 34862 17726 34914 17778
rect 35198 17726 35250 17778
rect 36430 17726 36482 17778
rect 1934 17614 1986 17666
rect 5742 17614 5794 17666
rect 6414 17614 6466 17666
rect 6974 17614 7026 17666
rect 7310 17614 7362 17666
rect 18062 17614 18114 17666
rect 18622 17614 18674 17666
rect 23774 17614 23826 17666
rect 24558 17614 24610 17666
rect 30158 17614 30210 17666
rect 35310 17614 35362 17666
rect 35534 17614 35586 17666
rect 40350 17614 40402 17666
rect 41582 17614 41634 17666
rect 5966 17502 6018 17554
rect 6526 17502 6578 17554
rect 18174 17502 18226 17554
rect 18286 17502 18338 17554
rect 23998 17502 24050 17554
rect 24110 17502 24162 17554
rect 25230 17502 25282 17554
rect 35758 17502 35810 17554
rect 35982 17502 36034 17554
rect 36990 17502 37042 17554
rect 37326 17502 37378 17554
rect 37438 17502 37490 17554
rect 40910 17502 40962 17554
rect 41134 17502 41186 17554
rect 6750 17390 6802 17442
rect 7086 17390 7138 17442
rect 17950 17390 18002 17442
rect 27806 17390 27858 17442
rect 28590 17390 28642 17442
rect 34750 17390 34802 17442
rect 37102 17390 37154 17442
rect 37214 17390 37266 17442
rect 40462 17390 40514 17442
rect 40686 17390 40738 17442
rect 41246 17390 41298 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 4958 17054 5010 17106
rect 17950 17054 18002 17106
rect 20638 17054 20690 17106
rect 13582 16942 13634 16994
rect 17502 16942 17554 16994
rect 22542 16942 22594 16994
rect 27694 16942 27746 16994
rect 31278 16942 31330 16994
rect 32510 16942 32562 16994
rect 36766 16942 36818 16994
rect 11678 16830 11730 16882
rect 16606 16830 16658 16882
rect 17838 16830 17890 16882
rect 19742 16830 19794 16882
rect 20974 16830 21026 16882
rect 22318 16830 22370 16882
rect 22990 16830 23042 16882
rect 28366 16830 28418 16882
rect 32062 16830 32114 16882
rect 33294 16830 33346 16882
rect 20078 16718 20130 16770
rect 28590 16718 28642 16770
rect 29150 16718 29202 16770
rect 17390 16606 17442 16658
rect 17950 16606 18002 16658
rect 19742 16606 19794 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 24782 16270 24834 16322
rect 9102 16158 9154 16210
rect 12350 16158 12402 16210
rect 18510 16158 18562 16210
rect 21422 16158 21474 16210
rect 34302 16158 34354 16210
rect 36430 16158 36482 16210
rect 37102 16158 37154 16210
rect 41246 16158 41298 16210
rect 43374 16158 43426 16210
rect 7422 16046 7474 16098
rect 7758 16046 7810 16098
rect 7870 16046 7922 16098
rect 8206 16046 8258 16098
rect 10782 16046 10834 16098
rect 12686 16046 12738 16098
rect 13022 16046 13074 16098
rect 15486 16046 15538 16098
rect 25566 16046 25618 16098
rect 26910 16046 26962 16098
rect 29150 16046 29202 16098
rect 32958 16046 33010 16098
rect 33630 16046 33682 16098
rect 40462 16046 40514 16098
rect 8542 15934 8594 15986
rect 8654 15934 8706 15986
rect 25230 15934 25282 15986
rect 25342 15934 25394 15986
rect 26126 15934 26178 15986
rect 26798 15934 26850 15986
rect 29262 15934 29314 15986
rect 32286 15934 32338 15986
rect 7534 15822 7586 15874
rect 10446 15822 10498 15874
rect 12798 15822 12850 15874
rect 26574 15822 26626 15874
rect 29374 15822 29426 15874
rect 40126 15822 40178 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 8878 15486 8930 15538
rect 9662 15486 9714 15538
rect 14366 15486 14418 15538
rect 21870 15486 21922 15538
rect 30270 15486 30322 15538
rect 30606 15486 30658 15538
rect 33294 15486 33346 15538
rect 2718 15374 2770 15426
rect 5742 15374 5794 15426
rect 7758 15374 7810 15426
rect 9886 15374 9938 15426
rect 14030 15374 14082 15426
rect 30158 15374 30210 15426
rect 37438 15374 37490 15426
rect 1934 15262 1986 15314
rect 6862 15262 6914 15314
rect 7310 15262 7362 15314
rect 9550 15262 9602 15314
rect 9998 15262 10050 15314
rect 13694 15262 13746 15314
rect 30382 15262 30434 15314
rect 4846 15150 4898 15202
rect 13134 15150 13186 15202
rect 14814 15150 14866 15202
rect 21758 15150 21810 15202
rect 29598 15150 29650 15202
rect 29822 15150 29874 15202
rect 22094 15038 22146 15090
rect 29262 15038 29314 15090
rect 37550 15038 37602 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 9998 14702 10050 14754
rect 29486 14702 29538 14754
rect 29934 14702 29986 14754
rect 15934 14590 15986 14642
rect 18062 14590 18114 14642
rect 18510 14590 18562 14642
rect 25790 14590 25842 14642
rect 29934 14590 29986 14642
rect 38110 14590 38162 14642
rect 40238 14590 40290 14642
rect 9998 14478 10050 14530
rect 15262 14478 15314 14530
rect 37326 14478 37378 14530
rect 9662 14366 9714 14418
rect 5070 14254 5122 14306
rect 13470 14254 13522 14306
rect 13806 14254 13858 14306
rect 14254 14254 14306 14306
rect 36430 14254 36482 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 7758 13918 7810 13970
rect 8094 13918 8146 13970
rect 19518 13918 19570 13970
rect 34414 13918 34466 13970
rect 20638 13806 20690 13858
rect 26126 13806 26178 13858
rect 19854 13694 19906 13746
rect 24670 13694 24722 13746
rect 26350 13694 26402 13746
rect 22766 13582 22818 13634
rect 24334 13582 24386 13634
rect 24670 13470 24722 13522
rect 25230 13470 25282 13522
rect 25342 13470 25394 13522
rect 25566 13470 25618 13522
rect 25678 13470 25730 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 29486 13134 29538 13186
rect 22878 13022 22930 13074
rect 25006 13022 25058 13074
rect 35198 13022 35250 13074
rect 7758 12910 7810 12962
rect 7982 12910 8034 12962
rect 8094 12910 8146 12962
rect 25790 12910 25842 12962
rect 29710 12910 29762 12962
rect 29934 12910 29986 12962
rect 30382 12910 30434 12962
rect 30830 12910 30882 12962
rect 33294 12910 33346 12962
rect 33966 12910 34018 12962
rect 34750 12910 34802 12962
rect 29374 12798 29426 12850
rect 30270 12798 30322 12850
rect 30606 12798 30658 12850
rect 32846 12798 32898 12850
rect 33182 12798 33234 12850
rect 8542 12686 8594 12738
rect 26238 12686 26290 12738
rect 33070 12686 33122 12738
rect 33742 12686 33794 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 6302 12350 6354 12402
rect 9662 12350 9714 12402
rect 16046 12350 16098 12402
rect 16830 12350 16882 12402
rect 2606 12238 2658 12290
rect 7646 12238 7698 12290
rect 8766 12238 8818 12290
rect 12238 12238 12290 12290
rect 12798 12238 12850 12290
rect 28814 12238 28866 12290
rect 35198 12238 35250 12290
rect 1934 12126 1986 12178
rect 6078 12126 6130 12178
rect 7534 12126 7586 12178
rect 7870 12126 7922 12178
rect 8318 12126 8370 12178
rect 8654 12126 8706 12178
rect 11566 12126 11618 12178
rect 11902 12126 11954 12178
rect 15934 12126 15986 12178
rect 20526 12126 20578 12178
rect 25230 12126 25282 12178
rect 25454 12126 25506 12178
rect 28142 12126 28194 12178
rect 31390 12126 31442 12178
rect 35870 12126 35922 12178
rect 4734 12014 4786 12066
rect 5182 12014 5234 12066
rect 11790 12014 11842 12066
rect 14814 12014 14866 12066
rect 17726 12014 17778 12066
rect 19854 12014 19906 12066
rect 30942 12014 30994 12066
rect 33070 12014 33122 12066
rect 36430 12014 36482 12066
rect 8094 11902 8146 11954
rect 15038 11902 15090 11954
rect 15262 11902 15314 11954
rect 15710 11902 15762 11954
rect 16046 11902 16098 11954
rect 25790 11902 25842 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 13806 11566 13858 11618
rect 29934 11566 29986 11618
rect 8430 11454 8482 11506
rect 9326 11454 9378 11506
rect 17838 11454 17890 11506
rect 17950 11454 18002 11506
rect 32958 11454 33010 11506
rect 6638 11342 6690 11394
rect 6974 11342 7026 11394
rect 7422 11342 7474 11394
rect 7870 11342 7922 11394
rect 8878 11342 8930 11394
rect 12238 11342 12290 11394
rect 16830 11342 16882 11394
rect 17054 11342 17106 11394
rect 17390 11342 17442 11394
rect 17614 11342 17666 11394
rect 18062 11342 18114 11394
rect 18286 11342 18338 11394
rect 30718 11342 30770 11394
rect 32510 11342 32562 11394
rect 32846 11342 32898 11394
rect 33518 11342 33570 11394
rect 7198 11230 7250 11282
rect 8430 11230 8482 11282
rect 12350 11230 12402 11282
rect 13694 11230 13746 11282
rect 16718 11230 16770 11282
rect 18622 11230 18674 11282
rect 30382 11230 30434 11282
rect 30494 11230 30546 11282
rect 33070 11230 33122 11282
rect 6750 11118 6802 11170
rect 7534 11118 7586 11170
rect 7646 11118 7698 11170
rect 8318 11118 8370 11170
rect 8654 11118 8706 11170
rect 12574 11118 12626 11170
rect 13806 11118 13858 11170
rect 18846 11118 18898 11170
rect 18958 11118 19010 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 8318 10782 8370 10834
rect 8542 10782 8594 10834
rect 8654 10782 8706 10834
rect 9102 10782 9154 10834
rect 10222 10670 10274 10722
rect 11790 10670 11842 10722
rect 15150 10670 15202 10722
rect 15934 10670 15986 10722
rect 30382 10670 30434 10722
rect 7198 10558 7250 10610
rect 7422 10558 7474 10610
rect 7870 10558 7922 10610
rect 8094 10558 8146 10610
rect 10446 10558 10498 10610
rect 11230 10558 11282 10610
rect 11342 10558 11394 10610
rect 11566 10558 11618 10610
rect 12574 10558 12626 10610
rect 12686 10558 12738 10610
rect 13806 10558 13858 10610
rect 14366 10558 14418 10610
rect 15262 10558 15314 10610
rect 15710 10558 15762 10610
rect 16382 10558 16434 10610
rect 30046 10558 30098 10610
rect 7310 10446 7362 10498
rect 11454 10446 11506 10498
rect 15822 10446 15874 10498
rect 10782 10334 10834 10386
rect 12910 10334 12962 10386
rect 13022 10334 13074 10386
rect 15374 10334 15426 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 6750 9998 6802 10050
rect 29598 9998 29650 10050
rect 29822 9998 29874 10050
rect 16270 9886 16322 9938
rect 23550 9886 23602 9938
rect 24110 9886 24162 9938
rect 7310 9774 7362 9826
rect 12126 9774 12178 9826
rect 12462 9774 12514 9826
rect 12798 9774 12850 9826
rect 13694 9774 13746 9826
rect 14478 9774 14530 9826
rect 16606 9774 16658 9826
rect 19070 9774 19122 9826
rect 19182 9774 19234 9826
rect 19406 9774 19458 9826
rect 29374 9774 29426 9826
rect 6526 9662 6578 9714
rect 7086 9662 7138 9714
rect 13470 9662 13522 9714
rect 14590 9662 14642 9714
rect 18174 9662 18226 9714
rect 23214 9662 23266 9714
rect 29934 9662 29986 9714
rect 6638 9550 6690 9602
rect 7982 9550 8034 9602
rect 12350 9550 12402 9602
rect 18622 9550 18674 9602
rect 19854 9550 19906 9602
rect 23438 9550 23490 9602
rect 23662 9550 23714 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 14254 9214 14306 9266
rect 16382 9214 16434 9266
rect 21422 9214 21474 9266
rect 27470 9214 27522 9266
rect 28926 9214 28978 9266
rect 4510 9102 4562 9154
rect 16494 9102 16546 9154
rect 25342 9102 25394 9154
rect 27582 9102 27634 9154
rect 28366 9102 28418 9154
rect 3838 8990 3890 9042
rect 7086 8990 7138 9042
rect 14590 8990 14642 9042
rect 21870 8990 21922 9042
rect 25678 8990 25730 9042
rect 27134 8990 27186 9042
rect 27806 8990 27858 9042
rect 28254 8990 28306 9042
rect 28478 8990 28530 9042
rect 6638 8878 6690 8930
rect 22542 8878 22594 8930
rect 24670 8878 24722 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 12350 8430 12402 8482
rect 10782 8318 10834 8370
rect 11118 8318 11170 8370
rect 11566 8318 11618 8370
rect 12686 8318 12738 8370
rect 23102 8318 23154 8370
rect 29486 8318 29538 8370
rect 31614 8318 31666 8370
rect 18286 8206 18338 8258
rect 22654 8206 22706 8258
rect 22990 8206 23042 8258
rect 23326 8206 23378 8258
rect 23550 8206 23602 8258
rect 27806 8206 27858 8258
rect 32398 8206 32450 8258
rect 32958 8206 33010 8258
rect 10894 8094 10946 8146
rect 12574 8094 12626 8146
rect 27582 8094 27634 8146
rect 13582 7982 13634 8034
rect 18510 7982 18562 8034
rect 22430 7982 22482 8034
rect 22542 7982 22594 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 22990 7646 23042 7698
rect 27582 7646 27634 7698
rect 19518 7534 19570 7586
rect 26686 7534 26738 7586
rect 28702 7534 28754 7586
rect 20302 7422 20354 7474
rect 27694 7422 27746 7474
rect 28254 7422 28306 7474
rect 17390 7310 17442 7362
rect 20750 7310 20802 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 26798 6862 26850 6914
rect 10670 6750 10722 6802
rect 12798 6750 12850 6802
rect 9998 6638 10050 6690
rect 13582 6638 13634 6690
rect 25902 6638 25954 6690
rect 26798 6638 26850 6690
rect 27470 6638 27522 6690
rect 26238 6526 26290 6578
rect 26350 6526 26402 6578
rect 27134 6526 27186 6578
rect 27806 6526 27858 6578
rect 26574 6414 26626 6466
rect 27582 6414 27634 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 15374 6078 15426 6130
rect 25902 6078 25954 6130
rect 12798 5966 12850 6018
rect 26462 5966 26514 6018
rect 27134 5966 27186 6018
rect 27358 5966 27410 6018
rect 28030 5966 28082 6018
rect 12126 5854 12178 5906
rect 23102 5854 23154 5906
rect 25678 5854 25730 5906
rect 26014 5854 26066 5906
rect 14926 5742 14978 5794
rect 23326 5742 23378 5794
rect 27470 5742 27522 5794
rect 22766 5630 22818 5682
rect 26350 5630 26402 5682
rect 27806 5630 27858 5682
rect 28142 5630 28194 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 24558 5182 24610 5234
rect 20862 5070 20914 5122
rect 21646 5070 21698 5122
rect 22430 4958 22482 5010
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 22430 4510 22482 4562
rect 30270 4510 30322 4562
rect 22766 4398 22818 4450
rect 27694 4398 27746 4450
rect 27022 4286 27074 4338
rect 29822 4174 29874 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 1792 45200 1904 46000
rect 5600 45200 5712 46000
rect 9408 45200 9520 46000
rect 13216 45200 13328 46000
rect 17024 45200 17136 46000
rect 17388 45276 17892 45332
rect 1820 43708 1876 45200
rect 1708 43652 1876 43708
rect 5628 43708 5684 45200
rect 9436 43708 9492 45200
rect 5628 43652 5908 43708
rect 9436 43652 9716 43708
rect 1708 22372 1764 43652
rect 5068 41972 5124 41982
rect 5852 41972 5908 43652
rect 5068 41970 5908 41972
rect 5068 41918 5070 41970
rect 5122 41918 5854 41970
rect 5906 41918 5908 41970
rect 5068 41916 5908 41918
rect 5068 41906 5124 41916
rect 5852 41906 5908 41916
rect 6188 42082 6244 42094
rect 6188 42030 6190 42082
rect 6242 42030 6244 42082
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 5628 40516 5684 40526
rect 5628 40422 5684 40460
rect 4956 40404 5012 40414
rect 4956 40310 5012 40348
rect 5740 40404 5796 40414
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4732 39732 4788 39742
rect 4732 39638 4788 39676
rect 5740 39730 5796 40348
rect 5740 39678 5742 39730
rect 5794 39678 5796 39730
rect 1820 39618 1876 39630
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1820 38164 1876 39566
rect 2604 39506 2660 39518
rect 2604 39454 2606 39506
rect 2658 39454 2660 39506
rect 1820 38098 1876 38108
rect 2268 38164 2324 38174
rect 2268 38050 2324 38108
rect 2268 37998 2270 38050
rect 2322 37998 2324 38050
rect 2268 34914 2324 37998
rect 2604 37492 2660 39454
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 5068 38164 5124 38174
rect 5740 38164 5796 39678
rect 5068 38162 5348 38164
rect 5068 38110 5070 38162
rect 5122 38110 5348 38162
rect 5068 38108 5348 38110
rect 5068 38098 5124 38108
rect 2940 37940 2996 37950
rect 2940 37846 2996 37884
rect 5068 37940 5124 37950
rect 2604 37426 2660 37436
rect 4620 37492 4676 37502
rect 4620 37398 4676 37436
rect 5068 37490 5124 37884
rect 5068 37438 5070 37490
rect 5122 37438 5124 37490
rect 5068 37426 5124 37438
rect 4396 37268 4452 37278
rect 2268 34862 2270 34914
rect 2322 34862 2324 34914
rect 2268 32562 2324 34862
rect 4284 37212 4396 37268
rect 2940 34802 2996 34814
rect 2940 34750 2942 34802
rect 2994 34750 2996 34802
rect 2940 33908 2996 34750
rect 2940 33842 2996 33852
rect 2268 32510 2270 32562
rect 2322 32510 2324 32562
rect 2268 31948 2324 32510
rect 3052 32452 3108 32462
rect 3052 32358 3108 32396
rect 4284 31948 4340 37212
rect 4396 37174 4452 37212
rect 5180 37154 5236 37166
rect 5180 37102 5182 37154
rect 5234 37102 5236 37154
rect 4732 37044 4788 37054
rect 4732 37042 4900 37044
rect 4732 36990 4734 37042
rect 4786 36990 4900 37042
rect 4732 36988 4900 36990
rect 4732 36978 4788 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 36708 4900 36988
rect 4844 36642 4900 36652
rect 5180 35364 5236 37102
rect 5292 35476 5348 38108
rect 5628 37268 5684 37278
rect 5628 37174 5684 37212
rect 5292 35410 5348 35420
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 5180 35298 5236 35308
rect 4476 35242 4740 35252
rect 5068 35026 5124 35038
rect 5068 34974 5070 35026
rect 5122 34974 5124 35026
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 5068 33012 5124 34974
rect 5740 35026 5796 38108
rect 6188 36484 6244 42030
rect 8876 41972 8932 41982
rect 9660 41972 9716 43652
rect 8876 41970 9716 41972
rect 8876 41918 8878 41970
rect 8930 41918 9662 41970
rect 9714 41918 9716 41970
rect 8876 41916 9716 41918
rect 8876 41906 8932 41916
rect 9660 41906 9716 41916
rect 9996 42082 10052 42094
rect 9996 42030 9998 42082
rect 10050 42030 10052 42082
rect 8764 40516 8820 40526
rect 8764 40422 8820 40460
rect 8316 40404 8372 40414
rect 8316 40310 8372 40348
rect 9772 40404 9828 40414
rect 9996 40404 10052 42030
rect 12684 41972 12740 41982
rect 10444 40404 10500 40414
rect 9996 40348 10276 40404
rect 9772 40310 9828 40348
rect 7756 40290 7812 40302
rect 7756 40238 7758 40290
rect 7810 40238 7812 40290
rect 6188 36418 6244 36428
rect 6972 39732 7028 39742
rect 6972 36594 7028 39676
rect 7756 39732 7812 40238
rect 7756 39666 7812 39676
rect 8764 39732 8820 39742
rect 8764 39638 8820 39676
rect 8876 39394 8932 39406
rect 8876 39342 8878 39394
rect 8930 39342 8932 39394
rect 7756 38162 7812 38174
rect 7756 38110 7758 38162
rect 7810 38110 7812 38162
rect 7420 36708 7476 36718
rect 7420 36614 7476 36652
rect 7756 36708 7812 38110
rect 7756 36642 7812 36652
rect 6972 36542 6974 36594
rect 7026 36542 7028 36594
rect 6972 36372 7028 36542
rect 6972 36306 7028 36316
rect 7756 36482 7812 36494
rect 7756 36430 7758 36482
rect 7810 36430 7812 36482
rect 6972 35476 7028 35486
rect 6972 35028 7028 35420
rect 5740 34974 5742 35026
rect 5794 34974 5796 35026
rect 5740 33572 5796 34974
rect 5068 32946 5124 32956
rect 5628 33516 5740 33572
rect 5628 32788 5684 33516
rect 5740 33506 5796 33516
rect 6748 35026 7364 35028
rect 6748 34974 6974 35026
rect 7026 34974 7364 35026
rect 6748 34972 7364 34974
rect 5068 32786 5684 32788
rect 5068 32734 5630 32786
rect 5682 32734 5684 32786
rect 5068 32732 5684 32734
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 1820 31892 2324 31948
rect 4172 31892 4340 31948
rect 1820 29426 1876 31892
rect 1820 29374 1822 29426
rect 1874 29374 1876 29426
rect 1820 26290 1876 29374
rect 2604 29314 2660 29326
rect 2604 29262 2606 29314
rect 2658 29262 2660 29314
rect 2604 26964 2660 29262
rect 2604 26898 2660 26908
rect 3724 26964 3780 26974
rect 1820 26238 1822 26290
rect 1874 26238 1876 26290
rect 1820 26226 1876 26238
rect 2604 26180 2660 26190
rect 2604 26086 2660 26124
rect 3724 24162 3780 26908
rect 4060 26180 4116 26190
rect 4060 25730 4116 26124
rect 4060 25678 4062 25730
rect 4114 25678 4116 25730
rect 4060 25666 4116 25678
rect 4172 25284 4228 31892
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5068 29652 5124 32732
rect 5628 32722 5684 32732
rect 6636 33124 6692 33134
rect 6636 32786 6692 33068
rect 6636 32734 6638 32786
rect 6690 32734 6692 32786
rect 6636 32722 6692 32734
rect 6748 32564 6804 34972
rect 6972 34962 7028 34972
rect 7308 34914 7364 34972
rect 7308 34862 7310 34914
rect 7362 34862 7364 34914
rect 7308 34850 7364 34862
rect 7644 34914 7700 34926
rect 7644 34862 7646 34914
rect 7698 34862 7700 34914
rect 7644 34356 7700 34862
rect 7756 34916 7812 36430
rect 7980 36372 8036 36382
rect 7980 36278 8036 36316
rect 8540 36372 8596 36382
rect 8540 36370 8708 36372
rect 8540 36318 8542 36370
rect 8594 36318 8708 36370
rect 8540 36316 8708 36318
rect 8540 36306 8596 36316
rect 7756 34850 7812 34860
rect 8428 35588 8484 35598
rect 8428 34914 8484 35532
rect 8540 35364 8596 35374
rect 8540 35026 8596 35308
rect 8540 34974 8542 35026
rect 8594 34974 8596 35026
rect 8540 34962 8596 34974
rect 8428 34862 8430 34914
rect 8482 34862 8484 34914
rect 6972 33908 7028 33918
rect 6972 33458 7028 33852
rect 6972 33406 6974 33458
rect 7026 33406 7028 33458
rect 6972 33394 7028 33406
rect 7308 33348 7364 33358
rect 7308 33234 7364 33292
rect 7308 33182 7310 33234
rect 7362 33182 7364 33234
rect 6636 32508 6804 32564
rect 6860 32674 6916 32686
rect 6860 32622 6862 32674
rect 6914 32622 6916 32674
rect 5180 32450 5236 32462
rect 5180 32398 5182 32450
rect 5234 32398 5236 32450
rect 5180 31668 5236 32398
rect 6636 32116 6692 32508
rect 6748 32116 6804 32126
rect 6636 32060 6748 32116
rect 6188 31892 6244 31902
rect 6188 31798 6244 31836
rect 6076 31668 6132 31678
rect 5180 31666 6132 31668
rect 5180 31614 6078 31666
rect 6130 31614 6132 31666
rect 5180 31612 6132 31614
rect 5852 30322 5908 30334
rect 5852 30270 5854 30322
rect 5906 30270 5908 30322
rect 5180 29652 5236 29662
rect 5068 29650 5236 29652
rect 5068 29598 5182 29650
rect 5234 29598 5236 29650
rect 5068 29596 5236 29598
rect 4732 29428 4788 29438
rect 4732 29314 4788 29372
rect 4732 29262 4734 29314
rect 4786 29262 4788 29314
rect 4732 29250 4788 29262
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 5180 26514 5236 29596
rect 5852 26908 5908 30270
rect 6076 30210 6132 31612
rect 6636 31220 6692 32060
rect 6748 32050 6804 32060
rect 6860 31892 6916 32622
rect 7084 32562 7140 32574
rect 7084 32510 7086 32562
rect 7138 32510 7140 32562
rect 6972 32452 7028 32462
rect 6972 32358 7028 32396
rect 7084 31948 7140 32510
rect 7308 32562 7364 33182
rect 7308 32510 7310 32562
rect 7362 32510 7364 32562
rect 7308 32498 7364 32510
rect 7420 33234 7476 33246
rect 7420 33182 7422 33234
rect 7474 33182 7476 33234
rect 7084 31892 7252 31948
rect 6860 31826 6916 31836
rect 6636 31218 7028 31220
rect 6636 31166 6638 31218
rect 6690 31166 7028 31218
rect 6636 31164 7028 31166
rect 6636 31154 6692 31164
rect 6860 30660 6916 30670
rect 6076 30158 6078 30210
rect 6130 30158 6132 30210
rect 6076 30146 6132 30158
rect 6636 30212 6692 30222
rect 6636 30118 6692 30156
rect 5964 29428 6020 29438
rect 5964 29334 6020 29372
rect 6636 29428 6692 29438
rect 6412 29316 6468 29326
rect 6188 29260 6412 29316
rect 5852 26852 6020 26908
rect 5180 26462 5182 26514
rect 5234 26462 5236 26514
rect 5180 26450 5236 26462
rect 4732 26180 4788 26190
rect 4732 26086 4788 26124
rect 5964 26180 6020 26852
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4396 25620 4452 25630
rect 4396 25526 4452 25564
rect 5852 25620 5908 25630
rect 5852 25526 5908 25564
rect 5852 25396 5908 25406
rect 5964 25396 6020 26124
rect 5852 25394 6020 25396
rect 5852 25342 5854 25394
rect 5906 25342 6020 25394
rect 5852 25340 6020 25342
rect 4844 25284 4900 25294
rect 4172 25282 5012 25284
rect 4172 25230 4174 25282
rect 4226 25230 4846 25282
rect 4898 25230 5012 25282
rect 4172 25228 5012 25230
rect 4172 25218 4228 25228
rect 4844 25218 4900 25228
rect 3724 24110 3726 24162
rect 3778 24110 3780 24162
rect 3724 24098 3780 24110
rect 4060 24612 4116 24622
rect 4060 24162 4116 24556
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4060 24110 4062 24162
rect 4114 24110 4116 24162
rect 4060 24098 4116 24110
rect 1708 22306 1764 22316
rect 3836 23714 3892 23726
rect 3836 23662 3838 23714
rect 3890 23662 3892 23714
rect 3836 22370 3892 23662
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 22484 4228 22494
rect 4172 22390 4228 22428
rect 3836 22318 3838 22370
rect 3890 22318 3892 22370
rect 2604 22148 2660 22158
rect 2604 21698 2660 22092
rect 2604 21646 2606 21698
rect 2658 21646 2660 21698
rect 2604 21634 2660 21646
rect 1932 21586 1988 21598
rect 1932 21534 1934 21586
rect 1986 21534 1988 21586
rect 1932 20020 1988 21534
rect 3836 20580 3892 22318
rect 4060 22148 4116 22158
rect 4060 22054 4116 22092
rect 4844 22148 4900 22158
rect 4844 21810 4900 22092
rect 4844 21758 4846 21810
rect 4898 21758 4900 21810
rect 4844 21746 4900 21758
rect 4956 21588 5012 25228
rect 5740 25282 5796 25294
rect 5740 25230 5742 25282
rect 5794 25230 5796 25282
rect 5740 25172 5796 25230
rect 5404 25116 5796 25172
rect 5404 24724 5460 25116
rect 5852 25060 5908 25340
rect 6076 25284 6132 25294
rect 5516 25004 5908 25060
rect 5964 25282 6132 25284
rect 5964 25230 6078 25282
rect 6130 25230 6132 25282
rect 5964 25228 6132 25230
rect 5516 24834 5572 25004
rect 5516 24782 5518 24834
rect 5570 24782 5572 24834
rect 5516 24770 5572 24782
rect 5404 22372 5460 24668
rect 5628 24498 5684 24510
rect 5628 24446 5630 24498
rect 5682 24446 5684 24498
rect 5628 23156 5684 24446
rect 5964 23380 6020 25228
rect 6076 25218 6132 25228
rect 6076 24724 6132 24734
rect 6076 24630 6132 24668
rect 6188 24722 6244 29260
rect 6412 29222 6468 29260
rect 6636 28754 6692 29372
rect 6748 28868 6804 28878
rect 6748 28774 6804 28812
rect 6636 28702 6638 28754
rect 6690 28702 6692 28754
rect 6636 28690 6692 28702
rect 6860 26908 6916 30604
rect 6972 30210 7028 31164
rect 7196 30436 7252 31892
rect 7420 30660 7476 33182
rect 7532 33122 7588 33134
rect 7532 33070 7534 33122
rect 7586 33070 7588 33122
rect 7532 32900 7588 33070
rect 7644 33124 7700 34300
rect 8204 33348 8260 33358
rect 8204 33254 8260 33292
rect 7756 33124 7812 33134
rect 7644 33068 7756 33124
rect 7756 33030 7812 33068
rect 7532 32844 7924 32900
rect 7868 32788 7924 32844
rect 7868 32786 8148 32788
rect 7868 32734 7870 32786
rect 7922 32734 8148 32786
rect 7868 32732 8148 32734
rect 7868 32722 7924 32732
rect 7756 32676 7812 32686
rect 7756 32582 7812 32620
rect 8092 31780 8148 32732
rect 8092 31714 8148 31724
rect 7420 30594 7476 30604
rect 7196 30380 7588 30436
rect 6972 30158 6974 30210
rect 7026 30158 7028 30210
rect 6972 30146 7028 30158
rect 7420 30210 7476 30222
rect 7420 30158 7422 30210
rect 7474 30158 7476 30210
rect 7084 30100 7140 30110
rect 7084 30006 7140 30044
rect 7420 29316 7476 30158
rect 7420 29250 7476 29260
rect 7532 26908 7588 30380
rect 6860 26852 7140 26908
rect 7308 26852 7364 26862
rect 7084 26514 7140 26852
rect 7084 26462 7086 26514
rect 7138 26462 7140 26514
rect 7084 26450 7140 26462
rect 7196 26850 7364 26852
rect 7196 26798 7310 26850
rect 7362 26798 7364 26850
rect 7196 26796 7364 26798
rect 6972 26402 7028 26414
rect 6972 26350 6974 26402
rect 7026 26350 7028 26402
rect 6524 26292 6580 26302
rect 6748 26292 6804 26302
rect 6524 26290 6692 26292
rect 6524 26238 6526 26290
rect 6578 26238 6692 26290
rect 6524 26236 6692 26238
rect 6524 26226 6580 26236
rect 6636 26180 6692 26236
rect 6748 26198 6804 26236
rect 6300 25396 6356 25406
rect 6524 25396 6580 25406
rect 6300 25394 6524 25396
rect 6300 25342 6302 25394
rect 6354 25342 6524 25394
rect 6300 25340 6524 25342
rect 6300 25330 6356 25340
rect 6188 24670 6190 24722
rect 6242 24670 6244 24722
rect 6188 23716 6244 24670
rect 6412 24722 6468 24734
rect 6412 24670 6414 24722
rect 6466 24670 6468 24722
rect 6300 24612 6356 24622
rect 6300 24518 6356 24556
rect 6188 23650 6244 23660
rect 6412 23492 6468 24670
rect 6188 23436 6468 23492
rect 6076 23380 6132 23390
rect 6188 23380 6244 23436
rect 5964 23324 6076 23380
rect 6132 23324 6244 23380
rect 5852 23156 5908 23166
rect 5628 23154 6020 23156
rect 5628 23102 5854 23154
rect 5906 23102 6020 23154
rect 5628 23100 6020 23102
rect 5852 23090 5908 23100
rect 5740 22484 5796 22494
rect 5740 22390 5796 22428
rect 5628 22372 5684 22382
rect 5404 22370 5684 22372
rect 5404 22318 5630 22370
rect 5682 22318 5684 22370
rect 5404 22316 5684 22318
rect 4844 21532 5012 21588
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 3836 20514 3892 20524
rect 1932 17666 1988 19964
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 2604 18228 2660 18238
rect 2604 17778 2660 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 2604 17726 2606 17778
rect 2658 17726 2660 17778
rect 2604 17714 2660 17726
rect 4732 17778 4788 17790
rect 4732 17726 4734 17778
rect 4786 17726 4788 17778
rect 1932 17614 1934 17666
rect 1986 17614 1988 17666
rect 1932 15314 1988 17614
rect 4732 17668 4788 17726
rect 4732 17602 4788 17612
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 2716 15876 2772 15886
rect 2716 15426 2772 15820
rect 4844 15764 4900 21532
rect 5516 21474 5572 21486
rect 5516 21422 5518 21474
rect 5570 21422 5572 21474
rect 5292 19908 5348 19918
rect 5516 19908 5572 21422
rect 5180 19852 5292 19908
rect 5348 19852 5572 19908
rect 4956 18452 5012 18490
rect 4956 18386 5012 18396
rect 4956 18228 5012 18238
rect 5180 18228 5236 19852
rect 5292 19842 5348 19852
rect 5628 19796 5684 22316
rect 5852 22148 5908 22158
rect 5852 22054 5908 22092
rect 5964 21140 6020 23100
rect 6076 22370 6132 23324
rect 6300 23268 6356 23278
rect 6524 23268 6580 25340
rect 6636 24834 6692 26124
rect 6748 25506 6804 25518
rect 6748 25454 6750 25506
rect 6802 25454 6804 25506
rect 6748 25396 6804 25454
rect 6748 25330 6804 25340
rect 6972 25284 7028 26350
rect 7084 26292 7140 26302
rect 7084 25506 7140 26236
rect 7084 25454 7086 25506
rect 7138 25454 7140 25506
rect 7084 25442 7140 25454
rect 7196 25284 7252 26796
rect 7308 26786 7364 26796
rect 7420 26852 7588 26908
rect 7756 28868 7812 28878
rect 7308 26180 7364 26190
rect 7308 26086 7364 26124
rect 7420 25730 7476 26852
rect 7756 26290 7812 28812
rect 7756 26238 7758 26290
rect 7810 26238 7812 26290
rect 7756 26226 7812 26238
rect 8204 26180 8260 26190
rect 8204 26178 8372 26180
rect 8204 26126 8206 26178
rect 8258 26126 8372 26178
rect 8204 26124 8372 26126
rect 8204 26114 8260 26124
rect 7420 25678 7422 25730
rect 7474 25678 7476 25730
rect 7420 25666 7476 25678
rect 7308 25284 7364 25294
rect 6972 25228 7308 25284
rect 7308 25190 7364 25228
rect 7756 25284 7812 25294
rect 7756 25190 7812 25228
rect 8316 24948 8372 26124
rect 8428 25844 8484 34862
rect 8652 34580 8708 36316
rect 8876 35140 8932 39342
rect 9884 37938 9940 37950
rect 9884 37886 9886 37938
rect 9938 37886 9940 37938
rect 9548 36708 9604 36718
rect 9548 35140 9604 36652
rect 9884 35924 9940 37886
rect 9884 35858 9940 35868
rect 9660 35588 9716 35598
rect 9884 35588 9940 35598
rect 9716 35586 9940 35588
rect 9716 35534 9886 35586
rect 9938 35534 9940 35586
rect 9716 35532 9940 35534
rect 9660 35522 9716 35532
rect 9884 35522 9940 35532
rect 9548 35084 9716 35140
rect 8876 35074 8932 35084
rect 9324 35028 9380 35038
rect 9324 34914 9380 34972
rect 9324 34862 9326 34914
rect 9378 34862 9380 34914
rect 9324 34850 9380 34862
rect 9548 34914 9604 34926
rect 9548 34862 9550 34914
rect 9602 34862 9604 34914
rect 8764 34580 8820 34590
rect 8652 34524 8764 34580
rect 8540 34356 8596 34366
rect 8540 34262 8596 34300
rect 8764 34354 8820 34524
rect 9548 34580 9604 34862
rect 9548 34514 9604 34524
rect 8764 34302 8766 34354
rect 8818 34302 8820 34354
rect 8764 34290 8820 34302
rect 9660 34244 9716 35084
rect 9772 34916 9828 34926
rect 9772 34822 9828 34860
rect 10108 34804 10164 34814
rect 9996 34692 10052 34730
rect 10108 34710 10164 34748
rect 9996 34626 10052 34636
rect 10220 34356 10276 40348
rect 10444 38052 10500 40348
rect 10556 40292 10612 40302
rect 10556 40198 10612 40236
rect 12684 40290 12740 41916
rect 13244 41860 13300 45200
rect 17052 45108 17108 45200
rect 17388 45108 17444 45276
rect 17052 45052 17444 45108
rect 17836 43708 17892 45276
rect 20832 45200 20944 46000
rect 21196 45276 21700 45332
rect 20860 45108 20916 45200
rect 21196 45108 21252 45276
rect 20860 45052 21252 45108
rect 17836 43652 18340 43708
rect 18284 42194 18340 43652
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 18284 42142 18286 42194
rect 18338 42142 18340 42194
rect 18284 42130 18340 42142
rect 13468 41972 13524 41982
rect 13468 41878 13524 41916
rect 16156 41972 16212 41982
rect 13244 41794 13300 41804
rect 14476 41860 14532 41870
rect 14476 41766 14532 41804
rect 13356 40404 13412 40414
rect 13356 40310 13412 40348
rect 12684 40238 12686 40290
rect 12738 40238 12740 40290
rect 12684 40226 12740 40238
rect 14028 40292 14084 40302
rect 14028 40290 14644 40292
rect 14028 40238 14030 40290
rect 14082 40238 14644 40290
rect 14028 40236 14644 40238
rect 14028 40226 14084 40236
rect 14588 39506 14644 40236
rect 16156 40290 16212 41916
rect 17276 41972 17332 41982
rect 21084 41972 21140 41982
rect 17276 41878 17332 41916
rect 20524 41970 21140 41972
rect 20524 41918 21086 41970
rect 21138 41918 21140 41970
rect 20524 41916 21140 41918
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 16940 40404 16996 40414
rect 16156 40238 16158 40290
rect 16210 40238 16212 40290
rect 16156 40226 16212 40238
rect 16716 40348 16940 40404
rect 14588 39454 14590 39506
rect 14642 39454 14644 39506
rect 14588 39442 14644 39454
rect 14924 39506 14980 39518
rect 14924 39454 14926 39506
rect 14978 39454 14980 39506
rect 12908 39394 12964 39406
rect 12908 39342 12910 39394
rect 12962 39342 12964 39394
rect 10556 38052 10612 38062
rect 11116 38052 11172 38062
rect 10444 38050 11116 38052
rect 10444 37998 10558 38050
rect 10610 37998 11116 38050
rect 10444 37996 11116 37998
rect 10556 37986 10612 37996
rect 11004 37266 11060 37996
rect 11116 37958 11172 37996
rect 12908 38052 12964 39342
rect 14924 38612 14980 39454
rect 14924 38546 14980 38556
rect 16380 39396 16436 39406
rect 16716 39396 16772 40348
rect 16940 40310 16996 40348
rect 17612 40404 17668 40414
rect 17612 40310 17668 40348
rect 20076 40404 20132 40414
rect 18396 40290 18452 40302
rect 18396 40238 18398 40290
rect 18450 40238 18452 40290
rect 18396 39730 18452 40238
rect 18396 39678 18398 39730
rect 18450 39678 18452 39730
rect 18396 39666 18452 39678
rect 18956 40292 19012 40302
rect 18956 39730 19012 40236
rect 20076 39732 20132 40348
rect 20524 40290 20580 41916
rect 21084 41906 21140 41916
rect 21644 41860 21700 45276
rect 24640 45200 24752 46000
rect 28448 45200 28560 46000
rect 32256 45200 32368 46000
rect 32620 45276 33124 45332
rect 22092 41860 22148 41870
rect 21644 41858 22148 41860
rect 21644 41806 22094 41858
rect 22146 41806 22148 41858
rect 21644 41804 22148 41806
rect 22092 41794 22148 41804
rect 24668 41860 24724 45200
rect 24892 41972 24948 41982
rect 24668 41794 24724 41804
rect 24780 41970 24948 41972
rect 24780 41918 24894 41970
rect 24946 41918 24948 41970
rect 24780 41916 24948 41918
rect 24780 40852 24836 41916
rect 24892 41906 24948 41916
rect 25900 41860 25956 41870
rect 28476 41860 28532 45200
rect 32284 45108 32340 45200
rect 32620 45108 32676 45276
rect 32284 45052 32676 45108
rect 33068 43708 33124 45276
rect 36064 45200 36176 46000
rect 36428 45276 36932 45332
rect 36092 45108 36148 45200
rect 36428 45108 36484 45276
rect 36092 45052 36484 45108
rect 33068 43652 33572 43708
rect 33516 42194 33572 43652
rect 33516 42142 33518 42194
rect 33570 42142 33572 42194
rect 33516 42130 33572 42142
rect 30828 41972 30884 41982
rect 30604 41970 30884 41972
rect 30604 41918 30830 41970
rect 30882 41918 30884 41970
rect 30604 41916 30884 41918
rect 28924 41860 28980 41870
rect 28476 41858 28980 41860
rect 28476 41806 28926 41858
rect 28978 41806 28980 41858
rect 28476 41804 28980 41806
rect 25900 41766 25956 41804
rect 28924 41794 28980 41804
rect 23548 40796 24836 40852
rect 20524 40238 20526 40290
rect 20578 40238 20580 40290
rect 20524 40226 20580 40238
rect 20636 40516 20692 40526
rect 20188 39732 20244 39742
rect 18956 39678 18958 39730
rect 19010 39678 19012 39730
rect 18956 39666 19012 39678
rect 19516 39730 20244 39732
rect 19516 39678 20190 39730
rect 20242 39678 20244 39730
rect 19516 39676 20244 39678
rect 16380 39394 16772 39396
rect 16380 39342 16382 39394
rect 16434 39342 16772 39394
rect 16380 39340 16772 39342
rect 17948 39618 18004 39630
rect 17948 39566 17950 39618
rect 18002 39566 18004 39618
rect 12908 37986 12964 37996
rect 14252 38052 14308 38062
rect 14252 37490 14308 37996
rect 14252 37438 14254 37490
rect 14306 37438 14308 37490
rect 14252 37426 14308 37438
rect 15820 38050 15876 38062
rect 15820 37998 15822 38050
rect 15874 37998 15876 38050
rect 15820 37828 15876 37998
rect 11004 37214 11006 37266
rect 11058 37214 11060 37266
rect 11004 37202 11060 37214
rect 11676 37154 11732 37166
rect 11676 37102 11678 37154
rect 11730 37102 11732 37154
rect 10892 35924 10948 35934
rect 10108 34300 10276 34356
rect 10332 34692 10388 34702
rect 10668 34692 10724 34702
rect 10388 34690 10724 34692
rect 10388 34638 10670 34690
rect 10722 34638 10724 34690
rect 10388 34636 10724 34638
rect 9996 34244 10052 34254
rect 9100 34242 10052 34244
rect 9100 34190 9998 34242
rect 10050 34190 10052 34242
rect 9100 34188 10052 34190
rect 8876 34130 8932 34142
rect 8876 34078 8878 34130
rect 8930 34078 8932 34130
rect 8876 34020 8932 34078
rect 8876 33954 8932 33964
rect 8540 33460 8596 33470
rect 8540 32786 8596 33404
rect 8540 32734 8542 32786
rect 8594 32734 8596 32786
rect 8540 32722 8596 32734
rect 9100 31948 9156 34188
rect 9996 34178 10052 34188
rect 9660 34020 9716 34030
rect 9660 33926 9716 33964
rect 8540 31892 8596 31902
rect 8540 31798 8596 31836
rect 8764 31892 9156 31948
rect 9772 32676 9828 32686
rect 8764 31778 8820 31892
rect 8988 31780 9044 31790
rect 8764 31726 8766 31778
rect 8818 31726 8820 31778
rect 8764 28644 8820 31726
rect 8876 31724 8988 31780
rect 8876 30210 8932 31724
rect 8988 31686 9044 31724
rect 9436 31556 9492 31566
rect 9436 31462 9492 31500
rect 8876 30158 8878 30210
rect 8930 30158 8932 30210
rect 8876 30146 8932 30158
rect 9212 30212 9268 30222
rect 9212 30118 9268 30156
rect 9772 29652 9828 32620
rect 10108 31948 10164 34300
rect 10220 34132 10276 34142
rect 10332 34132 10388 34636
rect 10668 34626 10724 34636
rect 10892 34354 10948 35868
rect 11676 35364 11732 37102
rect 13804 37156 13860 37166
rect 13804 37154 13972 37156
rect 13804 37102 13806 37154
rect 13858 37102 13972 37154
rect 13804 37100 13972 37102
rect 13804 37090 13860 37100
rect 11676 35308 11956 35364
rect 11004 35028 11060 35038
rect 11060 34972 11284 35028
rect 11004 34934 11060 34972
rect 10892 34302 10894 34354
rect 10946 34302 10948 34354
rect 10892 34290 10948 34302
rect 11116 34804 11172 34814
rect 10220 34130 10388 34132
rect 10220 34078 10222 34130
rect 10274 34078 10388 34130
rect 10220 34076 10388 34078
rect 10556 34244 10612 34254
rect 10556 34130 10612 34188
rect 10556 34078 10558 34130
rect 10610 34078 10612 34130
rect 10220 34020 10276 34076
rect 10556 34066 10612 34078
rect 10668 34130 10724 34142
rect 10668 34078 10670 34130
rect 10722 34078 10724 34130
rect 10220 33124 10276 33964
rect 10332 33908 10388 33918
rect 10668 33908 10724 34078
rect 10332 33906 10724 33908
rect 10332 33854 10334 33906
rect 10386 33854 10724 33906
rect 10332 33852 10724 33854
rect 11004 34130 11060 34142
rect 11004 34078 11006 34130
rect 11058 34078 11060 34130
rect 10332 33842 10388 33852
rect 10668 33124 10724 33134
rect 10220 33122 10724 33124
rect 10220 33070 10670 33122
rect 10722 33070 10724 33122
rect 10220 33068 10724 33070
rect 10444 32228 10500 32238
rect 10108 31892 10276 31948
rect 10220 31218 10276 31892
rect 10220 31166 10222 31218
rect 10274 31166 10276 31218
rect 10220 31154 10276 31166
rect 10108 30994 10164 31006
rect 10108 30942 10110 30994
rect 10162 30942 10164 30994
rect 9884 30884 9940 30894
rect 10108 30884 10164 30942
rect 9884 30882 10164 30884
rect 9884 30830 9886 30882
rect 9938 30830 10164 30882
rect 9884 30828 10164 30830
rect 9884 30818 9940 30828
rect 9996 29652 10052 29662
rect 9772 29650 10052 29652
rect 9772 29598 9998 29650
rect 10050 29598 10052 29650
rect 9772 29596 10052 29598
rect 9996 29586 10052 29596
rect 10108 29540 10164 30828
rect 10220 30772 10276 30782
rect 10220 30678 10276 30716
rect 10108 29474 10164 29484
rect 10444 29538 10500 32172
rect 10668 31668 10724 33068
rect 11004 33012 11060 34078
rect 10892 32956 11060 33012
rect 10668 31602 10724 31612
rect 10780 31780 10836 31790
rect 10444 29486 10446 29538
rect 10498 29486 10500 29538
rect 10444 29474 10500 29486
rect 9436 29428 9492 29438
rect 9436 28866 9492 29372
rect 9436 28814 9438 28866
rect 9490 28814 9492 28866
rect 9436 28802 9492 28814
rect 9772 29426 9828 29438
rect 9772 29374 9774 29426
rect 9826 29374 9828 29426
rect 9772 28868 9828 29374
rect 10220 29428 10276 29438
rect 10220 29334 10276 29372
rect 9772 28802 9828 28812
rect 9996 29314 10052 29326
rect 9996 29262 9998 29314
rect 10050 29262 10052 29314
rect 9324 28756 9380 28766
rect 9324 28662 9380 28700
rect 8764 28578 8820 28588
rect 9996 27972 10052 29262
rect 10780 28868 10836 31724
rect 10668 28812 10836 28868
rect 10332 28754 10388 28766
rect 10332 28702 10334 28754
rect 10386 28702 10388 28754
rect 10108 28644 10164 28654
rect 10108 28550 10164 28588
rect 9996 27906 10052 27916
rect 8428 25778 8484 25788
rect 8764 25284 8820 25294
rect 8652 24948 8708 24958
rect 8316 24946 8708 24948
rect 8316 24894 8654 24946
rect 8706 24894 8708 24946
rect 8316 24892 8708 24894
rect 8652 24882 8708 24892
rect 6636 24782 6638 24834
rect 6690 24782 6692 24834
rect 6636 24770 6692 24782
rect 8204 23380 8260 23390
rect 8204 23286 8260 23324
rect 6300 23266 6580 23268
rect 6300 23214 6302 23266
rect 6354 23214 6580 23266
rect 6300 23212 6580 23214
rect 6300 23202 6356 23212
rect 6076 22318 6078 22370
rect 6130 22318 6132 22370
rect 6076 22306 6132 22318
rect 6188 23154 6244 23166
rect 6188 23102 6190 23154
rect 6242 23102 6244 23154
rect 6188 22484 6244 23102
rect 7980 23154 8036 23166
rect 7980 23102 7982 23154
rect 8034 23102 8036 23154
rect 6188 21252 6244 22428
rect 6972 23044 7028 23054
rect 6300 22260 6356 22270
rect 6300 22166 6356 22204
rect 6188 21196 6356 21252
rect 5964 21084 6244 21140
rect 5516 19740 5684 19796
rect 5516 18564 5572 19740
rect 6076 19346 6132 19358
rect 6076 19294 6078 19346
rect 6130 19294 6132 19346
rect 6076 18788 6132 19294
rect 6188 19124 6244 21084
rect 6300 19348 6356 21196
rect 6412 19348 6468 19358
rect 6300 19346 6692 19348
rect 6300 19294 6414 19346
rect 6466 19294 6692 19346
rect 6300 19292 6692 19294
rect 6412 19282 6468 19292
rect 6188 19122 6580 19124
rect 6188 19070 6190 19122
rect 6242 19070 6580 19122
rect 6188 19068 6580 19070
rect 6188 19058 6244 19068
rect 6524 18900 6580 19068
rect 6412 18844 6580 18900
rect 5628 18732 6356 18788
rect 5628 18674 5684 18732
rect 5628 18622 5630 18674
rect 5682 18622 5684 18674
rect 5628 18610 5684 18622
rect 5516 18498 5572 18508
rect 5852 18450 5908 18462
rect 6188 18452 6244 18462
rect 5852 18398 5854 18450
rect 5906 18398 5908 18450
rect 5740 18338 5796 18350
rect 5740 18286 5742 18338
rect 5794 18286 5796 18338
rect 4956 18134 5012 18172
rect 5068 18172 5236 18228
rect 5292 18228 5348 18238
rect 5740 18228 5796 18286
rect 5292 18226 5796 18228
rect 5292 18174 5294 18226
rect 5346 18174 5796 18226
rect 5292 18172 5796 18174
rect 5852 18340 5908 18398
rect 4956 17108 5012 17118
rect 5068 17108 5124 18172
rect 5292 18162 5348 18172
rect 4956 17106 5124 17108
rect 4956 17054 4958 17106
rect 5010 17054 5124 17106
rect 4956 17052 5124 17054
rect 4956 17042 5012 17052
rect 4844 15698 4900 15708
rect 2716 15374 2718 15426
rect 2770 15374 2772 15426
rect 2716 15362 2772 15374
rect 4844 15428 4900 15438
rect 1932 15262 1934 15314
rect 1986 15262 1988 15314
rect 1932 12178 1988 15262
rect 4844 15202 4900 15372
rect 4844 15150 4846 15202
rect 4898 15150 4900 15202
rect 4844 15138 4900 15150
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 5068 14308 5124 17052
rect 5740 17668 5796 17678
rect 5740 15426 5796 17612
rect 5852 17556 5908 18284
rect 5964 18450 6244 18452
rect 5964 18398 6190 18450
rect 6242 18398 6244 18450
rect 5964 18396 6244 18398
rect 5964 17780 6020 18396
rect 6188 18386 6244 18396
rect 5964 17714 6020 17724
rect 6300 17668 6356 18732
rect 6412 18228 6468 18844
rect 6524 18564 6580 18574
rect 6524 18450 6580 18508
rect 6524 18398 6526 18450
rect 6578 18398 6580 18450
rect 6524 18386 6580 18398
rect 6412 18162 6468 18172
rect 6636 18116 6692 19292
rect 6860 19012 6916 19022
rect 6860 18918 6916 18956
rect 6972 18674 7028 22988
rect 7980 23044 8036 23102
rect 7980 22978 8036 22988
rect 8428 22484 8484 22494
rect 8428 22390 8484 22428
rect 6972 18622 6974 18674
rect 7026 18622 7028 18674
rect 6972 18610 7028 18622
rect 7084 18900 7140 18910
rect 6636 18050 6692 18060
rect 6748 18450 6804 18462
rect 6748 18398 6750 18450
rect 6802 18398 6804 18450
rect 6748 18340 6804 18398
rect 6860 18452 6916 18462
rect 6860 18358 6916 18396
rect 6748 17892 6804 18284
rect 6524 17836 7028 17892
rect 6412 17668 6468 17678
rect 6300 17666 6468 17668
rect 6300 17614 6414 17666
rect 6466 17614 6468 17666
rect 6300 17612 6468 17614
rect 6412 17602 6468 17612
rect 5964 17556 6020 17566
rect 5852 17554 6020 17556
rect 5852 17502 5966 17554
rect 6018 17502 6020 17554
rect 5852 17500 6020 17502
rect 5964 17490 6020 17500
rect 6524 17554 6580 17836
rect 6972 17666 7028 17836
rect 7084 17780 7140 18844
rect 7084 17714 7140 17724
rect 7196 18450 7252 18462
rect 7532 18452 7588 18462
rect 7196 18398 7198 18450
rect 7250 18398 7252 18450
rect 6972 17614 6974 17666
rect 7026 17614 7028 17666
rect 6972 17602 7028 17614
rect 6524 17502 6526 17554
rect 6578 17502 6580 17554
rect 6524 17490 6580 17502
rect 6748 17444 6804 17454
rect 6748 17350 6804 17388
rect 7084 17442 7140 17454
rect 7084 17390 7086 17442
rect 7138 17390 7140 17442
rect 5740 15374 5742 15426
rect 5794 15374 5796 15426
rect 5740 15362 5796 15374
rect 6860 15428 6916 15438
rect 7084 15428 7140 17390
rect 7196 17444 7252 18398
rect 7308 18450 7588 18452
rect 7308 18398 7534 18450
rect 7586 18398 7588 18450
rect 7308 18396 7588 18398
rect 7308 17666 7364 18396
rect 7532 18386 7588 18396
rect 7756 18226 7812 18238
rect 7756 18174 7758 18226
rect 7810 18174 7812 18226
rect 7756 18116 7812 18174
rect 7980 18228 8036 18238
rect 7980 18134 8036 18172
rect 8092 18226 8148 18238
rect 8092 18174 8094 18226
rect 8146 18174 8148 18226
rect 7756 18050 7812 18060
rect 7308 17614 7310 17666
rect 7362 17614 7364 17666
rect 7308 17602 7364 17614
rect 7980 17780 8036 17790
rect 7420 17444 7476 17454
rect 7196 17388 7420 17444
rect 7420 16098 7476 17388
rect 7420 16046 7422 16098
rect 7474 16046 7476 16098
rect 7420 16034 7476 16046
rect 7756 16098 7812 16110
rect 7756 16046 7758 16098
rect 7810 16046 7812 16098
rect 7756 15988 7812 16046
rect 7868 16100 7924 16110
rect 7868 16006 7924 16044
rect 7756 15922 7812 15932
rect 7532 15876 7588 15886
rect 7532 15782 7588 15820
rect 7980 15540 8036 17724
rect 7868 15484 8036 15540
rect 6916 15372 7140 15428
rect 7756 15426 7812 15438
rect 7756 15374 7758 15426
rect 7810 15374 7812 15426
rect 6860 15314 6916 15372
rect 6860 15262 6862 15314
rect 6914 15262 6916 15314
rect 6860 15250 6916 15262
rect 7308 15316 7364 15326
rect 7308 15222 7364 15260
rect 7756 15148 7812 15374
rect 7644 15092 7812 15148
rect 6860 14420 6916 14430
rect 6748 14364 6860 14420
rect 5068 14306 5236 14308
rect 5068 14254 5070 14306
rect 5122 14254 5236 14306
rect 5068 14252 5236 14254
rect 5068 14242 5124 14252
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2604 12292 2660 12302
rect 2604 12198 2660 12236
rect 1932 12126 1934 12178
rect 1986 12126 1988 12178
rect 1932 12114 1988 12126
rect 4732 12180 4788 12190
rect 4732 12066 4788 12124
rect 4732 12014 4734 12066
rect 4786 12014 4788 12066
rect 4732 12002 4788 12014
rect 5180 12066 5236 14252
rect 6076 13076 6132 13086
rect 6076 12180 6132 13020
rect 6300 12852 6356 12862
rect 6300 12402 6356 12796
rect 6300 12350 6302 12402
rect 6354 12350 6356 12402
rect 6300 12338 6356 12350
rect 6076 12086 6132 12124
rect 5180 12014 5182 12066
rect 5234 12014 5236 12066
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4508 9604 4564 9614
rect 4508 9154 4564 9548
rect 4508 9102 4510 9154
rect 4562 9102 4564 9154
rect 4508 9090 4564 9102
rect 3836 9044 3892 9054
rect 3836 8950 3892 8988
rect 5180 9044 5236 12014
rect 6636 11396 6692 11406
rect 6748 11396 6804 14364
rect 6860 14354 6916 14364
rect 7644 13076 7700 15092
rect 7756 14420 7812 14430
rect 7756 13970 7812 14364
rect 7756 13918 7758 13970
rect 7810 13918 7812 13970
rect 7756 13906 7812 13918
rect 7644 13010 7700 13020
rect 7756 12962 7812 12974
rect 7756 12910 7758 12962
rect 7810 12910 7812 12962
rect 7756 12852 7812 12910
rect 7756 12786 7812 12796
rect 7868 12404 7924 15484
rect 7756 12348 7924 12404
rect 7980 15316 8036 15326
rect 7980 12962 8036 15260
rect 7980 12910 7982 12962
rect 8034 12910 8036 12962
rect 7644 12292 7700 12302
rect 7644 12198 7700 12236
rect 7532 12178 7588 12190
rect 7532 12126 7534 12178
rect 7586 12126 7588 12178
rect 6636 11394 6804 11396
rect 6636 11342 6638 11394
rect 6690 11342 6804 11394
rect 6636 11340 6804 11342
rect 6972 11452 7364 11508
rect 6972 11394 7028 11452
rect 6972 11342 6974 11394
rect 7026 11342 7028 11394
rect 6524 11172 6580 11182
rect 6524 9714 6580 11116
rect 6636 10724 6692 11340
rect 6972 11330 7028 11342
rect 7308 11396 7364 11452
rect 7420 11396 7476 11406
rect 7532 11396 7588 12126
rect 7308 11394 7588 11396
rect 7308 11342 7422 11394
rect 7474 11342 7588 11394
rect 7308 11340 7588 11342
rect 7420 11330 7476 11340
rect 7196 11284 7252 11294
rect 7196 11190 7252 11228
rect 6748 11170 6804 11182
rect 6748 11118 6750 11170
rect 6802 11118 6804 11170
rect 6748 10948 6804 11118
rect 7532 11172 7588 11182
rect 7532 11078 7588 11116
rect 7644 11170 7700 11182
rect 7644 11118 7646 11170
rect 7698 11118 7700 11170
rect 7644 10948 7700 11118
rect 6748 10892 7644 10948
rect 6636 10668 7252 10724
rect 7196 10612 7252 10668
rect 7196 10518 7252 10556
rect 7420 10610 7476 10892
rect 7644 10882 7700 10892
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 7308 10498 7364 10510
rect 7308 10446 7310 10498
rect 7362 10446 7364 10498
rect 7308 10164 7364 10446
rect 6748 10108 7364 10164
rect 6748 10050 6804 10108
rect 7420 10052 7476 10558
rect 7756 10612 7812 12348
rect 7868 12180 7924 12190
rect 7868 12086 7924 12124
rect 7868 11394 7924 11406
rect 7868 11342 7870 11394
rect 7922 11342 7924 11394
rect 7868 11172 7924 11342
rect 7868 11106 7924 11116
rect 7868 10612 7924 10622
rect 7756 10610 7924 10612
rect 7756 10558 7870 10610
rect 7922 10558 7924 10610
rect 7756 10556 7924 10558
rect 6748 9998 6750 10050
rect 6802 9998 6804 10050
rect 6748 9986 6804 9998
rect 7084 9996 7476 10052
rect 6524 9662 6526 9714
rect 6578 9662 6580 9714
rect 6524 9650 6580 9662
rect 6748 9828 6804 9838
rect 6636 9604 6692 9614
rect 6636 9510 6692 9548
rect 5180 8978 5236 8988
rect 6636 8932 6692 8942
rect 6748 8932 6804 9772
rect 7084 9714 7140 9996
rect 7308 9828 7364 9838
rect 7308 9734 7364 9772
rect 7084 9662 7086 9714
rect 7138 9662 7140 9714
rect 7084 9650 7140 9662
rect 7868 9604 7924 10556
rect 7980 9828 8036 12910
rect 8092 13970 8148 18174
rect 8204 16212 8260 16222
rect 8204 16100 8260 16156
rect 8204 16098 8484 16100
rect 8204 16046 8206 16098
rect 8258 16046 8484 16098
rect 8204 16044 8484 16046
rect 8204 16034 8260 16044
rect 8092 13918 8094 13970
rect 8146 13918 8148 13970
rect 8092 12962 8148 13918
rect 8092 12910 8094 12962
rect 8146 12910 8148 12962
rect 8092 12898 8148 12910
rect 8428 12404 8484 16044
rect 8540 15988 8596 15998
rect 8540 15894 8596 15932
rect 8652 15986 8708 15998
rect 8652 15934 8654 15986
rect 8706 15934 8708 15986
rect 8652 15428 8708 15934
rect 8652 15362 8708 15372
rect 8764 15204 8820 25228
rect 8876 24834 8932 24846
rect 8876 24782 8878 24834
rect 8930 24782 8932 24834
rect 8876 23940 8932 24782
rect 8988 24722 9044 24734
rect 8988 24670 8990 24722
rect 9042 24670 9044 24722
rect 8988 24276 9044 24670
rect 8988 24220 9380 24276
rect 9212 24050 9268 24062
rect 9212 23998 9214 24050
rect 9266 23998 9268 24050
rect 9100 23940 9156 23950
rect 8876 23884 9100 23940
rect 9100 23846 9156 23884
rect 8876 23716 8932 23726
rect 8876 23622 8932 23660
rect 9212 23156 9268 23998
rect 9324 24052 9380 24220
rect 9436 24052 9492 24062
rect 9324 23996 9436 24052
rect 9436 23938 9492 23996
rect 9436 23886 9438 23938
rect 9490 23886 9492 23938
rect 9436 23874 9492 23886
rect 9212 23090 9268 23100
rect 9660 23716 9716 23726
rect 9660 22932 9716 23660
rect 9884 23156 9940 23166
rect 10220 23156 10276 23166
rect 10332 23156 10388 28702
rect 10668 26908 10724 28812
rect 10780 28644 10836 28654
rect 10780 28550 10836 28588
rect 10668 26852 10836 26908
rect 9884 23042 9940 23100
rect 9884 22990 9886 23042
rect 9938 22990 9940 23042
rect 9884 22978 9940 22990
rect 9996 23154 10388 23156
rect 9996 23102 10222 23154
rect 10274 23102 10388 23154
rect 9996 23100 10388 23102
rect 10668 26290 10724 26302
rect 10668 26238 10670 26290
rect 10722 26238 10724 26290
rect 9660 22876 9828 22932
rect 9772 22370 9828 22876
rect 9772 22318 9774 22370
rect 9826 22318 9828 22370
rect 9772 22306 9828 22318
rect 9884 22260 9940 22270
rect 9996 22260 10052 23100
rect 10220 23090 10276 23100
rect 9884 22258 10052 22260
rect 9884 22206 9886 22258
rect 9938 22206 10052 22258
rect 9884 22204 10052 22206
rect 10220 22932 10276 22942
rect 10668 22932 10724 26238
rect 10780 25956 10836 26852
rect 10892 26178 10948 32956
rect 11116 32900 11172 34748
rect 11004 32844 11172 32900
rect 11004 29204 11060 32844
rect 11228 31948 11284 34972
rect 11676 34804 11732 34814
rect 11676 34354 11732 34748
rect 11676 34302 11678 34354
rect 11730 34302 11732 34354
rect 11676 34290 11732 34302
rect 11340 34130 11396 34142
rect 11340 34078 11342 34130
rect 11394 34078 11396 34130
rect 11340 34020 11396 34078
rect 11340 33954 11396 33964
rect 11900 33458 11956 35308
rect 13804 35026 13860 35038
rect 13804 34974 13806 35026
rect 13858 34974 13860 35026
rect 12012 34244 12068 34254
rect 12068 34188 12180 34244
rect 12012 34150 12068 34188
rect 12124 33684 12180 34188
rect 12460 34020 12516 34030
rect 12796 34020 12852 34030
rect 12460 34018 12796 34020
rect 12460 33966 12462 34018
rect 12514 33966 12796 34018
rect 12460 33964 12796 33966
rect 12460 33908 12516 33964
rect 12124 33618 12180 33628
rect 12348 33852 12516 33908
rect 11900 33406 11902 33458
rect 11954 33406 11956 33458
rect 11900 33394 11956 33406
rect 12012 33572 12068 33582
rect 11788 33234 11844 33246
rect 11788 33182 11790 33234
rect 11842 33182 11844 33234
rect 11788 32786 11844 33182
rect 11788 32734 11790 32786
rect 11842 32734 11844 32786
rect 11788 32722 11844 32734
rect 11900 32674 11956 32686
rect 11900 32622 11902 32674
rect 11954 32622 11956 32674
rect 11900 32228 11956 32622
rect 11900 32162 11956 32172
rect 11116 31892 11284 31948
rect 11116 31780 11172 31892
rect 11116 31714 11172 31724
rect 11452 31668 11508 31678
rect 11116 31554 11172 31566
rect 11116 31502 11118 31554
rect 11170 31502 11172 31554
rect 11116 31444 11172 31502
rect 11116 30772 11172 31388
rect 11116 29764 11172 30716
rect 11452 31554 11508 31612
rect 11452 31502 11454 31554
rect 11506 31502 11508 31554
rect 11452 30324 11508 31502
rect 12012 31106 12068 33516
rect 12348 33346 12404 33852
rect 12348 33294 12350 33346
rect 12402 33294 12404 33346
rect 12348 33282 12404 33294
rect 12460 33684 12516 33694
rect 12124 33236 12180 33246
rect 12460 33236 12516 33628
rect 12796 33458 12852 33964
rect 12796 33406 12798 33458
rect 12850 33406 12852 33458
rect 12796 33394 12852 33406
rect 13804 33348 13860 34974
rect 13804 33282 13860 33292
rect 12124 33234 12292 33236
rect 12124 33182 12126 33234
rect 12178 33182 12292 33234
rect 12124 33180 12292 33182
rect 12124 33170 12180 33180
rect 12124 32788 12180 32798
rect 12124 32694 12180 32732
rect 12012 31054 12014 31106
rect 12066 31054 12068 31106
rect 12012 31042 12068 31054
rect 11452 30268 11956 30324
rect 11228 30212 11284 30222
rect 11228 30118 11284 30156
rect 11564 30100 11620 30110
rect 11564 30006 11620 30044
rect 11676 29988 11732 29998
rect 11676 29894 11732 29932
rect 11116 29708 11284 29764
rect 11228 29652 11284 29708
rect 11228 29596 11508 29652
rect 11116 29538 11172 29550
rect 11116 29486 11118 29538
rect 11170 29486 11172 29538
rect 11116 29428 11172 29486
rect 11116 29362 11172 29372
rect 11228 29426 11284 29438
rect 11228 29374 11230 29426
rect 11282 29374 11284 29426
rect 11116 29204 11172 29214
rect 11004 29202 11172 29204
rect 11004 29150 11118 29202
rect 11170 29150 11172 29202
rect 11004 29148 11172 29150
rect 11116 29138 11172 29148
rect 11228 27076 11284 29374
rect 11452 28532 11508 29596
rect 11676 29428 11732 29438
rect 11676 29334 11732 29372
rect 11452 28476 11732 28532
rect 11004 27020 11284 27076
rect 11004 26516 11060 27020
rect 11676 26908 11732 28476
rect 11004 26422 11060 26460
rect 11452 26852 11732 26908
rect 10892 26126 10894 26178
rect 10946 26126 10948 26178
rect 10892 26114 10948 26126
rect 11228 26402 11284 26414
rect 11228 26350 11230 26402
rect 11282 26350 11284 26402
rect 11228 25956 11284 26350
rect 10780 25900 11060 25956
rect 10892 24052 10948 24062
rect 10780 23940 10836 23950
rect 10780 23846 10836 23884
rect 10220 22930 10724 22932
rect 10220 22878 10222 22930
rect 10274 22878 10724 22930
rect 10220 22876 10724 22878
rect 10220 22260 10276 22876
rect 9884 22148 9940 22204
rect 10220 22194 10276 22204
rect 10892 22258 10948 23996
rect 10892 22206 10894 22258
rect 10946 22206 10948 22258
rect 10892 22194 10948 22206
rect 9884 22082 9940 22092
rect 11004 22036 11060 25900
rect 11228 25284 11284 25900
rect 11228 25218 11284 25228
rect 11340 25730 11396 25742
rect 11340 25678 11342 25730
rect 11394 25678 11396 25730
rect 11228 24052 11284 24062
rect 11228 23938 11284 23996
rect 11228 23886 11230 23938
rect 11282 23886 11284 23938
rect 11228 23874 11284 23886
rect 11340 24052 11396 25678
rect 11452 25508 11508 26852
rect 11788 26516 11844 26526
rect 11788 26422 11844 26460
rect 11564 26290 11620 26302
rect 11564 26238 11566 26290
rect 11618 26238 11620 26290
rect 11564 25730 11620 26238
rect 11564 25678 11566 25730
rect 11618 25678 11620 25730
rect 11564 25666 11620 25678
rect 11452 25452 11732 25508
rect 11452 25284 11508 25294
rect 11452 25190 11508 25228
rect 11452 24052 11508 24062
rect 11340 24050 11508 24052
rect 11340 23998 11454 24050
rect 11506 23998 11508 24050
rect 11340 23996 11508 23998
rect 11340 23716 11396 23996
rect 11452 23986 11508 23996
rect 11116 23660 11396 23716
rect 11452 23828 11508 23838
rect 11116 23154 11172 23660
rect 11228 23380 11284 23390
rect 11228 23286 11284 23324
rect 11452 23380 11508 23772
rect 11452 23286 11508 23324
rect 11116 23102 11118 23154
rect 11170 23102 11172 23154
rect 11116 23090 11172 23102
rect 11228 23156 11284 23166
rect 11564 23156 11620 23166
rect 11228 22370 11284 23100
rect 11452 23154 11620 23156
rect 11452 23102 11566 23154
rect 11618 23102 11620 23154
rect 11452 23100 11620 23102
rect 11228 22318 11230 22370
rect 11282 22318 11284 22370
rect 11228 22306 11284 22318
rect 11340 23042 11396 23054
rect 11340 22990 11342 23042
rect 11394 22990 11396 23042
rect 10780 21980 11060 22036
rect 10556 20914 10612 20926
rect 10556 20862 10558 20914
rect 10610 20862 10612 20914
rect 9100 20804 9156 20814
rect 9100 16212 9156 20748
rect 10556 20130 10612 20862
rect 10668 20580 10724 20590
rect 10668 20486 10724 20524
rect 10556 20078 10558 20130
rect 10610 20078 10612 20130
rect 10556 20066 10612 20078
rect 10780 20132 10836 21980
rect 11340 21812 11396 22990
rect 10892 21756 11396 21812
rect 10892 21026 10948 21756
rect 10892 20974 10894 21026
rect 10946 20974 10948 21026
rect 10892 20962 10948 20974
rect 11452 21588 11508 23100
rect 11564 23090 11620 23100
rect 10892 20132 10948 20142
rect 10780 20076 10892 20132
rect 10892 20066 10948 20076
rect 9884 20018 9940 20030
rect 9884 19966 9886 20018
rect 9938 19966 9940 20018
rect 9884 19908 9940 19966
rect 9884 19842 9940 19852
rect 11228 19234 11284 19246
rect 11228 19182 11230 19234
rect 11282 19182 11284 19234
rect 9548 18562 9604 18574
rect 9548 18510 9550 18562
rect 9602 18510 9604 18562
rect 9548 18452 9604 18510
rect 9548 18386 9604 18396
rect 9884 18452 9940 18462
rect 9884 18358 9940 18396
rect 11228 18452 11284 19182
rect 11452 19122 11508 21532
rect 11452 19070 11454 19122
rect 11506 19070 11508 19122
rect 11452 19058 11508 19070
rect 11228 18228 11284 18396
rect 11676 18450 11732 25452
rect 11900 19572 11956 30268
rect 12124 30100 12180 30110
rect 12124 28868 12180 30044
rect 12124 28802 12180 28812
rect 12236 26908 12292 33180
rect 12460 32562 12516 33180
rect 13020 33124 13076 33134
rect 13020 32788 13076 33068
rect 12684 32564 12740 32574
rect 12460 32510 12462 32562
rect 12514 32510 12516 32562
rect 12460 32498 12516 32510
rect 12572 32562 12740 32564
rect 12572 32510 12686 32562
rect 12738 32510 12740 32562
rect 12572 32508 12740 32510
rect 12572 31444 12628 32508
rect 12684 32498 12740 32508
rect 13020 31948 13076 32732
rect 13916 32786 13972 37100
rect 15148 36372 15204 36382
rect 15036 33236 15092 33246
rect 15036 33142 15092 33180
rect 14700 33124 14756 33134
rect 14700 33030 14756 33068
rect 13916 32734 13918 32786
rect 13970 32734 13972 32786
rect 13580 32674 13636 32686
rect 13580 32622 13582 32674
rect 13634 32622 13636 32674
rect 13580 32228 13636 32622
rect 13580 32162 13636 32172
rect 13916 31948 13972 32734
rect 15148 32900 15204 36316
rect 15820 34692 15876 37772
rect 16380 37828 16436 39340
rect 16604 38724 16660 38734
rect 16604 38162 16660 38668
rect 17948 38724 18004 39566
rect 19516 39618 19572 39676
rect 20188 39666 20244 39676
rect 19516 39566 19518 39618
rect 19570 39566 19572 39618
rect 19516 39554 19572 39566
rect 18508 39508 18564 39518
rect 18508 39414 18564 39452
rect 19068 39508 19124 39518
rect 19068 39414 19124 39452
rect 19852 39508 19908 39518
rect 19852 39414 19908 39452
rect 20188 39508 20244 39518
rect 18284 39396 18340 39406
rect 18284 39302 18340 39340
rect 18844 39396 18900 39406
rect 18844 39302 18900 39340
rect 20076 39396 20132 39434
rect 20076 39330 20132 39340
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20188 39060 20244 39452
rect 20300 39396 20356 39406
rect 20300 39394 20468 39396
rect 20300 39342 20302 39394
rect 20354 39342 20468 39394
rect 20300 39340 20468 39342
rect 20300 39330 20356 39340
rect 20300 39060 20356 39070
rect 17948 38658 18004 38668
rect 19740 39058 20356 39060
rect 19740 39006 20302 39058
rect 20354 39006 20356 39058
rect 19740 39004 20356 39006
rect 16604 38110 16606 38162
rect 16658 38110 16660 38162
rect 16604 38098 16660 38110
rect 18732 38162 18788 38174
rect 18732 38110 18734 38162
rect 18786 38110 18788 38162
rect 16380 37762 16436 37772
rect 18732 36372 18788 38110
rect 19740 37938 19796 39004
rect 20300 38994 20356 39004
rect 20188 38836 20244 38846
rect 20412 38836 20468 39340
rect 20524 38948 20580 38958
rect 20524 38854 20580 38892
rect 20244 38780 20468 38836
rect 19740 37886 19742 37938
rect 19794 37886 19796 37938
rect 19740 37874 19796 37886
rect 20076 37940 20132 37950
rect 20076 37846 20132 37884
rect 19180 37828 19236 37838
rect 19180 37734 19236 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 38780
rect 20636 38724 20692 40460
rect 23548 39730 23604 40796
rect 24332 40628 24388 40638
rect 23884 40626 24388 40628
rect 23884 40574 24334 40626
rect 24386 40574 24388 40626
rect 23884 40572 24388 40574
rect 23660 40404 23716 40414
rect 23660 40310 23716 40348
rect 23548 39678 23550 39730
rect 23602 39678 23604 39730
rect 23548 39666 23604 39678
rect 23772 39508 23828 39518
rect 20412 38668 20692 38724
rect 23660 39452 23772 39508
rect 20412 38276 20468 38668
rect 23548 38612 23604 38622
rect 23548 38518 23604 38556
rect 20412 38182 20468 38220
rect 23548 38164 23604 38174
rect 23660 38164 23716 39452
rect 23772 39442 23828 39452
rect 23548 38162 23716 38164
rect 23548 38110 23550 38162
rect 23602 38110 23716 38162
rect 23548 38108 23716 38110
rect 23772 38836 23828 38846
rect 23548 38098 23604 38108
rect 20524 37940 20580 37950
rect 20524 37846 20580 37884
rect 21420 37940 21476 37950
rect 20412 37492 20468 37502
rect 20188 37490 20468 37492
rect 20188 37438 20414 37490
rect 20466 37438 20468 37490
rect 20188 37436 20468 37438
rect 20412 37426 20468 37436
rect 20748 37268 20804 37278
rect 20748 37266 21364 37268
rect 20748 37214 20750 37266
rect 20802 37214 21364 37266
rect 20748 37212 21364 37214
rect 20748 37202 20804 37212
rect 21308 36706 21364 37212
rect 21308 36654 21310 36706
rect 21362 36654 21364 36706
rect 21308 36642 21364 36654
rect 19740 36484 19796 36494
rect 19740 36390 19796 36428
rect 20188 36484 20244 36494
rect 18732 36306 18788 36316
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19852 35812 19908 35822
rect 20076 35812 20132 35822
rect 20188 35812 20244 36428
rect 20524 36372 20580 36382
rect 20412 36260 20468 36270
rect 20412 36166 20468 36204
rect 19852 35810 20244 35812
rect 19852 35758 19854 35810
rect 19906 35758 20078 35810
rect 20130 35758 20244 35810
rect 19852 35756 20244 35758
rect 19852 35746 19908 35756
rect 20076 35718 20132 35756
rect 20188 35474 20244 35486
rect 20188 35422 20190 35474
rect 20242 35422 20244 35474
rect 16604 34914 16660 34926
rect 16604 34862 16606 34914
rect 16658 34862 16660 34914
rect 15820 34626 15876 34636
rect 15932 34802 15988 34814
rect 15932 34750 15934 34802
rect 15986 34750 15988 34802
rect 15932 34468 15988 34750
rect 16604 34692 16660 34862
rect 20188 34916 20244 35422
rect 20188 34822 20244 34860
rect 20412 35140 20468 35150
rect 20412 34914 20468 35084
rect 20412 34862 20414 34914
rect 20466 34862 20468 34914
rect 20412 34850 20468 34862
rect 16604 34626 16660 34636
rect 17164 34692 17220 34702
rect 17164 34598 17220 34636
rect 18284 34692 18340 34702
rect 15596 34412 15988 34468
rect 15596 34354 15652 34412
rect 15596 34302 15598 34354
rect 15650 34302 15652 34354
rect 15596 34290 15652 34302
rect 15372 34130 15428 34142
rect 15372 34078 15374 34130
rect 15426 34078 15428 34130
rect 15372 33458 15428 34078
rect 15372 33406 15374 33458
rect 15426 33406 15428 33458
rect 15372 33394 15428 33406
rect 15708 34130 15764 34142
rect 15708 34078 15710 34130
rect 15762 34078 15764 34130
rect 15484 33348 15540 33358
rect 15484 33234 15540 33292
rect 15484 33182 15486 33234
rect 15538 33182 15540 33234
rect 15484 33170 15540 33182
rect 15260 33124 15316 33134
rect 15260 33030 15316 33068
rect 15148 32844 15540 32900
rect 15036 32450 15092 32462
rect 15036 32398 15038 32450
rect 15090 32398 15092 32450
rect 15036 32340 15092 32398
rect 12684 31892 13076 31948
rect 13804 31892 13972 31948
rect 14588 32116 14644 32126
rect 15036 32116 15092 32284
rect 14644 32060 15092 32116
rect 12684 31890 12740 31892
rect 12684 31838 12686 31890
rect 12738 31838 12740 31890
rect 12684 31826 12740 31838
rect 12572 31378 12628 31388
rect 13804 30210 13860 31892
rect 13804 30158 13806 30210
rect 13858 30158 13860 30210
rect 13804 30146 13860 30158
rect 14588 30212 14644 32060
rect 15036 31220 15092 31230
rect 14588 30118 14644 30156
rect 14924 30322 14980 30334
rect 14924 30270 14926 30322
rect 14978 30270 14980 30322
rect 14700 30100 14756 30110
rect 13916 29986 13972 29998
rect 13916 29934 13918 29986
rect 13970 29934 13972 29986
rect 13468 28756 13524 28766
rect 12124 26852 12292 26908
rect 12908 28084 12964 28094
rect 12908 27074 12964 28028
rect 12908 27022 12910 27074
rect 12962 27022 12964 27074
rect 12908 26964 12964 27022
rect 12908 26898 12964 26908
rect 13244 27748 13300 27758
rect 12124 26514 12180 26852
rect 12572 26850 12628 26862
rect 12572 26798 12574 26850
rect 12626 26798 12628 26850
rect 12124 26462 12126 26514
rect 12178 26462 12180 26514
rect 12124 26450 12180 26462
rect 12348 26516 12404 26526
rect 12572 26516 12628 26798
rect 12404 26460 12628 26516
rect 12348 26422 12404 26460
rect 12012 26402 12068 26414
rect 12012 26350 12014 26402
rect 12066 26350 12068 26402
rect 12012 25956 12068 26350
rect 12684 26402 12740 26414
rect 12684 26350 12686 26402
rect 12738 26350 12740 26402
rect 12684 26292 12740 26350
rect 12684 26226 12740 26236
rect 12012 25890 12068 25900
rect 13132 26178 13188 26190
rect 13132 26126 13134 26178
rect 13186 26126 13188 26178
rect 13132 25956 13188 26126
rect 13132 25890 13188 25900
rect 12012 23380 12068 23390
rect 12012 23286 12068 23324
rect 12348 23380 12404 23390
rect 12348 23286 12404 23324
rect 12684 23380 12740 23390
rect 12684 19906 12740 23324
rect 12684 19854 12686 19906
rect 12738 19854 12740 19906
rect 12684 19842 12740 19854
rect 11900 19516 12292 19572
rect 11676 18398 11678 18450
rect 11730 18398 11732 18450
rect 11676 18386 11732 18398
rect 11900 18452 11956 18462
rect 11900 18358 11956 18396
rect 11340 18228 11396 18238
rect 11228 18226 11396 18228
rect 11228 18174 11342 18226
rect 11394 18174 11396 18226
rect 11228 18172 11396 18174
rect 9100 16118 9156 16156
rect 9660 16100 9716 16110
rect 8876 15540 8932 15550
rect 8876 15446 8932 15484
rect 9660 15538 9716 16044
rect 10780 16100 10836 16110
rect 11340 16100 11396 18172
rect 11676 16884 11732 16894
rect 11676 16790 11732 16828
rect 12236 16212 12292 19516
rect 12348 18452 12404 18462
rect 12348 18358 12404 18396
rect 12348 16212 12404 16222
rect 12236 16210 12740 16212
rect 12236 16158 12350 16210
rect 12402 16158 12740 16210
rect 12236 16156 12740 16158
rect 12348 16146 12404 16156
rect 10780 16098 11396 16100
rect 10780 16046 10782 16098
rect 10834 16046 11396 16098
rect 10780 16044 11396 16046
rect 12684 16098 12740 16156
rect 12684 16046 12686 16098
rect 12738 16046 12740 16098
rect 10780 16034 10836 16044
rect 12684 16034 12740 16046
rect 13020 16100 13076 16110
rect 13020 16006 13076 16044
rect 9660 15486 9662 15538
rect 9714 15486 9716 15538
rect 9660 15474 9716 15486
rect 10444 15874 10500 15886
rect 10444 15822 10446 15874
rect 10498 15822 10500 15874
rect 9884 15428 9940 15438
rect 9884 15334 9940 15372
rect 9548 15316 9604 15326
rect 9548 15222 9604 15260
rect 9996 15314 10052 15326
rect 9996 15262 9998 15314
rect 10050 15262 10052 15314
rect 8764 15138 8820 15148
rect 9436 15204 9492 15214
rect 8764 12852 8820 12862
rect 8540 12740 8596 12750
rect 8540 12646 8596 12684
rect 8316 12180 8372 12190
rect 8428 12180 8484 12348
rect 8764 12290 8820 12796
rect 8764 12238 8766 12290
rect 8818 12238 8820 12290
rect 8316 12178 8484 12180
rect 8316 12126 8318 12178
rect 8370 12126 8484 12178
rect 8316 12124 8484 12126
rect 8652 12180 8708 12190
rect 8316 12114 8372 12124
rect 8652 12086 8708 12124
rect 8092 11956 8148 11966
rect 8092 11954 8372 11956
rect 8092 11902 8094 11954
rect 8146 11902 8372 11954
rect 8092 11900 8372 11902
rect 8092 11890 8148 11900
rect 8316 11508 8372 11900
rect 8428 11508 8484 11518
rect 8764 11508 8820 12238
rect 9100 12068 9156 12078
rect 8316 11506 8484 11508
rect 8316 11454 8430 11506
rect 8482 11454 8484 11506
rect 8316 11452 8484 11454
rect 8428 11442 8484 11452
rect 8540 11452 8820 11508
rect 8876 11508 8932 11518
rect 8428 11284 8484 11294
rect 8540 11284 8596 11452
rect 8428 11282 8596 11284
rect 8428 11230 8430 11282
rect 8482 11230 8596 11282
rect 8428 11228 8596 11230
rect 8428 11218 8484 11228
rect 8316 11172 8372 11182
rect 8316 11078 8372 11116
rect 8092 10948 8148 10958
rect 8148 10892 8372 10948
rect 8092 10882 8148 10892
rect 8316 10834 8372 10892
rect 8316 10782 8318 10834
rect 8370 10782 8372 10834
rect 8316 10770 8372 10782
rect 8540 10834 8596 11228
rect 8876 11394 8932 11452
rect 8876 11342 8878 11394
rect 8930 11342 8932 11394
rect 8876 11284 8932 11342
rect 8876 11218 8932 11228
rect 8540 10782 8542 10834
rect 8594 10782 8596 10834
rect 8540 10770 8596 10782
rect 8652 11170 8708 11182
rect 8652 11118 8654 11170
rect 8706 11118 8708 11170
rect 8652 11060 8708 11118
rect 9100 11060 9156 12012
rect 9324 11508 9380 11518
rect 9436 11508 9492 15148
rect 9996 14754 10052 15262
rect 9996 14702 9998 14754
rect 10050 14702 10052 14754
rect 9996 14690 10052 14702
rect 10220 15316 10276 15326
rect 10220 15148 10276 15260
rect 10444 15148 10500 15822
rect 12796 15874 12852 15886
rect 12796 15822 12798 15874
rect 12850 15822 12852 15874
rect 10220 15092 10500 15148
rect 12460 15764 12516 15774
rect 12460 15316 12516 15708
rect 9996 14530 10052 14542
rect 9996 14478 9998 14530
rect 10050 14478 10052 14530
rect 9660 14420 9716 14430
rect 9660 14326 9716 14364
rect 9996 14308 10052 14478
rect 9996 14242 10052 14252
rect 9660 12404 9716 12414
rect 9660 12310 9716 12348
rect 8652 11004 9156 11060
rect 9212 11452 9324 11508
rect 9380 11452 9492 11508
rect 8652 10834 8708 11004
rect 8652 10782 8654 10834
rect 8706 10782 8708 10834
rect 8652 10770 8708 10782
rect 9100 10836 9156 10846
rect 9212 10836 9268 11452
rect 9324 11414 9380 11452
rect 9100 10834 9268 10836
rect 9100 10782 9102 10834
rect 9154 10782 9268 10834
rect 9100 10780 9268 10782
rect 10220 11172 10276 15092
rect 11564 12740 11620 12750
rect 11564 12180 11620 12684
rect 12236 12292 12292 12302
rect 12236 12198 12292 12236
rect 9100 10770 9156 10780
rect 10220 10722 10276 11116
rect 10220 10670 10222 10722
rect 10274 10670 10276 10722
rect 10220 10658 10276 10670
rect 11340 12178 11620 12180
rect 11340 12126 11566 12178
rect 11618 12126 11620 12178
rect 11340 12124 11620 12126
rect 11340 11396 11396 12124
rect 11564 12114 11620 12124
rect 11900 12178 11956 12190
rect 11900 12126 11902 12178
rect 11954 12126 11956 12178
rect 11788 12066 11844 12078
rect 11788 12014 11790 12066
rect 11842 12014 11844 12066
rect 11788 11844 11844 12014
rect 8092 10612 8148 10622
rect 8092 10518 8148 10556
rect 10444 10612 10500 10622
rect 11228 10612 11284 10622
rect 10444 10610 11228 10612
rect 10444 10558 10446 10610
rect 10498 10558 11228 10610
rect 10444 10556 11228 10558
rect 10444 10546 10500 10556
rect 11228 10518 11284 10556
rect 11340 10610 11396 11340
rect 11676 11788 11844 11844
rect 11340 10558 11342 10610
rect 11394 10558 11396 10610
rect 11340 10546 11396 10558
rect 11564 10610 11620 10622
rect 11564 10558 11566 10610
rect 11618 10558 11620 10610
rect 11452 10498 11508 10510
rect 11452 10446 11454 10498
rect 11506 10446 11508 10498
rect 10780 10386 10836 10398
rect 10780 10334 10782 10386
rect 10834 10334 10836 10386
rect 10780 10052 10836 10334
rect 10780 9986 10836 9996
rect 7980 9762 8036 9772
rect 8092 9940 8148 9950
rect 7980 9604 8036 9614
rect 8092 9604 8148 9884
rect 7868 9602 8148 9604
rect 7868 9550 7982 9602
rect 8034 9550 8148 9602
rect 7868 9548 8148 9550
rect 7980 9538 8036 9548
rect 11452 9268 11508 10446
rect 11564 10052 11620 10558
rect 11676 10612 11732 11788
rect 11788 11284 11844 11294
rect 11900 11284 11956 12126
rect 11844 11228 11956 11284
rect 12236 11396 12292 11406
rect 11788 10722 11844 11228
rect 11788 10670 11790 10722
rect 11842 10670 11844 10722
rect 11788 10658 11844 10670
rect 11676 10546 11732 10556
rect 12236 10612 12292 11340
rect 12348 11284 12404 11294
rect 12348 11190 12404 11228
rect 12236 10546 12292 10556
rect 12460 10276 12516 15260
rect 12796 14308 12852 15822
rect 13244 15540 13300 27692
rect 13468 26964 13524 28700
rect 13692 27972 13748 27982
rect 13692 27878 13748 27916
rect 13580 27858 13636 27870
rect 13580 27806 13582 27858
rect 13634 27806 13636 27858
rect 13580 27300 13636 27806
rect 13580 27244 13860 27300
rect 13804 27186 13860 27244
rect 13804 27134 13806 27186
rect 13858 27134 13860 27186
rect 13804 27122 13860 27134
rect 13916 27074 13972 29934
rect 14700 29650 14756 30044
rect 14700 29598 14702 29650
rect 14754 29598 14756 29650
rect 14700 29586 14756 29598
rect 14252 29540 14308 29550
rect 14588 29540 14644 29550
rect 14252 29538 14588 29540
rect 14252 29486 14254 29538
rect 14306 29486 14588 29538
rect 14252 29484 14588 29486
rect 14252 29474 14308 29484
rect 14588 29446 14644 29484
rect 14364 28756 14420 28766
rect 14028 27858 14084 27870
rect 14028 27806 14030 27858
rect 14082 27806 14084 27858
rect 14028 27748 14084 27806
rect 14028 27682 14084 27692
rect 13916 27022 13918 27074
rect 13970 27022 13972 27074
rect 13916 27010 13972 27022
rect 14364 27074 14420 28700
rect 14924 28084 14980 30270
rect 14924 28018 14980 28028
rect 15036 29986 15092 31164
rect 15036 29934 15038 29986
rect 15090 29934 15092 29986
rect 14924 27860 14980 27870
rect 14924 27766 14980 27804
rect 15036 27634 15092 29934
rect 15148 29540 15204 32844
rect 15484 32788 15540 32844
rect 15484 32694 15540 32732
rect 15708 31948 15764 34078
rect 15932 34130 15988 34142
rect 15932 34078 15934 34130
rect 15986 34078 15988 34130
rect 15932 34020 15988 34078
rect 15932 33954 15988 33964
rect 16380 34020 16436 34030
rect 16380 33926 16436 33964
rect 15820 33348 15876 33358
rect 15820 32676 15876 33292
rect 17276 33236 17332 33246
rect 17052 33124 17108 33134
rect 17052 33030 17108 33068
rect 16380 32788 16436 32798
rect 16436 32732 16548 32788
rect 16380 32722 16436 32732
rect 15820 32582 15876 32620
rect 16044 32564 16100 32574
rect 16044 32470 16100 32508
rect 16492 32562 16548 32732
rect 16492 32510 16494 32562
rect 16546 32510 16548 32562
rect 16492 32498 16548 32510
rect 16716 32676 16772 32686
rect 16268 32340 16324 32350
rect 16268 32246 16324 32284
rect 15708 31892 16212 31948
rect 15484 31780 15540 31790
rect 15260 30098 15316 30110
rect 15260 30046 15262 30098
rect 15314 30046 15316 30098
rect 15260 29876 15316 30046
rect 15484 29876 15540 31724
rect 15596 31778 15652 31790
rect 15596 31726 15598 31778
rect 15650 31726 15652 31778
rect 15596 30996 15652 31726
rect 15820 30996 15876 31006
rect 15596 30994 15876 30996
rect 15596 30942 15822 30994
rect 15874 30942 15876 30994
rect 15596 30940 15876 30942
rect 15820 30884 15876 30940
rect 15820 30818 15876 30828
rect 16044 30212 16100 30222
rect 16044 30118 16100 30156
rect 15596 30100 15652 30110
rect 15596 30006 15652 30044
rect 15820 29986 15876 29998
rect 15820 29934 15822 29986
rect 15874 29934 15876 29986
rect 15260 29820 15764 29876
rect 15148 29092 15204 29484
rect 15260 29428 15316 29438
rect 15260 29426 15540 29428
rect 15260 29374 15262 29426
rect 15314 29374 15540 29426
rect 15260 29372 15540 29374
rect 15260 29362 15316 29372
rect 15148 29036 15428 29092
rect 15260 28642 15316 28654
rect 15260 28590 15262 28642
rect 15314 28590 15316 28642
rect 15260 27860 15316 28590
rect 15260 27794 15316 27804
rect 15372 27972 15428 29036
rect 15484 28866 15540 29372
rect 15708 29202 15764 29820
rect 15708 29150 15710 29202
rect 15762 29150 15764 29202
rect 15708 29138 15764 29150
rect 15484 28814 15486 28866
rect 15538 28814 15540 28866
rect 15484 28802 15540 28814
rect 15820 28756 15876 29934
rect 15932 29986 15988 29998
rect 15932 29934 15934 29986
rect 15986 29934 15988 29986
rect 15932 29426 15988 29934
rect 16156 29988 16212 31892
rect 16380 30884 16436 30894
rect 16380 30790 16436 30828
rect 16268 30212 16324 30222
rect 16268 30210 16660 30212
rect 16268 30158 16270 30210
rect 16322 30158 16660 30210
rect 16268 30156 16660 30158
rect 16268 30146 16324 30156
rect 16492 29988 16548 29998
rect 16156 29932 16436 29988
rect 16268 29764 16324 29774
rect 15932 29374 15934 29426
rect 15986 29374 15988 29426
rect 15932 29362 15988 29374
rect 16156 29708 16268 29764
rect 15596 28700 15876 28756
rect 16156 28756 16212 29708
rect 16268 29698 16324 29708
rect 16268 29538 16324 29550
rect 16268 29486 16270 29538
rect 16322 29486 16324 29538
rect 16268 28756 16324 29486
rect 16380 29204 16436 29932
rect 16492 29426 16548 29932
rect 16492 29374 16494 29426
rect 16546 29374 16548 29426
rect 16492 29362 16548 29374
rect 16380 29148 16548 29204
rect 16268 28700 16436 28756
rect 15484 28644 15540 28654
rect 15484 28550 15540 28588
rect 15036 27582 15038 27634
rect 15090 27582 15092 27634
rect 15036 27570 15092 27582
rect 15372 27186 15428 27916
rect 15372 27134 15374 27186
rect 15426 27134 15428 27186
rect 15372 27122 15428 27134
rect 14364 27022 14366 27074
rect 14418 27022 14420 27074
rect 14364 27010 14420 27022
rect 13804 26964 13860 26974
rect 13356 26962 13860 26964
rect 13356 26910 13806 26962
rect 13858 26910 13860 26962
rect 13356 26908 13860 26910
rect 13356 23380 13412 26908
rect 13804 26898 13860 26908
rect 14140 26852 14196 26862
rect 14140 26758 14196 26796
rect 15372 26852 15428 26862
rect 13692 26740 13748 26750
rect 13748 26684 13860 26740
rect 13692 26674 13748 26684
rect 13580 24388 13636 24398
rect 13580 23828 13636 24332
rect 13804 24162 13860 26684
rect 15372 26514 15428 26796
rect 15596 26628 15652 28700
rect 16156 28644 16212 28700
rect 16156 28588 16324 28644
rect 15820 28532 15876 28542
rect 15820 28438 15876 28476
rect 16268 28530 16324 28588
rect 16268 28478 16270 28530
rect 16322 28478 16324 28530
rect 16268 28466 16324 28478
rect 16156 28420 16212 28430
rect 15932 28418 16212 28420
rect 15932 28366 16158 28418
rect 16210 28366 16212 28418
rect 15932 28364 16212 28366
rect 15820 28084 15876 28094
rect 15932 28084 15988 28364
rect 16156 28354 16212 28364
rect 15820 28082 15988 28084
rect 15820 28030 15822 28082
rect 15874 28030 15988 28082
rect 15820 28028 15988 28030
rect 16044 28140 16324 28196
rect 16044 28082 16100 28140
rect 16044 28030 16046 28082
rect 16098 28030 16100 28082
rect 15820 28018 15876 28028
rect 16044 28018 16100 28030
rect 16156 27972 16212 27982
rect 15596 26562 15652 26572
rect 15708 27858 15764 27870
rect 15708 27806 15710 27858
rect 15762 27806 15764 27858
rect 15372 26462 15374 26514
rect 15426 26462 15428 26514
rect 15372 24724 15428 26462
rect 15484 26292 15540 26302
rect 15708 26292 15764 27806
rect 15484 26290 15764 26292
rect 15484 26238 15486 26290
rect 15538 26238 15764 26290
rect 15484 26236 15764 26238
rect 15484 26226 15540 26236
rect 15596 24724 15652 24734
rect 15372 24722 15652 24724
rect 15372 24670 15598 24722
rect 15650 24670 15652 24722
rect 15372 24668 15652 24670
rect 15596 24658 15652 24668
rect 13804 24110 13806 24162
rect 13858 24110 13860 24162
rect 13804 24098 13860 24110
rect 14252 24388 14308 24398
rect 14252 24050 14308 24332
rect 14252 23998 14254 24050
rect 14306 23998 14308 24050
rect 14252 23986 14308 23998
rect 15708 23940 15764 26236
rect 13356 23314 13412 23324
rect 13468 23826 13636 23828
rect 13468 23774 13582 23826
rect 13634 23774 13636 23826
rect 13468 23772 13636 23774
rect 13244 15474 13300 15484
rect 13468 18452 13524 23772
rect 13580 23762 13636 23772
rect 15484 23884 15708 23940
rect 13692 23714 13748 23726
rect 13692 23662 13694 23714
rect 13746 23662 13748 23714
rect 13692 23044 13748 23662
rect 13692 21924 13748 22988
rect 13692 21858 13748 21868
rect 14588 21924 14644 21934
rect 14364 20914 14420 20926
rect 14364 20862 14366 20914
rect 14418 20862 14420 20914
rect 13132 15316 13188 15326
rect 13132 15202 13188 15260
rect 13132 15150 13134 15202
rect 13186 15150 13188 15202
rect 13132 15138 13188 15150
rect 12796 14242 12852 14252
rect 13468 14306 13524 18396
rect 13468 14254 13470 14306
rect 13522 14254 13524 14306
rect 13468 13412 13524 14254
rect 12796 12292 12852 12302
rect 12796 12198 12852 12236
rect 13468 12292 13524 13356
rect 13468 12226 13524 12236
rect 13580 20578 13636 20590
rect 13580 20526 13582 20578
rect 13634 20526 13636 20578
rect 13580 19908 13636 20526
rect 13804 20580 13860 20590
rect 13692 20020 13748 20030
rect 13692 19926 13748 19964
rect 13580 16994 13636 19852
rect 13804 19122 13860 20524
rect 14364 20130 14420 20862
rect 14588 20804 14644 21868
rect 15484 21810 15540 23884
rect 15708 23874 15764 23884
rect 15820 27860 15876 27870
rect 16044 27860 16100 27870
rect 15484 21758 15486 21810
rect 15538 21758 15540 21810
rect 15484 21746 15540 21758
rect 15260 21588 15316 21598
rect 15260 21494 15316 21532
rect 15708 21586 15764 21598
rect 15708 21534 15710 21586
rect 15762 21534 15764 21586
rect 14700 21476 14756 21486
rect 14700 21026 14756 21420
rect 15596 21476 15652 21486
rect 15596 21382 15652 21420
rect 14700 20974 14702 21026
rect 14754 20974 14756 21026
rect 14700 20962 14756 20974
rect 14588 20748 14756 20804
rect 14476 20580 14532 20590
rect 14476 20486 14532 20524
rect 14364 20078 14366 20130
rect 14418 20078 14420 20130
rect 14364 20066 14420 20078
rect 13804 19070 13806 19122
rect 13858 19070 13860 19122
rect 13804 19058 13860 19070
rect 13580 16942 13582 16994
rect 13634 16942 13636 16994
rect 13468 11284 13524 11294
rect 12572 11170 12628 11182
rect 12572 11118 12574 11170
rect 12626 11118 12628 11170
rect 12572 10610 12628 11118
rect 12572 10558 12574 10610
rect 12626 10558 12628 10610
rect 12572 10546 12628 10558
rect 12684 10724 12740 10734
rect 12684 10610 12740 10668
rect 12684 10558 12686 10610
rect 12738 10558 12740 10610
rect 12684 10546 12740 10558
rect 12908 10386 12964 10398
rect 12908 10334 12910 10386
rect 12962 10334 12964 10386
rect 12460 10220 12628 10276
rect 11564 9986 11620 9996
rect 12124 10052 12180 10062
rect 12124 9826 12180 9996
rect 12124 9774 12126 9826
rect 12178 9774 12180 9826
rect 12124 9762 12180 9774
rect 12460 10052 12516 10062
rect 12460 9826 12516 9996
rect 12460 9774 12462 9826
rect 12514 9774 12516 9826
rect 12460 9762 12516 9774
rect 11116 9212 11508 9268
rect 12348 9602 12404 9614
rect 12348 9550 12350 9602
rect 12402 9550 12404 9602
rect 7084 9044 7140 9054
rect 7084 8950 7140 8988
rect 6636 8930 6804 8932
rect 6636 8878 6638 8930
rect 6690 8878 6804 8930
rect 6636 8876 6804 8878
rect 6636 8866 6692 8876
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 10780 8370 10836 8382
rect 10780 8318 10782 8370
rect 10834 8318 10836 8370
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 10668 6804 10724 6814
rect 10780 6804 10836 8318
rect 10892 8372 10948 8382
rect 10892 8146 10948 8316
rect 11116 8370 11172 9212
rect 12348 8482 12404 9550
rect 12348 8430 12350 8482
rect 12402 8430 12404 8482
rect 12348 8418 12404 8430
rect 11116 8318 11118 8370
rect 11170 8318 11172 8370
rect 11116 8306 11172 8318
rect 11564 8372 11620 8382
rect 11564 8278 11620 8316
rect 12572 8372 12628 10220
rect 12908 10052 12964 10334
rect 12908 9986 12964 9996
rect 13020 10386 13076 10398
rect 13020 10334 13022 10386
rect 13074 10334 13076 10386
rect 12796 9828 12852 9838
rect 13020 9828 13076 10334
rect 12796 9826 13076 9828
rect 12796 9774 12798 9826
rect 12850 9774 13076 9826
rect 12796 9772 13076 9774
rect 12796 9762 12852 9772
rect 13468 9714 13524 11228
rect 13468 9662 13470 9714
rect 13522 9662 13524 9714
rect 13468 9650 13524 9662
rect 12796 9604 12852 9614
rect 10892 8094 10894 8146
rect 10946 8094 10948 8146
rect 10892 8082 10948 8094
rect 12572 8146 12628 8316
rect 12572 8094 12574 8146
rect 12626 8094 12628 8146
rect 12572 8036 12628 8094
rect 12572 7970 12628 7980
rect 12684 8370 12740 8382
rect 12684 8318 12686 8370
rect 12738 8318 12740 8370
rect 10668 6802 10836 6804
rect 10668 6750 10670 6802
rect 10722 6750 10836 6802
rect 10668 6748 10836 6750
rect 10668 6738 10724 6748
rect 9996 6692 10052 6702
rect 9996 6598 10052 6636
rect 12124 6692 12180 6702
rect 12124 5906 12180 6636
rect 12684 6020 12740 8318
rect 12796 6802 12852 9548
rect 13580 8260 13636 16942
rect 14140 19012 14196 19022
rect 14588 19012 14644 19022
rect 14140 19010 14644 19012
rect 14140 18958 14142 19010
rect 14194 18958 14590 19010
rect 14642 18958 14644 19010
rect 14140 18956 14644 18958
rect 14140 18564 14196 18956
rect 14588 18946 14644 18956
rect 14028 15428 14084 15438
rect 14028 15334 14084 15372
rect 13692 15316 13748 15326
rect 13692 15314 13972 15316
rect 13692 15262 13694 15314
rect 13746 15262 13972 15314
rect 13692 15260 13972 15262
rect 13692 15250 13748 15260
rect 13916 15204 13972 15260
rect 14140 15204 14196 18508
rect 14588 18452 14644 18462
rect 14700 18452 14756 20748
rect 15708 20188 15764 21534
rect 15820 21476 15876 27804
rect 15932 27804 16044 27860
rect 15932 27746 15988 27804
rect 16044 27794 16100 27804
rect 16156 27858 16212 27916
rect 16156 27806 16158 27858
rect 16210 27806 16212 27858
rect 16156 27794 16212 27806
rect 15932 27694 15934 27746
rect 15986 27694 15988 27746
rect 15932 27682 15988 27694
rect 16268 26516 16324 28140
rect 16380 27860 16436 28700
rect 16380 27794 16436 27804
rect 16268 26450 16324 26460
rect 16268 26290 16324 26302
rect 16268 26238 16270 26290
rect 16322 26238 16324 26290
rect 16044 24722 16100 24734
rect 16044 24670 16046 24722
rect 16098 24670 16100 24722
rect 16044 23380 16100 24670
rect 16268 24612 16324 26238
rect 16492 26178 16548 29148
rect 16604 28866 16660 30156
rect 16716 29764 16772 32620
rect 17276 32562 17332 33180
rect 17612 33124 17668 33134
rect 17612 32786 17668 33068
rect 17612 32734 17614 32786
rect 17666 32734 17668 32786
rect 17612 32722 17668 32734
rect 17276 32510 17278 32562
rect 17330 32510 17332 32562
rect 17276 32498 17332 32510
rect 17836 32674 17892 32686
rect 17836 32622 17838 32674
rect 17890 32622 17892 32674
rect 17836 32564 17892 32622
rect 16940 32338 16996 32350
rect 16940 32286 16942 32338
rect 16994 32286 16996 32338
rect 16940 30996 16996 32286
rect 16940 30930 16996 30940
rect 16716 29698 16772 29708
rect 16604 28814 16606 28866
rect 16658 28814 16660 28866
rect 16604 28802 16660 28814
rect 16716 28868 16772 28878
rect 16716 28756 16772 28812
rect 17164 28756 17220 28766
rect 16716 28754 17220 28756
rect 16716 28702 16718 28754
rect 16770 28702 17166 28754
rect 17218 28702 17220 28754
rect 16716 28700 17220 28702
rect 16716 28690 16772 28700
rect 16828 26404 16884 26414
rect 16828 26310 16884 26348
rect 16604 26292 16660 26302
rect 16604 26198 16660 26236
rect 16492 26126 16494 26178
rect 16546 26126 16548 26178
rect 16492 26114 16548 26126
rect 16044 23314 16100 23324
rect 16156 24610 16324 24612
rect 16156 24558 16270 24610
rect 16322 24558 16324 24610
rect 16156 24556 16324 24558
rect 15932 21700 15988 21710
rect 16156 21700 16212 24556
rect 16268 24546 16324 24556
rect 16716 25396 16772 25406
rect 16268 24052 16324 24062
rect 16268 23958 16324 23996
rect 15932 21698 16212 21700
rect 15932 21646 15934 21698
rect 15986 21646 16212 21698
rect 15932 21644 16212 21646
rect 16492 23940 16548 23950
rect 15932 21634 15988 21644
rect 15820 21420 16212 21476
rect 16044 20244 16100 20254
rect 15708 20132 16100 20188
rect 16156 20188 16212 21420
rect 16156 20132 16324 20188
rect 14588 18450 14756 18452
rect 14588 18398 14590 18450
rect 14642 18398 14756 18450
rect 14588 18396 14756 18398
rect 14812 18562 14868 18574
rect 14812 18510 14814 18562
rect 14866 18510 14868 18562
rect 14588 18386 14644 18396
rect 14812 17444 14868 18510
rect 14812 17378 14868 17388
rect 15708 17444 15764 20132
rect 15708 17378 15764 17388
rect 15484 16884 15540 16894
rect 15484 16098 15540 16828
rect 15484 16046 15486 16098
rect 15538 16046 15540 16098
rect 15484 16034 15540 16046
rect 15932 16660 15988 16670
rect 14364 15876 14420 15886
rect 14364 15538 14420 15820
rect 14364 15486 14366 15538
rect 14418 15486 14420 15538
rect 14364 15474 14420 15486
rect 14812 15204 14868 15214
rect 13916 15202 14868 15204
rect 13916 15150 14814 15202
rect 14866 15150 14868 15202
rect 13916 15148 14868 15150
rect 14812 15138 14868 15148
rect 15260 14644 15316 14654
rect 15260 14530 15316 14588
rect 15932 14642 15988 16604
rect 15932 14590 15934 14642
rect 15986 14590 15988 14642
rect 15932 14578 15988 14590
rect 16044 15876 16100 15886
rect 15260 14478 15262 14530
rect 15314 14478 15316 14530
rect 15260 14466 15316 14478
rect 13804 14308 13860 14318
rect 13860 14252 13972 14308
rect 13804 14214 13860 14252
rect 13804 11956 13860 11966
rect 13804 11618 13860 11900
rect 13804 11566 13806 11618
rect 13858 11566 13860 11618
rect 13804 11554 13860 11566
rect 13692 11284 13748 11294
rect 13916 11284 13972 14252
rect 14252 14306 14308 14318
rect 14252 14254 14254 14306
rect 14306 14254 14308 14306
rect 14252 13412 14308 14254
rect 14252 13346 14308 13356
rect 16044 12402 16100 15820
rect 16044 12350 16046 12402
rect 16098 12350 16100 12402
rect 16044 12338 16100 12350
rect 15932 12178 15988 12190
rect 15932 12126 15934 12178
rect 15986 12126 15988 12178
rect 14812 12068 14868 12078
rect 14812 11974 14868 12012
rect 15036 11956 15092 11966
rect 15036 11862 15092 11900
rect 15260 11954 15316 11966
rect 15260 11902 15262 11954
rect 15314 11902 15316 11954
rect 15260 11732 15316 11902
rect 15260 11666 15316 11676
rect 15708 11954 15764 11966
rect 15708 11902 15710 11954
rect 15762 11902 15764 11954
rect 15708 11396 15764 11902
rect 15708 11330 15764 11340
rect 13916 11228 14084 11284
rect 13692 11190 13748 11228
rect 13804 11172 13860 11182
rect 13804 11170 13972 11172
rect 13804 11118 13806 11170
rect 13858 11118 13972 11170
rect 13804 11116 13972 11118
rect 13804 11106 13860 11116
rect 13804 10612 13860 10622
rect 13916 10612 13972 11116
rect 14028 10836 14084 11228
rect 15932 11060 15988 12126
rect 16044 11954 16100 11966
rect 16044 11902 16046 11954
rect 16098 11902 16100 11954
rect 16044 11732 16100 11902
rect 16044 11666 16100 11676
rect 14028 10770 14084 10780
rect 15708 11004 15988 11060
rect 15148 10722 15204 10734
rect 15148 10670 15150 10722
rect 15202 10670 15204 10722
rect 14364 10612 14420 10622
rect 13916 10610 14420 10612
rect 13916 10558 14366 10610
rect 14418 10558 14420 10610
rect 13916 10556 14420 10558
rect 13804 10518 13860 10556
rect 14364 10052 14420 10556
rect 15148 10388 15204 10670
rect 15260 10612 15316 10622
rect 15260 10518 15316 10556
rect 15708 10610 15764 11004
rect 15932 10724 15988 10734
rect 15932 10630 15988 10668
rect 15708 10558 15710 10610
rect 15762 10558 15764 10610
rect 13692 9826 13748 9838
rect 13692 9774 13694 9826
rect 13746 9774 13748 9826
rect 13692 9604 13748 9774
rect 13692 9538 13748 9548
rect 14252 9268 14308 9278
rect 14364 9268 14420 9996
rect 14588 10332 15204 10388
rect 15372 10388 15428 10398
rect 15708 10388 15764 10558
rect 15372 10386 15764 10388
rect 15372 10334 15374 10386
rect 15426 10334 15764 10386
rect 15372 10332 15764 10334
rect 15820 10498 15876 10510
rect 15820 10446 15822 10498
rect 15874 10446 15876 10498
rect 14252 9266 14420 9268
rect 14252 9214 14254 9266
rect 14306 9214 14420 9266
rect 14252 9212 14420 9214
rect 14476 9826 14532 9838
rect 14476 9774 14478 9826
rect 14530 9774 14532 9826
rect 14252 9202 14308 9212
rect 14476 9044 14532 9774
rect 14588 9714 14644 10332
rect 15372 10322 15428 10332
rect 15820 10052 15876 10446
rect 15820 9986 15876 9996
rect 16268 9938 16324 20132
rect 16492 19906 16548 23884
rect 16716 23938 16772 25340
rect 17164 25172 17220 28700
rect 17836 27076 17892 32508
rect 17948 32338 18004 32350
rect 17948 32286 17950 32338
rect 18002 32286 18004 32338
rect 17948 30324 18004 32286
rect 17948 30258 18004 30268
rect 18284 31890 18340 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 18284 31838 18286 31890
rect 18338 31838 18340 31890
rect 18284 28756 18340 31838
rect 18508 34020 18564 34030
rect 18284 28690 18340 28700
rect 18396 29986 18452 29998
rect 18396 29934 18398 29986
rect 18450 29934 18452 29986
rect 17836 27010 17892 27020
rect 17276 26628 17332 26638
rect 17276 25396 17332 26572
rect 17388 26516 17444 26526
rect 17388 26422 17444 26460
rect 17948 26404 18004 26414
rect 17948 26310 18004 26348
rect 17276 25302 17332 25340
rect 17500 26178 17556 26190
rect 17500 26126 17502 26178
rect 17554 26126 17556 26178
rect 17500 25284 17556 26126
rect 18060 25396 18116 25406
rect 17612 25284 17668 25294
rect 17500 25282 17668 25284
rect 17500 25230 17614 25282
rect 17666 25230 17668 25282
rect 17500 25228 17668 25230
rect 16716 23886 16718 23938
rect 16770 23886 16772 23938
rect 16716 23874 16772 23886
rect 16940 25116 17220 25172
rect 16940 23938 16996 25116
rect 16940 23886 16942 23938
rect 16994 23886 16996 23938
rect 16940 23492 16996 23886
rect 17164 23938 17220 23950
rect 17164 23886 17166 23938
rect 17218 23886 17220 23938
rect 17164 23604 17220 23886
rect 17276 23940 17332 23950
rect 17276 23846 17332 23884
rect 17164 23548 17556 23604
rect 16940 23426 16996 23436
rect 17388 23380 17444 23390
rect 17388 23286 17444 23324
rect 17500 23268 17556 23548
rect 17500 23174 17556 23212
rect 17612 23044 17668 25228
rect 17724 23714 17780 23726
rect 17724 23662 17726 23714
rect 17778 23662 17780 23714
rect 17724 23492 17780 23662
rect 17724 23426 17780 23436
rect 17724 23156 17780 23166
rect 17948 23156 18004 23166
rect 17724 23062 17780 23100
rect 17836 23154 18004 23156
rect 17836 23102 17950 23154
rect 18002 23102 18004 23154
rect 17836 23100 18004 23102
rect 17500 22988 17668 23044
rect 17500 21812 17556 22988
rect 17500 21746 17556 21756
rect 17612 22148 17668 22158
rect 17836 22148 17892 23100
rect 17948 23090 18004 23100
rect 18060 22932 18116 25340
rect 18396 24388 18452 29934
rect 18508 27972 18564 33964
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20412 32900 20468 32910
rect 20300 32788 20356 32798
rect 20300 32694 20356 32732
rect 19404 32450 19460 32462
rect 19404 32398 19406 32450
rect 19458 32398 19460 32450
rect 19404 31668 19460 32398
rect 19628 32338 19684 32350
rect 19628 32286 19630 32338
rect 19682 32286 19684 32338
rect 19068 31556 19124 31566
rect 18956 31218 19012 31230
rect 18956 31166 18958 31218
rect 19010 31166 19012 31218
rect 18956 30660 19012 31166
rect 19068 30996 19124 31500
rect 19292 30996 19348 31006
rect 19068 30994 19236 30996
rect 19068 30942 19070 30994
rect 19122 30942 19236 30994
rect 19068 30940 19236 30942
rect 19068 30930 19124 30940
rect 18508 27906 18564 27916
rect 18620 30324 18676 30334
rect 18844 30324 18900 30334
rect 18620 27860 18676 30268
rect 18732 30268 18844 30324
rect 18732 30210 18788 30268
rect 18844 30258 18900 30268
rect 18732 30158 18734 30210
rect 18786 30158 18788 30210
rect 18732 30146 18788 30158
rect 18956 27972 19012 30604
rect 19180 30434 19236 30940
rect 19180 30382 19182 30434
rect 19234 30382 19236 30434
rect 19180 30370 19236 30382
rect 19292 30436 19348 30940
rect 19404 30772 19460 31612
rect 19516 32228 19572 32238
rect 19516 30996 19572 32172
rect 19628 31892 19684 32286
rect 19628 31220 19684 31836
rect 19852 32338 19908 32350
rect 19852 32286 19854 32338
rect 19906 32286 19908 32338
rect 19852 31780 19908 32286
rect 20076 31892 20132 31902
rect 20076 31798 20132 31836
rect 20412 31890 20468 32844
rect 20412 31838 20414 31890
rect 20466 31838 20468 31890
rect 20412 31826 20468 31838
rect 20524 31892 20580 36316
rect 21420 35138 21476 37884
rect 23660 37940 23716 37950
rect 23772 37940 23828 38780
rect 23660 37938 23828 37940
rect 23660 37886 23662 37938
rect 23714 37886 23828 37938
rect 23660 37884 23828 37886
rect 23884 38722 23940 40572
rect 24332 40562 24388 40572
rect 23884 38670 23886 38722
rect 23938 38670 23940 38722
rect 23660 37874 23716 37884
rect 23436 37826 23492 37838
rect 23436 37774 23438 37826
rect 23490 37774 23492 37826
rect 21644 36484 21700 36494
rect 21644 36390 21700 36428
rect 21868 36482 21924 36494
rect 21868 36430 21870 36482
rect 21922 36430 21924 36482
rect 21868 36260 21924 36430
rect 21868 35364 21924 36204
rect 23436 36484 23492 37774
rect 23884 37492 23940 38670
rect 24108 40402 24164 40414
rect 24108 40350 24110 40402
rect 24162 40350 24164 40402
rect 24108 38948 24164 40350
rect 25788 40404 25844 40414
rect 24220 40292 24276 40302
rect 24220 40198 24276 40236
rect 25452 40290 25508 40302
rect 25452 40238 25454 40290
rect 25506 40238 25508 40290
rect 24780 39060 24836 39070
rect 24780 38966 24836 39004
rect 25452 39060 25508 40238
rect 25676 40292 25732 40302
rect 25676 39730 25732 40236
rect 25676 39678 25678 39730
rect 25730 39678 25732 39730
rect 25676 39666 25732 39678
rect 25452 39004 25732 39060
rect 24444 38948 24500 38958
rect 24108 38946 24500 38948
rect 24108 38894 24110 38946
rect 24162 38894 24446 38946
rect 24498 38894 24500 38946
rect 24108 38892 24500 38894
rect 24108 38050 24164 38892
rect 24108 37998 24110 38050
rect 24162 37998 24164 38050
rect 24108 37986 24164 37998
rect 24220 38276 24276 38286
rect 24220 38050 24276 38220
rect 24444 38274 24500 38892
rect 24556 38948 24612 38958
rect 24556 38854 24612 38892
rect 24444 38222 24446 38274
rect 24498 38222 24500 38274
rect 24444 38210 24500 38222
rect 25452 38276 25508 39004
rect 25452 38210 25508 38220
rect 25564 38834 25620 38846
rect 25564 38782 25566 38834
rect 25618 38782 25620 38834
rect 25564 38274 25620 38782
rect 25676 38836 25732 39004
rect 25788 39058 25844 40348
rect 27804 40402 27860 40414
rect 27804 40350 27806 40402
rect 27858 40350 27860 40402
rect 26460 39620 26516 39630
rect 26460 39526 26516 39564
rect 26908 39620 26964 39630
rect 26908 39526 26964 39564
rect 27804 39620 27860 40350
rect 28476 40404 28532 40414
rect 28476 40310 28532 40348
rect 30604 40290 30660 41916
rect 30828 41906 30884 41916
rect 32620 41970 32676 41982
rect 36316 41972 36372 41982
rect 32620 41918 32622 41970
rect 32674 41918 32676 41970
rect 30604 40238 30606 40290
rect 30658 40238 30660 40290
rect 30604 40226 30660 40238
rect 31164 40404 31220 40414
rect 27804 39554 27860 39564
rect 29820 39620 29876 39630
rect 25788 39006 25790 39058
rect 25842 39006 25844 39058
rect 25788 38994 25844 39006
rect 26460 39396 26516 39406
rect 26460 39058 26516 39340
rect 26460 39006 26462 39058
rect 26514 39006 26516 39058
rect 26460 38994 26516 39006
rect 27132 39396 27188 39406
rect 27132 38946 27188 39340
rect 27132 38894 27134 38946
rect 27186 38894 27188 38946
rect 27132 38882 27188 38894
rect 25788 38836 25844 38846
rect 25676 38834 25844 38836
rect 25676 38782 25790 38834
rect 25842 38782 25844 38834
rect 25676 38780 25844 38782
rect 25788 38770 25844 38780
rect 26124 38836 26180 38846
rect 26124 38742 26180 38780
rect 26684 38834 26740 38846
rect 26684 38782 26686 38834
rect 26738 38782 26740 38834
rect 25564 38222 25566 38274
rect 25618 38222 25620 38274
rect 24220 37998 24222 38050
rect 24274 37998 24276 38050
rect 23884 37426 23940 37436
rect 24108 37492 24164 37502
rect 24220 37492 24276 37998
rect 24108 37490 24276 37492
rect 24108 37438 24110 37490
rect 24162 37438 24276 37490
rect 24108 37436 24276 37438
rect 25228 37492 25284 37502
rect 24108 37426 24164 37436
rect 25228 37398 25284 37436
rect 21868 35298 21924 35308
rect 22988 35364 23044 35374
rect 21420 35086 21422 35138
rect 21474 35086 21476 35138
rect 21420 35074 21476 35086
rect 20636 35028 20692 35038
rect 20636 35026 21364 35028
rect 20636 34974 20638 35026
rect 20690 34974 21364 35026
rect 20636 34972 21364 34974
rect 20636 34962 20692 34972
rect 21308 34914 21364 34972
rect 21308 34862 21310 34914
rect 21362 34862 21364 34914
rect 21308 34850 21364 34862
rect 20748 34802 20804 34814
rect 20748 34750 20750 34802
rect 20802 34750 20804 34802
rect 20636 34692 20692 34702
rect 20636 34132 20692 34636
rect 20748 34132 20804 34750
rect 21420 34692 21476 34702
rect 21420 34690 21588 34692
rect 21420 34638 21422 34690
rect 21474 34638 21588 34690
rect 21420 34636 21588 34638
rect 21420 34626 21476 34636
rect 21084 34132 21140 34142
rect 20748 34130 21140 34132
rect 20748 34078 21086 34130
rect 21138 34078 21140 34130
rect 20748 34076 21140 34078
rect 20636 34038 20692 34076
rect 21084 33572 21140 34076
rect 21084 32788 21140 33516
rect 21532 32788 21588 34636
rect 22764 34244 22820 34254
rect 22204 34130 22260 34142
rect 22204 34078 22206 34130
rect 22258 34078 22260 34130
rect 22204 33572 22260 34078
rect 22764 34130 22820 34188
rect 22764 34078 22766 34130
rect 22818 34078 22820 34130
rect 22764 34066 22820 34078
rect 22260 33516 22484 33572
rect 22204 33506 22260 33516
rect 21756 32788 21812 32798
rect 21532 32786 21812 32788
rect 21532 32734 21758 32786
rect 21810 32734 21812 32786
rect 21532 32732 21812 32734
rect 21084 32722 21140 32732
rect 21756 32722 21812 32732
rect 22204 32564 22260 32574
rect 22204 32470 22260 32508
rect 22428 32562 22484 33516
rect 22428 32510 22430 32562
rect 22482 32510 22484 32562
rect 22428 32498 22484 32510
rect 22652 32452 22708 32462
rect 22652 32358 22708 32396
rect 20636 31892 20692 31902
rect 20524 31890 20692 31892
rect 20524 31838 20638 31890
rect 20690 31838 20692 31890
rect 20524 31836 20692 31838
rect 20636 31826 20692 31836
rect 19852 31686 19908 31724
rect 20412 31668 20468 31678
rect 20412 31574 20468 31612
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19628 31154 19684 31164
rect 19516 30994 19796 30996
rect 19516 30942 19518 30994
rect 19570 30942 19796 30994
rect 19516 30940 19796 30942
rect 19516 30930 19572 30940
rect 19404 30716 19572 30772
rect 19404 30436 19460 30446
rect 19292 30434 19460 30436
rect 19292 30382 19406 30434
rect 19458 30382 19460 30434
rect 19292 30380 19460 30382
rect 19404 30370 19460 30380
rect 19516 30324 19572 30716
rect 19516 30212 19572 30268
rect 19628 30212 19684 30222
rect 19516 30210 19684 30212
rect 19516 30158 19630 30210
rect 19682 30158 19684 30210
rect 19516 30156 19684 30158
rect 19628 30146 19684 30156
rect 19740 30210 19796 30940
rect 20636 30884 20692 30894
rect 20636 30790 20692 30828
rect 19964 30324 20020 30334
rect 19964 30322 20244 30324
rect 19964 30270 19966 30322
rect 20018 30270 20244 30322
rect 19964 30268 20244 30270
rect 19964 30258 20020 30268
rect 19740 30158 19742 30210
rect 19794 30158 19796 30210
rect 19740 30146 19796 30158
rect 20188 29988 20244 30268
rect 20412 29988 20468 29998
rect 20188 29986 20468 29988
rect 20188 29934 20414 29986
rect 20466 29934 20468 29986
rect 20188 29932 20468 29934
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20412 29316 20468 29932
rect 20412 29250 20468 29260
rect 19404 28756 19460 28766
rect 19460 28700 19684 28756
rect 19404 28662 19460 28700
rect 18844 27916 19012 27972
rect 19292 27972 19348 27982
rect 18732 27860 18788 27870
rect 18620 27858 18788 27860
rect 18620 27806 18734 27858
rect 18786 27806 18788 27858
rect 18620 27804 18788 27806
rect 18732 27794 18788 27804
rect 18732 26404 18788 26414
rect 18732 26310 18788 26348
rect 18844 26068 18900 27916
rect 19068 27858 19124 27870
rect 19068 27806 19070 27858
rect 19122 27806 19124 27858
rect 18956 27748 19012 27758
rect 18956 27654 19012 27692
rect 18956 26292 19012 26302
rect 18956 26198 19012 26236
rect 19068 26178 19124 27806
rect 19292 27860 19348 27916
rect 19628 27860 19684 28700
rect 21308 28532 21364 28542
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19740 27860 19796 27870
rect 19292 27858 19572 27860
rect 19292 27806 19294 27858
rect 19346 27806 19572 27858
rect 19292 27804 19572 27806
rect 19628 27858 19796 27860
rect 19628 27806 19742 27858
rect 19794 27806 19796 27858
rect 19628 27804 19796 27806
rect 19292 27794 19348 27804
rect 19516 27636 19572 27804
rect 19740 27794 19796 27804
rect 20524 27748 20580 27758
rect 20524 27654 20580 27692
rect 19516 27580 19796 27636
rect 19740 27188 19796 27580
rect 19740 27094 19796 27132
rect 21308 27186 21364 28476
rect 21308 27134 21310 27186
rect 21362 27134 21364 27186
rect 21308 27122 21364 27134
rect 22652 27746 22708 27758
rect 22652 27694 22654 27746
rect 22706 27694 22708 27746
rect 21420 27074 21476 27086
rect 21420 27022 21422 27074
rect 21474 27022 21476 27074
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26404 19684 26414
rect 19628 26310 19684 26348
rect 19068 26126 19070 26178
rect 19122 26126 19124 26178
rect 19068 26114 19124 26126
rect 19292 26290 19348 26302
rect 19292 26238 19294 26290
rect 19346 26238 19348 26290
rect 18844 26012 19012 26068
rect 18396 24322 18452 24332
rect 18396 23492 18452 23502
rect 18452 23436 18564 23492
rect 18396 23426 18452 23436
rect 17948 22876 18116 22932
rect 18396 23156 18452 23166
rect 17948 22484 18004 22876
rect 17948 22428 18340 22484
rect 17948 22370 18004 22428
rect 17948 22318 17950 22370
rect 18002 22318 18004 22370
rect 17948 22306 18004 22318
rect 18284 22370 18340 22428
rect 18284 22318 18286 22370
rect 18338 22318 18340 22370
rect 18284 22306 18340 22318
rect 17612 22146 17892 22148
rect 17612 22094 17614 22146
rect 17666 22094 17892 22146
rect 17612 22092 17892 22094
rect 18396 22258 18452 23100
rect 18396 22206 18398 22258
rect 18450 22206 18452 22258
rect 17612 20188 17668 22092
rect 18396 22036 18452 22206
rect 18508 22148 18564 23436
rect 18844 23042 18900 23054
rect 18844 22990 18846 23042
rect 18898 22990 18900 23042
rect 18844 22708 18900 22990
rect 18620 22652 18900 22708
rect 18620 22370 18676 22652
rect 18620 22318 18622 22370
rect 18674 22318 18676 22370
rect 18620 22306 18676 22318
rect 18956 22148 19012 26012
rect 19180 23828 19236 23838
rect 19180 23156 19236 23772
rect 19180 23062 19236 23100
rect 19292 22930 19348 26238
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 21420 24052 21476 27022
rect 21756 27076 21812 27086
rect 21756 26982 21812 27020
rect 22652 27076 22708 27694
rect 22652 27010 22708 27020
rect 22988 26852 23044 35308
rect 23324 34244 23380 34254
rect 23324 34150 23380 34188
rect 23436 34242 23492 36428
rect 24556 37044 24612 37054
rect 23660 36372 23716 36382
rect 23660 35810 23716 36316
rect 24556 35922 24612 36988
rect 25564 37044 25620 38222
rect 25564 36950 25620 36988
rect 25788 38162 25844 38174
rect 25788 38110 25790 38162
rect 25842 38110 25844 38162
rect 25788 37154 25844 38110
rect 25788 37102 25790 37154
rect 25842 37102 25844 37154
rect 25788 36932 25844 37102
rect 25788 36866 25844 36876
rect 26012 37938 26068 37950
rect 26012 37886 26014 37938
rect 26066 37886 26068 37938
rect 26012 37828 26068 37886
rect 26572 37828 26628 37838
rect 26012 37826 26628 37828
rect 26012 37774 26574 37826
rect 26626 37774 26628 37826
rect 26012 37772 26628 37774
rect 24556 35870 24558 35922
rect 24610 35870 24612 35922
rect 24556 35858 24612 35870
rect 23660 35758 23662 35810
rect 23714 35758 23716 35810
rect 23660 35746 23716 35758
rect 23436 34190 23438 34242
rect 23490 34190 23492 34242
rect 23436 34178 23492 34190
rect 23548 35698 23604 35710
rect 23548 35646 23550 35698
rect 23602 35646 23604 35698
rect 23548 34132 23604 35646
rect 24668 35700 24724 35710
rect 24668 35698 25172 35700
rect 24668 35646 24670 35698
rect 24722 35646 25172 35698
rect 24668 35644 25172 35646
rect 24668 35634 24724 35644
rect 24444 34916 24500 34926
rect 24444 34822 24500 34860
rect 24220 34692 24276 34702
rect 23548 34066 23604 34076
rect 24108 34636 24220 34692
rect 23884 34020 23940 34030
rect 23884 33926 23940 33964
rect 23100 33906 23156 33918
rect 23100 33854 23102 33906
rect 23154 33854 23156 33906
rect 23100 32900 23156 33854
rect 23660 33908 23716 33918
rect 23660 33814 23716 33852
rect 23100 32834 23156 32844
rect 22988 26516 23044 26796
rect 23212 26516 23268 26526
rect 22988 26514 23268 26516
rect 22988 26462 23214 26514
rect 23266 26462 23268 26514
rect 22988 26460 23268 26462
rect 23212 26450 23268 26460
rect 23772 26180 23828 26190
rect 23772 25844 23828 26124
rect 23772 25778 23828 25788
rect 20748 24050 21476 24052
rect 20748 23998 21422 24050
rect 21474 23998 21476 24050
rect 20748 23996 21476 23998
rect 20748 23938 20804 23996
rect 21420 23986 21476 23996
rect 20748 23886 20750 23938
rect 20802 23886 20804 23938
rect 20748 23874 20804 23886
rect 20412 23828 20468 23838
rect 20412 23734 20468 23772
rect 21756 23828 21812 23838
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19292 22878 19294 22930
rect 19346 22878 19348 22930
rect 19292 22370 19348 22878
rect 19292 22318 19294 22370
rect 19346 22318 19348 22370
rect 19292 22306 19348 22318
rect 19740 23156 19796 23166
rect 19740 22370 19796 23100
rect 21756 22594 21812 23772
rect 23548 23828 23604 23838
rect 23548 23734 23604 23772
rect 21756 22542 21758 22594
rect 21810 22542 21812 22594
rect 21756 22530 21812 22542
rect 19852 22484 19908 22494
rect 19852 22390 19908 22428
rect 21420 22484 21476 22494
rect 21420 22390 21476 22428
rect 19740 22318 19742 22370
rect 19794 22318 19796 22370
rect 19740 22306 19796 22318
rect 21980 22372 22036 22382
rect 22204 22372 22260 22382
rect 22036 22370 22260 22372
rect 22036 22318 22206 22370
rect 22258 22318 22260 22370
rect 22036 22316 22260 22318
rect 18508 22092 18900 22148
rect 18956 22092 19348 22148
rect 18284 21980 18452 22036
rect 18284 20692 18340 21980
rect 17612 20132 18004 20188
rect 17612 20020 17668 20030
rect 17612 19926 17668 19964
rect 17948 20020 18004 20132
rect 17948 20018 18228 20020
rect 17948 19966 17950 20018
rect 18002 19966 18228 20018
rect 17948 19964 18228 19966
rect 17948 19954 18004 19964
rect 16492 19854 16494 19906
rect 16546 19854 16548 19906
rect 16492 19842 16548 19854
rect 18060 17668 18116 17678
rect 17500 17666 18116 17668
rect 17500 17614 18062 17666
rect 18114 17614 18116 17666
rect 17500 17612 18116 17614
rect 17500 16994 17556 17612
rect 18060 17602 18116 17612
rect 18172 17554 18228 19964
rect 18284 20018 18340 20636
rect 18284 19966 18286 20018
rect 18338 19966 18340 20018
rect 18284 19954 18340 19966
rect 18396 21812 18452 21822
rect 18172 17502 18174 17554
rect 18226 17502 18228 17554
rect 17948 17444 18004 17454
rect 17948 17350 18004 17388
rect 18172 17332 18228 17502
rect 18060 17276 18228 17332
rect 18284 17554 18340 17566
rect 18284 17502 18286 17554
rect 18338 17502 18340 17554
rect 17948 17108 18004 17118
rect 18060 17108 18116 17276
rect 18284 17220 18340 17502
rect 18284 17154 18340 17164
rect 17948 17106 18116 17108
rect 17948 17054 17950 17106
rect 18002 17054 18116 17106
rect 17948 17052 18116 17054
rect 17948 17042 18004 17052
rect 17500 16942 17502 16994
rect 17554 16942 17556 16994
rect 17500 16930 17556 16942
rect 16604 16884 16660 16894
rect 16604 16790 16660 16828
rect 17836 16882 17892 16894
rect 17836 16830 17838 16882
rect 17890 16830 17892 16882
rect 17388 16660 17444 16670
rect 17388 16566 17444 16604
rect 17836 16100 17892 16830
rect 17948 16884 18004 16894
rect 18396 16884 18452 21756
rect 18844 20916 18900 22092
rect 18844 20802 18900 20860
rect 18844 20750 18846 20802
rect 18898 20750 18900 20802
rect 18844 20738 18900 20750
rect 19180 20692 19236 20702
rect 19180 20356 19236 20636
rect 19180 20290 19236 20300
rect 18844 20132 18900 20142
rect 19180 20132 19236 20142
rect 18900 20130 19236 20132
rect 18900 20078 19182 20130
rect 19234 20078 19236 20130
rect 18900 20076 19236 20078
rect 18844 20038 18900 20076
rect 17948 16658 18004 16828
rect 17948 16606 17950 16658
rect 18002 16606 18004 16658
rect 17948 16594 18004 16606
rect 18060 16828 18452 16884
rect 18508 20020 18564 20030
rect 17892 16044 18004 16100
rect 17836 16034 17892 16044
rect 16716 14644 16772 14654
rect 16716 13524 16772 14588
rect 16716 13468 16884 13524
rect 16828 12402 16884 13468
rect 17948 12516 18004 16044
rect 18060 14642 18116 16828
rect 18060 14590 18062 14642
rect 18114 14590 18116 14642
rect 18060 14578 18116 14590
rect 18508 16210 18564 19964
rect 18956 19346 19012 20076
rect 19180 20066 19236 20076
rect 18956 19294 18958 19346
rect 19010 19294 19012 19346
rect 18956 19282 19012 19294
rect 18620 17780 18676 17790
rect 18620 17666 18676 17724
rect 19180 17780 19236 17790
rect 19180 17686 19236 17724
rect 18620 17614 18622 17666
rect 18674 17614 18676 17666
rect 18620 17602 18676 17614
rect 19292 17108 19348 22092
rect 19516 22146 19572 22158
rect 19852 22148 19908 22158
rect 19516 22094 19518 22146
rect 19570 22094 19572 22146
rect 19404 20244 19460 20254
rect 19404 20020 19460 20188
rect 19516 20020 19572 22094
rect 19628 22146 19908 22148
rect 19628 22094 19854 22146
rect 19906 22094 19908 22146
rect 19628 22092 19908 22094
rect 19628 21588 19684 22092
rect 19852 22082 19908 22092
rect 21644 22146 21700 22158
rect 21644 22094 21646 22146
rect 21698 22094 21700 22146
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19684 21532 19796 21588
rect 19628 21522 19684 21532
rect 19628 20916 19684 20926
rect 19628 20822 19684 20860
rect 19740 20580 19796 21532
rect 19852 20916 19908 20926
rect 19852 20580 19908 20860
rect 19852 20524 20244 20580
rect 19740 20514 19796 20524
rect 19836 20412 20100 20422
rect 19628 20356 19684 20366
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19628 20242 19684 20300
rect 19628 20190 19630 20242
rect 19682 20190 19684 20242
rect 19628 20178 19684 20190
rect 19740 20244 19796 20254
rect 19404 20018 19572 20020
rect 19404 19966 19406 20018
rect 19458 19966 19572 20018
rect 19404 19964 19572 19966
rect 19740 20018 19796 20188
rect 19740 19966 19742 20018
rect 19794 19966 19796 20018
rect 19404 19954 19460 19964
rect 19740 19954 19796 19966
rect 19628 19908 19684 19918
rect 19628 19814 19684 19852
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18674 20244 20524
rect 21644 20188 21700 22094
rect 21980 21810 22036 22316
rect 22204 22306 22260 22316
rect 21980 21758 21982 21810
rect 22034 21758 22036 21810
rect 21980 21746 22036 21758
rect 23772 20916 23828 20926
rect 24108 20916 24164 34636
rect 24220 34598 24276 34636
rect 25116 34244 25172 35644
rect 25228 34916 25284 34926
rect 25228 34822 25284 34860
rect 26012 34692 26068 37772
rect 26572 37762 26628 37772
rect 26684 36932 26740 38782
rect 27244 38836 27300 38846
rect 27244 38742 27300 38780
rect 29708 38836 29764 38846
rect 26684 36866 26740 36876
rect 27132 36932 27188 36942
rect 27132 35026 27188 36876
rect 29708 35810 29764 38780
rect 29820 38724 29876 39564
rect 30492 39508 30548 39518
rect 30492 39414 30548 39452
rect 29820 38658 29876 38668
rect 30492 38724 30548 38734
rect 29708 35758 29710 35810
rect 29762 35758 29764 35810
rect 29708 35746 29764 35758
rect 30492 35700 30548 38668
rect 31164 38724 31220 40348
rect 32620 39730 32676 41918
rect 35980 41970 36372 41972
rect 35980 41918 36318 41970
rect 36370 41918 36372 41970
rect 35980 41916 36372 41918
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 33180 40404 33236 40414
rect 32620 39678 32622 39730
rect 32674 39678 32676 39730
rect 32620 39666 32676 39678
rect 33068 40348 33180 40404
rect 33068 39730 33124 40348
rect 33180 40310 33236 40348
rect 33068 39678 33070 39730
rect 33122 39678 33124 39730
rect 33068 39666 33124 39678
rect 33852 40290 33908 40302
rect 33852 40238 33854 40290
rect 33906 40238 33908 40290
rect 33852 39060 33908 40238
rect 35980 40290 36036 41916
rect 36316 41906 36372 41916
rect 36876 41860 36932 45276
rect 39872 45200 39984 46000
rect 43680 45200 43792 46000
rect 37324 41860 37380 41870
rect 36876 41858 37380 41860
rect 36876 41806 37326 41858
rect 37378 41806 37380 41858
rect 36876 41804 37380 41806
rect 37324 41794 37380 41804
rect 39900 41860 39956 45200
rect 39900 41794 39956 41804
rect 40348 41970 40404 41982
rect 40348 41918 40350 41970
rect 40402 41918 40404 41970
rect 36428 40404 36484 40414
rect 36428 40310 36484 40348
rect 35980 40238 35982 40290
rect 36034 40238 36036 40290
rect 35980 40226 36036 40238
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 39228 39730 39284 39742
rect 39228 39678 39230 39730
rect 39282 39678 39284 39730
rect 38892 39396 38948 39406
rect 33852 38994 33908 39004
rect 38332 39060 38388 39070
rect 38332 38966 38388 39004
rect 37324 38948 37380 38958
rect 31164 38658 31220 38668
rect 34636 38722 34692 38734
rect 34636 38670 34638 38722
rect 34690 38670 34692 38722
rect 34636 37940 34692 38670
rect 36764 38722 36820 38734
rect 36764 38670 36766 38722
rect 36818 38670 36820 38722
rect 36764 38612 36820 38670
rect 36764 38546 36820 38556
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34636 37874 34692 37884
rect 37100 37938 37156 37950
rect 37100 37886 37102 37938
rect 37154 37886 37156 37938
rect 37100 37044 37156 37886
rect 37212 37940 37268 37950
rect 37212 37846 37268 37884
rect 37100 36978 37156 36988
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 37100 36484 37156 36494
rect 37100 36372 37156 36428
rect 36988 36370 37156 36372
rect 36988 36318 37102 36370
rect 37154 36318 37156 36370
rect 36988 36316 37156 36318
rect 30940 35700 30996 35710
rect 30492 35698 30996 35700
rect 30492 35646 30494 35698
rect 30546 35646 30942 35698
rect 30994 35646 30996 35698
rect 30492 35644 30996 35646
rect 30492 35634 30548 35644
rect 27132 34974 27134 35026
rect 27186 34974 27188 35026
rect 27132 34962 27188 34974
rect 27580 35586 27636 35598
rect 27580 35534 27582 35586
rect 27634 35534 27636 35586
rect 26684 34916 26740 34926
rect 27020 34916 27076 34926
rect 26012 34626 26068 34636
rect 26460 34914 26740 34916
rect 26460 34862 26686 34914
rect 26738 34862 26740 34914
rect 26460 34860 26740 34862
rect 25228 34244 25284 34254
rect 25116 34242 25284 34244
rect 25116 34190 25230 34242
rect 25282 34190 25284 34242
rect 25116 34188 25284 34190
rect 25228 34178 25284 34188
rect 25340 34132 25396 34142
rect 25340 34038 25396 34076
rect 25788 34130 25844 34142
rect 25788 34078 25790 34130
rect 25842 34078 25844 34130
rect 25788 34020 25844 34078
rect 24892 33908 24948 33918
rect 24892 32564 24948 33852
rect 25564 33908 25620 33918
rect 25564 33814 25620 33852
rect 25788 33572 25844 33964
rect 25788 33516 26180 33572
rect 25900 33346 25956 33358
rect 25900 33294 25902 33346
rect 25954 33294 25956 33346
rect 24892 31890 24948 32508
rect 25564 33234 25620 33246
rect 25564 33182 25566 33234
rect 25618 33182 25620 33234
rect 25564 32004 25620 33182
rect 25788 32674 25844 32686
rect 25788 32622 25790 32674
rect 25842 32622 25844 32674
rect 25676 32452 25732 32462
rect 25676 32358 25732 32396
rect 25676 32004 25732 32014
rect 25564 32002 25732 32004
rect 25564 31950 25678 32002
rect 25730 31950 25732 32002
rect 25564 31948 25732 31950
rect 25676 31938 25732 31948
rect 24892 31838 24894 31890
rect 24946 31838 24948 31890
rect 24892 31826 24948 31838
rect 25788 31892 25844 32622
rect 25228 31780 25284 31790
rect 25228 31686 25284 31724
rect 25452 31780 25508 31790
rect 25788 31780 25844 31836
rect 25452 31778 25844 31780
rect 25452 31726 25454 31778
rect 25506 31726 25844 31778
rect 25452 31724 25844 31726
rect 25452 31714 25508 31724
rect 25564 31444 25620 31454
rect 25564 30994 25620 31388
rect 25564 30942 25566 30994
rect 25618 30942 25620 30994
rect 25564 30772 25620 30942
rect 25788 30996 25844 31724
rect 25900 31218 25956 33294
rect 25900 31166 25902 31218
rect 25954 31166 25956 31218
rect 25900 31154 25956 31166
rect 26012 32338 26068 32350
rect 26012 32286 26014 32338
rect 26066 32286 26068 32338
rect 26012 31220 26068 32286
rect 26124 31948 26180 33516
rect 26460 33122 26516 34860
rect 26684 34850 26740 34860
rect 26796 34914 27076 34916
rect 26796 34862 27022 34914
rect 27074 34862 27076 34914
rect 26796 34860 27076 34862
rect 26796 34132 26852 34860
rect 27020 34850 27076 34860
rect 27580 34804 27636 35534
rect 30604 34914 30660 35644
rect 30940 35634 30996 35644
rect 36764 35700 36820 35710
rect 36764 35606 36820 35644
rect 33852 35586 33908 35598
rect 33852 35534 33854 35586
rect 33906 35534 33908 35586
rect 30604 34862 30606 34914
rect 30658 34862 30660 34914
rect 28028 34804 28084 34814
rect 27580 34802 28084 34804
rect 27580 34750 28030 34802
rect 28082 34750 28084 34802
rect 27580 34748 28084 34750
rect 28028 34738 28084 34748
rect 30604 34692 30660 34862
rect 33404 35140 33460 35150
rect 33404 35026 33460 35084
rect 33404 34974 33406 35026
rect 33458 34974 33460 35026
rect 31276 34804 31332 34814
rect 31276 34710 31332 34748
rect 32060 34804 32116 34814
rect 30604 34626 30660 34636
rect 32060 34354 32116 34748
rect 32060 34302 32062 34354
rect 32114 34302 32116 34354
rect 32060 34290 32116 34302
rect 30828 34244 30884 34254
rect 26796 33572 26852 34076
rect 30156 34132 30212 34142
rect 29708 34020 29764 34030
rect 26572 33516 26852 33572
rect 29596 33964 29708 34020
rect 26572 33346 26628 33516
rect 26572 33294 26574 33346
rect 26626 33294 26628 33346
rect 26572 33282 26628 33294
rect 26460 33070 26462 33122
rect 26514 33070 26516 33122
rect 26460 33058 26516 33070
rect 26124 31892 26292 31948
rect 26124 31778 26180 31790
rect 26124 31726 26126 31778
rect 26178 31726 26180 31778
rect 26124 31444 26180 31726
rect 26236 31556 26292 31892
rect 26348 31892 26404 31902
rect 26348 31798 26404 31836
rect 26460 31780 26516 31790
rect 26460 31556 26516 31724
rect 26572 31780 26628 31790
rect 26572 31778 26852 31780
rect 26572 31726 26574 31778
rect 26626 31726 26852 31778
rect 26572 31724 26852 31726
rect 26572 31714 26628 31724
rect 26236 31500 26404 31556
rect 26460 31500 26740 31556
rect 26124 31378 26180 31388
rect 26012 31164 26180 31220
rect 26012 30996 26068 31006
rect 25788 30940 26012 30996
rect 26012 30902 26068 30940
rect 25564 30210 25620 30716
rect 26124 30212 26180 31164
rect 26236 30996 26292 31006
rect 26348 30996 26404 31500
rect 26684 31218 26740 31500
rect 26684 31166 26686 31218
rect 26738 31166 26740 31218
rect 26684 31154 26740 31166
rect 26236 30994 26404 30996
rect 26236 30942 26238 30994
rect 26290 30942 26404 30994
rect 26236 30940 26404 30942
rect 26236 30930 26292 30940
rect 26236 30212 26292 30222
rect 25564 30158 25566 30210
rect 25618 30158 25620 30210
rect 25564 30146 25620 30158
rect 26012 30210 26292 30212
rect 26012 30158 26238 30210
rect 26290 30158 26292 30210
rect 26012 30156 26292 30158
rect 25900 30100 25956 30110
rect 25900 30006 25956 30044
rect 25788 29988 25844 29998
rect 25788 29894 25844 29932
rect 25564 29538 25620 29550
rect 25564 29486 25566 29538
rect 25618 29486 25620 29538
rect 25228 29426 25284 29438
rect 25228 29374 25230 29426
rect 25282 29374 25284 29426
rect 24668 29316 24724 29326
rect 25228 29316 25284 29374
rect 25564 29428 25620 29486
rect 26012 29538 26068 30156
rect 26236 30146 26292 30156
rect 26348 29986 26404 30940
rect 26796 30996 26852 31724
rect 29036 31108 29092 31118
rect 29036 31014 29092 31052
rect 26908 30996 26964 31006
rect 26796 30940 26908 30996
rect 26572 30882 26628 30894
rect 26572 30830 26574 30882
rect 26626 30830 26628 30882
rect 26460 30772 26516 30782
rect 26572 30772 26628 30830
rect 26516 30716 26628 30772
rect 26684 30884 26740 30894
rect 26460 30706 26516 30716
rect 26348 29934 26350 29986
rect 26402 29934 26404 29986
rect 26348 29922 26404 29934
rect 26460 30548 26516 30558
rect 26012 29486 26014 29538
rect 26066 29486 26068 29538
rect 26012 29474 26068 29486
rect 25564 29362 25620 29372
rect 26460 29426 26516 30492
rect 26460 29374 26462 29426
rect 26514 29374 26516 29426
rect 26460 29362 26516 29374
rect 24724 29260 25284 29316
rect 23772 20914 24164 20916
rect 23772 20862 23774 20914
rect 23826 20862 24110 20914
rect 24162 20862 24164 20914
rect 23772 20860 24164 20862
rect 23772 20850 23828 20860
rect 20972 20132 21700 20188
rect 23996 20244 24052 20860
rect 24108 20850 24164 20860
rect 24220 23938 24276 23950
rect 24220 23886 24222 23938
rect 24274 23886 24276 23938
rect 24220 21588 24276 23886
rect 23996 20178 24052 20188
rect 20972 20018 21028 20132
rect 20972 19966 20974 20018
rect 21026 19966 21028 20018
rect 20972 19954 21028 19966
rect 20636 19908 20692 19918
rect 20636 19814 20692 19852
rect 20188 18622 20190 18674
rect 20242 18622 20244 18674
rect 20188 18610 20244 18622
rect 20972 19794 21028 19806
rect 20972 19742 20974 19794
rect 21026 19742 21028 19794
rect 20972 18452 21028 19742
rect 20972 18386 21028 18396
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19292 17042 19348 17052
rect 19740 17108 19796 17118
rect 19740 16882 19796 17052
rect 20636 17108 20692 17118
rect 20636 17014 20692 17052
rect 19740 16830 19742 16882
rect 19794 16830 19796 16882
rect 19740 16818 19796 16830
rect 20188 16884 20244 16894
rect 20076 16772 20132 16782
rect 20188 16772 20244 16828
rect 20972 16884 21028 16894
rect 20972 16790 21028 16828
rect 20076 16770 20244 16772
rect 20076 16718 20078 16770
rect 20130 16718 20244 16770
rect 20076 16716 20244 16718
rect 21420 16772 21476 16782
rect 20076 16706 20132 16716
rect 18508 16158 18510 16210
rect 18562 16158 18564 16210
rect 18508 14644 18564 16158
rect 19740 16658 19796 16670
rect 19740 16606 19742 16658
rect 19794 16606 19796 16658
rect 19740 15876 19796 16606
rect 21420 16210 21476 16716
rect 21644 16660 21700 20132
rect 22988 20132 23044 20142
rect 22988 18564 23044 20076
rect 23660 20132 23716 20142
rect 23660 20038 23716 20076
rect 22428 18452 22484 18462
rect 22428 18358 22484 18396
rect 22540 16994 22596 17006
rect 22540 16942 22542 16994
rect 22594 16942 22596 16994
rect 22316 16884 22372 16894
rect 22316 16882 22484 16884
rect 22316 16830 22318 16882
rect 22370 16830 22484 16882
rect 22316 16828 22484 16830
rect 22316 16818 22372 16828
rect 21700 16604 21924 16660
rect 21644 16594 21700 16604
rect 21420 16158 21422 16210
rect 21474 16158 21476 16210
rect 21420 16146 21476 16158
rect 19740 15810 19796 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 21868 15538 21924 16604
rect 21868 15486 21870 15538
rect 21922 15486 21924 15538
rect 21868 15474 21924 15486
rect 22428 16436 22484 16828
rect 22540 16660 22596 16942
rect 22540 16594 22596 16604
rect 22988 16882 23044 18508
rect 23212 18450 23268 18462
rect 23212 18398 23214 18450
rect 23266 18398 23268 18450
rect 23212 18340 23268 18398
rect 23660 18340 23716 18350
rect 23212 18338 23716 18340
rect 23212 18286 23662 18338
rect 23714 18286 23716 18338
rect 23212 18284 23716 18286
rect 23660 17444 23716 18284
rect 23660 17378 23716 17388
rect 23772 17666 23828 17678
rect 23772 17614 23774 17666
rect 23826 17614 23828 17666
rect 22988 16830 22990 16882
rect 23042 16830 23044 16882
rect 22988 16436 23044 16830
rect 23772 16660 23828 17614
rect 24220 17668 24276 21532
rect 24444 20804 24500 20814
rect 24444 20690 24500 20748
rect 24444 20638 24446 20690
rect 24498 20638 24500 20690
rect 24444 20626 24500 20638
rect 24556 20244 24612 20282
rect 24556 20178 24612 20188
rect 24556 17668 24612 17678
rect 24220 17666 24612 17668
rect 24220 17614 24558 17666
rect 24610 17614 24612 17666
rect 24220 17612 24612 17614
rect 23996 17556 24052 17566
rect 23996 17462 24052 17500
rect 24108 17554 24164 17566
rect 24108 17502 24110 17554
rect 24162 17502 24164 17554
rect 24108 16996 24164 17502
rect 24556 17444 24612 17612
rect 24556 17378 24612 17388
rect 24108 16930 24164 16940
rect 23772 16594 23828 16604
rect 22428 16380 23044 16436
rect 20636 15204 20692 15214
rect 18508 14550 18564 14588
rect 19516 14644 19572 14654
rect 19516 13972 19572 14588
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19516 13970 19908 13972
rect 19516 13918 19518 13970
rect 19570 13918 19908 13970
rect 19516 13916 19908 13918
rect 19516 13906 19572 13916
rect 19852 13746 19908 13916
rect 20636 13858 20692 15148
rect 21756 15204 21812 15214
rect 21756 15110 21812 15148
rect 20636 13806 20638 13858
rect 20690 13806 20692 13858
rect 20636 13794 20692 13806
rect 22092 15090 22148 15102
rect 22092 15038 22094 15090
rect 22146 15038 22148 15090
rect 19852 13694 19854 13746
rect 19906 13694 19908 13746
rect 19852 13412 19908 13694
rect 22092 13636 22148 15038
rect 22092 13570 22148 13580
rect 19852 13346 19908 13356
rect 20524 13412 20580 13422
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 17948 12460 18116 12516
rect 19836 12506 20100 12516
rect 16828 12350 16830 12402
rect 16882 12350 16884 12402
rect 16828 12338 16884 12350
rect 17724 12066 17780 12078
rect 17724 12014 17726 12066
rect 17778 12014 17780 12066
rect 16828 11396 16884 11406
rect 17052 11396 17108 11406
rect 16828 11394 17108 11396
rect 16828 11342 16830 11394
rect 16882 11342 17054 11394
rect 17106 11342 17108 11394
rect 16828 11340 17108 11342
rect 16828 11330 16884 11340
rect 17052 11330 17108 11340
rect 17388 11396 17444 11406
rect 17388 11302 17444 11340
rect 17612 11396 17668 11434
rect 17612 11330 17668 11340
rect 16716 11284 16772 11294
rect 16604 11228 16716 11284
rect 16268 9886 16270 9938
rect 16322 9886 16324 9938
rect 16268 9874 16324 9886
rect 16380 10610 16436 10622
rect 16380 10558 16382 10610
rect 16434 10558 16436 10610
rect 14588 9662 14590 9714
rect 14642 9662 14644 9714
rect 14588 9604 14644 9662
rect 14588 9538 14644 9548
rect 16380 9266 16436 10558
rect 16604 10612 16660 11228
rect 16716 11190 16772 11228
rect 17724 11284 17780 12014
rect 17948 12068 18004 12078
rect 17836 11732 17892 11742
rect 17836 11506 17892 11676
rect 17836 11454 17838 11506
rect 17890 11454 17892 11506
rect 17836 11442 17892 11454
rect 17948 11506 18004 12012
rect 17948 11454 17950 11506
rect 18002 11454 18004 11506
rect 17948 11442 18004 11454
rect 17724 11218 17780 11228
rect 18060 11394 18116 12460
rect 20524 12178 20580 13356
rect 20524 12126 20526 12178
rect 20578 12126 20580 12178
rect 19852 12068 19908 12078
rect 19852 11974 19908 12012
rect 18060 11342 18062 11394
rect 18114 11342 18116 11394
rect 18060 11284 18116 11342
rect 18284 11732 18340 11742
rect 18284 11394 18340 11676
rect 18284 11342 18286 11394
rect 18338 11342 18340 11394
rect 18284 11330 18340 11342
rect 18060 11218 18116 11228
rect 18620 11284 18676 11294
rect 18620 11190 18676 11228
rect 16604 9826 16660 10556
rect 16604 9774 16606 9826
rect 16658 9774 16660 9826
rect 16604 9762 16660 9774
rect 18844 11170 18900 11182
rect 18844 11118 18846 11170
rect 18898 11118 18900 11170
rect 16380 9214 16382 9266
rect 16434 9214 16436 9266
rect 16380 9202 16436 9214
rect 17388 9716 17444 9726
rect 16492 9156 16548 9166
rect 16492 9062 16548 9100
rect 17388 9156 17444 9660
rect 18172 9716 18228 9726
rect 18172 9622 18228 9660
rect 18844 9716 18900 11118
rect 18956 11172 19012 11182
rect 18956 11170 19236 11172
rect 18956 11118 18958 11170
rect 19010 11118 19236 11170
rect 18956 11116 19236 11118
rect 18956 11106 19012 11116
rect 19068 10052 19124 10062
rect 19068 9826 19124 9996
rect 19068 9774 19070 9826
rect 19122 9774 19124 9826
rect 19068 9762 19124 9774
rect 19180 9826 19236 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19180 9774 19182 9826
rect 19234 9774 19236 9826
rect 19180 9762 19236 9774
rect 19404 9826 19460 9838
rect 19404 9774 19406 9826
rect 19458 9774 19460 9826
rect 18844 9650 18900 9660
rect 14588 9044 14644 9054
rect 14476 9042 14644 9044
rect 14476 8990 14590 9042
rect 14642 8990 14644 9042
rect 14476 8988 14644 8990
rect 13580 8204 13748 8260
rect 13580 8036 13636 8046
rect 13580 7942 13636 7980
rect 12796 6750 12798 6802
rect 12850 6750 12852 6802
rect 12796 6738 12852 6750
rect 13580 6692 13636 6702
rect 13692 6692 13748 8204
rect 13636 6636 13748 6692
rect 13580 6598 13636 6636
rect 13692 6132 13748 6636
rect 13692 6066 13748 6076
rect 12796 6020 12852 6030
rect 12684 6018 12852 6020
rect 12684 5966 12798 6018
rect 12850 5966 12852 6018
rect 12684 5964 12852 5966
rect 12796 5954 12852 5964
rect 12124 5854 12126 5906
rect 12178 5854 12180 5906
rect 12124 5842 12180 5854
rect 14588 5796 14644 8988
rect 17388 7362 17444 9100
rect 18620 9602 18676 9614
rect 18620 9550 18622 9602
rect 18674 9550 18676 9602
rect 18620 8428 18676 9550
rect 19404 9604 19460 9774
rect 19852 9604 19908 9614
rect 19404 9602 19908 9604
rect 19404 9550 19854 9602
rect 19906 9550 19908 9602
rect 19404 9548 19908 9550
rect 19628 9268 19684 9548
rect 19852 9538 19908 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 9202 19684 9212
rect 20524 9268 20580 12126
rect 18284 8372 18676 8428
rect 20524 8428 20580 9212
rect 21420 9268 21476 9278
rect 21420 9174 21476 9212
rect 21868 9268 21924 9278
rect 21868 9042 21924 9212
rect 21868 8990 21870 9042
rect 21922 8990 21924 9042
rect 21868 8978 21924 8990
rect 20524 8372 20804 8428
rect 18284 8258 18340 8372
rect 18284 8206 18286 8258
rect 18338 8206 18340 8258
rect 18284 8194 18340 8206
rect 18508 8036 18564 8046
rect 18508 8034 19572 8036
rect 18508 7982 18510 8034
rect 18562 7982 19572 8034
rect 18508 7980 19572 7982
rect 18508 7970 18564 7980
rect 19516 7586 19572 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19516 7534 19518 7586
rect 19570 7534 19572 7586
rect 19516 7522 19572 7534
rect 17388 7310 17390 7362
rect 17442 7310 17444 7362
rect 17388 7298 17444 7310
rect 20300 7474 20356 7486
rect 20300 7422 20302 7474
rect 20354 7422 20356 7474
rect 20300 7364 20356 7422
rect 20748 7364 20804 8372
rect 22428 8034 22484 16380
rect 24668 16324 24724 29260
rect 25228 27970 25284 27982
rect 25228 27918 25230 27970
rect 25282 27918 25284 27970
rect 25228 27188 25284 27918
rect 25452 27860 25508 27870
rect 26012 27860 26068 27870
rect 25228 27122 25284 27132
rect 25340 27858 26068 27860
rect 25340 27806 25454 27858
rect 25506 27806 26014 27858
rect 26066 27806 26068 27858
rect 25340 27804 26068 27806
rect 25228 26852 25284 26862
rect 24892 26180 24948 26190
rect 24780 23714 24836 23726
rect 24780 23662 24782 23714
rect 24834 23662 24836 23714
rect 24780 21588 24836 23662
rect 24780 21522 24836 21532
rect 24780 20578 24836 20590
rect 24780 20526 24782 20578
rect 24834 20526 24836 20578
rect 24780 20244 24836 20526
rect 24780 20178 24836 20188
rect 24780 16324 24836 16334
rect 24668 16322 24836 16324
rect 24668 16270 24782 16322
rect 24834 16270 24836 16322
rect 24668 16268 24836 16270
rect 24780 16258 24836 16268
rect 24892 13972 24948 26124
rect 25228 24946 25284 26796
rect 25228 24894 25230 24946
rect 25282 24894 25284 24946
rect 25228 24882 25284 24894
rect 25116 20578 25172 20590
rect 25116 20526 25118 20578
rect 25170 20526 25172 20578
rect 25116 20244 25172 20526
rect 25340 20580 25396 27804
rect 25452 27794 25508 27804
rect 26012 27794 26068 27804
rect 25900 27076 25956 27086
rect 25564 26962 25620 26974
rect 25564 26910 25566 26962
rect 25618 26910 25620 26962
rect 25564 26852 25620 26910
rect 25900 26962 25956 27020
rect 25900 26910 25902 26962
rect 25954 26910 25956 26962
rect 25900 26898 25956 26910
rect 25564 26786 25620 26796
rect 25788 24610 25844 24622
rect 25788 24558 25790 24610
rect 25842 24558 25844 24610
rect 25788 23268 25844 24558
rect 25788 22596 25844 23212
rect 25788 22540 25956 22596
rect 25676 22484 25732 22494
rect 25452 21588 25508 21598
rect 25452 21494 25508 21532
rect 25452 20580 25508 20590
rect 25340 20578 25508 20580
rect 25340 20526 25454 20578
rect 25506 20526 25508 20578
rect 25340 20524 25508 20526
rect 25452 20468 25508 20524
rect 25452 20402 25508 20412
rect 25116 20178 25172 20188
rect 25676 17668 25732 22428
rect 25228 17556 25284 17566
rect 25228 17462 25284 17500
rect 25676 16772 25732 17612
rect 25676 16706 25732 16716
rect 25788 20468 25844 20478
rect 25564 16098 25620 16110
rect 25564 16046 25566 16098
rect 25618 16046 25620 16098
rect 25228 15988 25284 15998
rect 25228 15894 25284 15932
rect 25340 15986 25396 15998
rect 25340 15934 25342 15986
rect 25394 15934 25396 15986
rect 25340 15092 25396 15934
rect 25564 15876 25620 16046
rect 25564 15810 25620 15820
rect 25340 14756 25396 15036
rect 25340 14700 25620 14756
rect 24108 13916 24948 13972
rect 22764 13636 22820 13646
rect 22764 13542 22820 13580
rect 22876 13076 22932 13086
rect 22876 12982 22932 13020
rect 23212 9940 23268 9950
rect 23548 9940 23604 9950
rect 23212 9714 23268 9884
rect 23212 9662 23214 9714
rect 23266 9662 23268 9714
rect 23212 9650 23268 9662
rect 23324 9938 23604 9940
rect 23324 9886 23550 9938
rect 23602 9886 23604 9938
rect 23324 9884 23604 9886
rect 23324 9492 23380 9884
rect 23548 9874 23604 9884
rect 24108 9940 24164 13916
rect 24668 13748 24724 13758
rect 24668 13746 24836 13748
rect 24668 13694 24670 13746
rect 24722 13694 24836 13746
rect 24668 13692 24836 13694
rect 24668 13682 24724 13692
rect 24332 13636 24388 13646
rect 24332 13542 24388 13580
rect 24668 13524 24724 13534
rect 24668 13430 24724 13468
rect 24780 13076 24836 13692
rect 25452 13636 25508 13646
rect 25228 13524 25284 13534
rect 24780 12180 24836 13020
rect 25004 13522 25284 13524
rect 25004 13470 25230 13522
rect 25282 13470 25284 13522
rect 25004 13468 25284 13470
rect 25004 13074 25060 13468
rect 25228 13458 25284 13468
rect 25340 13522 25396 13534
rect 25340 13470 25342 13522
rect 25394 13470 25396 13522
rect 25004 13022 25006 13074
rect 25058 13022 25060 13074
rect 25004 13010 25060 13022
rect 25340 13412 25396 13470
rect 25228 12180 25284 12190
rect 24780 12178 25284 12180
rect 24780 12126 25230 12178
rect 25282 12126 25284 12178
rect 24780 12124 25284 12126
rect 25228 12114 25284 12124
rect 25340 11396 25396 13356
rect 25452 12178 25508 13580
rect 25564 13524 25620 14700
rect 25788 14644 25844 20412
rect 25900 17780 25956 22540
rect 26684 22484 26740 30828
rect 26796 30548 26852 30940
rect 26908 30902 26964 30940
rect 29596 30772 29652 33964
rect 29708 33926 29764 33964
rect 30156 34018 30212 34076
rect 30828 34130 30884 34188
rect 31836 34242 31892 34254
rect 31836 34190 31838 34242
rect 31890 34190 31892 34242
rect 30828 34078 30830 34130
rect 30882 34078 30884 34130
rect 30828 34066 30884 34078
rect 30940 34132 30996 34142
rect 30940 34038 30996 34076
rect 31164 34130 31220 34142
rect 31164 34078 31166 34130
rect 31218 34078 31220 34130
rect 30156 33966 30158 34018
rect 30210 33966 30212 34018
rect 30156 33124 30212 33966
rect 31164 34020 31220 34078
rect 31388 34132 31444 34142
rect 31388 34038 31444 34076
rect 31724 34130 31780 34142
rect 31724 34078 31726 34130
rect 31778 34078 31780 34130
rect 31164 33954 31220 33964
rect 31276 34018 31332 34030
rect 31276 33966 31278 34018
rect 31330 33966 31332 34018
rect 31276 33908 31332 33966
rect 31724 33908 31780 34078
rect 31836 34020 31892 34190
rect 33404 34244 33460 34974
rect 33852 34916 33908 35534
rect 35980 35588 36036 35598
rect 35980 35494 36036 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 33852 34850 33908 34860
rect 35084 34916 35140 34926
rect 33852 34692 33908 34702
rect 33852 34598 33908 34636
rect 34636 34692 34692 34702
rect 33404 34178 33460 34188
rect 31836 33954 31892 33964
rect 32284 34132 32340 34142
rect 31276 33852 31780 33908
rect 30156 33058 30212 33068
rect 30492 32450 30548 32462
rect 30492 32398 30494 32450
rect 30546 32398 30548 32450
rect 30380 31780 30436 31790
rect 30380 31686 30436 31724
rect 30492 31780 30548 32398
rect 32284 31948 32340 34076
rect 32396 34020 32452 34030
rect 32396 33926 32452 33964
rect 34524 34020 34580 34030
rect 33740 32788 33796 32798
rect 33740 32694 33796 32732
rect 34188 32788 34244 32798
rect 34188 32562 34244 32732
rect 34188 32510 34190 32562
rect 34242 32510 34244 32562
rect 34188 31948 34244 32510
rect 34524 32452 34580 33964
rect 34636 33460 34692 34636
rect 34636 33458 35028 33460
rect 34636 33406 34638 33458
rect 34690 33406 35028 33458
rect 34636 33404 35028 33406
rect 34636 33394 34692 33404
rect 34972 32564 35028 33404
rect 34860 32562 35028 32564
rect 34860 32510 34974 32562
rect 35026 32510 35028 32562
rect 34860 32508 35028 32510
rect 34636 32452 34692 32462
rect 34524 32450 34692 32452
rect 34524 32398 34638 32450
rect 34690 32398 34692 32450
rect 34524 32396 34692 32398
rect 34636 31948 34692 32396
rect 32284 31892 32452 31948
rect 34188 31892 34468 31948
rect 34636 31892 34804 31948
rect 30716 31780 30772 31790
rect 30492 31778 30772 31780
rect 30492 31726 30718 31778
rect 30770 31726 30772 31778
rect 30492 31724 30772 31726
rect 29820 31556 29876 31566
rect 29596 30706 29652 30716
rect 29708 31554 29876 31556
rect 29708 31502 29822 31554
rect 29874 31502 29876 31554
rect 29708 31500 29876 31502
rect 26796 30482 26852 30492
rect 27356 30210 27412 30222
rect 27356 30158 27358 30210
rect 27410 30158 27412 30210
rect 27244 30098 27300 30110
rect 27244 30046 27246 30098
rect 27298 30046 27300 30098
rect 27244 29988 27300 30046
rect 26908 29932 27244 29988
rect 26908 29426 26964 29932
rect 27244 29922 27300 29932
rect 27356 30100 27412 30158
rect 26908 29374 26910 29426
rect 26962 29374 26964 29426
rect 26908 29362 26964 29374
rect 27356 29092 27412 30044
rect 29708 29988 29764 31500
rect 29820 31490 29876 31500
rect 29932 31554 29988 31566
rect 29932 31502 29934 31554
rect 29986 31502 29988 31554
rect 29820 30996 29876 31006
rect 29932 30996 29988 31502
rect 30044 31556 30100 31566
rect 30044 31554 30324 31556
rect 30044 31502 30046 31554
rect 30098 31502 30324 31554
rect 30044 31500 30324 31502
rect 30044 31490 30100 31500
rect 29820 30994 29988 30996
rect 29820 30942 29822 30994
rect 29874 30942 29988 30994
rect 29820 30940 29988 30942
rect 30268 30996 30324 31500
rect 29820 30930 29876 30940
rect 30268 30212 30324 30940
rect 30492 30884 30548 31724
rect 30716 31714 30772 31724
rect 31388 31780 31444 31790
rect 31444 31724 31780 31780
rect 31388 31714 31444 31724
rect 30492 30818 30548 30828
rect 30828 30994 30884 31006
rect 30828 30942 30830 30994
rect 30882 30942 30884 30994
rect 30380 30212 30436 30222
rect 30268 30210 30436 30212
rect 30268 30158 30382 30210
rect 30434 30158 30436 30210
rect 30268 30156 30436 30158
rect 30380 30146 30436 30156
rect 30604 30212 30660 30222
rect 30604 30118 30660 30156
rect 29708 29540 29764 29932
rect 29820 29540 29876 29550
rect 29708 29484 29820 29540
rect 29820 29474 29876 29484
rect 27356 29026 27412 29036
rect 30380 29092 30436 29102
rect 30380 27298 30436 29036
rect 30380 27246 30382 27298
rect 30434 27246 30436 27298
rect 30380 27234 30436 27246
rect 30716 27300 30772 27310
rect 30716 27206 30772 27244
rect 27020 26964 27076 26974
rect 27020 26290 27076 26908
rect 30044 26964 30100 26974
rect 30828 26908 30884 30942
rect 31276 30884 31332 30894
rect 31276 30790 31332 30828
rect 31276 30212 31332 30222
rect 31164 30156 31276 30212
rect 31052 29428 31108 29438
rect 31052 29334 31108 29372
rect 30044 26870 30100 26908
rect 30380 26852 30884 26908
rect 30940 26962 30996 26974
rect 30940 26910 30942 26962
rect 30994 26910 30996 26962
rect 30044 26404 30100 26414
rect 27020 26238 27022 26290
rect 27074 26238 27076 26290
rect 27020 26226 27076 26238
rect 29820 26292 29876 26302
rect 27692 26178 27748 26190
rect 27692 26126 27694 26178
rect 27746 26126 27748 26178
rect 27692 24948 27748 26126
rect 29484 26180 29540 26190
rect 27692 24882 27748 24892
rect 29260 24948 29316 24958
rect 29260 24854 29316 24892
rect 28700 24836 28756 24846
rect 28700 24742 28756 24780
rect 28588 24724 28644 24734
rect 28476 24668 28588 24724
rect 28252 23156 28308 23166
rect 27580 23044 27636 23054
rect 26684 22390 26740 22428
rect 27356 23042 27636 23044
rect 27356 22990 27582 23042
rect 27634 22990 27636 23042
rect 27356 22988 27636 22990
rect 26124 21476 26180 21486
rect 26124 21382 26180 21420
rect 27020 21476 27076 21486
rect 27020 21026 27076 21420
rect 27020 20974 27022 21026
rect 27074 20974 27076 21026
rect 27020 20962 27076 20974
rect 27356 21026 27412 22988
rect 27580 22978 27636 22988
rect 28252 21474 28308 23100
rect 28476 23154 28532 24668
rect 28588 24630 28644 24668
rect 28924 24724 28980 24734
rect 29148 24724 29204 24734
rect 28924 24722 29204 24724
rect 28924 24670 28926 24722
rect 28978 24670 29150 24722
rect 29202 24670 29204 24722
rect 28924 24668 29204 24670
rect 28924 24658 28980 24668
rect 29148 24658 29204 24668
rect 29484 24722 29540 26124
rect 29820 26180 29876 26236
rect 30044 26290 30100 26348
rect 30044 26238 30046 26290
rect 30098 26238 30100 26290
rect 30044 26226 30100 26238
rect 30268 26180 30324 26190
rect 29820 26178 29988 26180
rect 29820 26126 29822 26178
rect 29874 26126 29988 26178
rect 29820 26124 29988 26126
rect 29820 26114 29876 26124
rect 29484 24670 29486 24722
rect 29538 24670 29540 24722
rect 29484 24658 29540 24670
rect 29596 25394 29652 25406
rect 29596 25342 29598 25394
rect 29650 25342 29652 25394
rect 29596 24724 29652 25342
rect 29932 25394 29988 26124
rect 30268 26086 30324 26124
rect 29932 25342 29934 25394
rect 29986 25342 29988 25394
rect 29932 25330 29988 25342
rect 29932 24836 29988 24846
rect 29932 24742 29988 24780
rect 29596 24658 29652 24668
rect 28476 23102 28478 23154
rect 28530 23102 28532 23154
rect 28476 23090 28532 23102
rect 30380 23156 30436 26852
rect 30940 26516 30996 26910
rect 31164 26908 31220 30156
rect 31276 30118 31332 30156
rect 31724 30210 31780 31724
rect 31724 30158 31726 30210
rect 31778 30158 31780 30210
rect 31724 30146 31780 30158
rect 31948 30212 32004 30222
rect 31948 30098 32004 30156
rect 32396 30212 32452 31892
rect 34076 31668 34132 31678
rect 31948 30046 31950 30098
rect 32002 30046 32004 30098
rect 31948 30034 32004 30046
rect 32060 30100 32116 30110
rect 32060 30006 32116 30044
rect 32396 29650 32452 30156
rect 32396 29598 32398 29650
rect 32450 29598 32452 29650
rect 32396 29586 32452 29598
rect 33964 30772 34020 30782
rect 31276 29540 31332 29550
rect 31276 27186 31332 29484
rect 31724 29540 31780 29550
rect 33628 29540 33684 29550
rect 31724 29538 31892 29540
rect 31724 29486 31726 29538
rect 31778 29486 31892 29538
rect 31724 29484 31892 29486
rect 31724 29474 31780 29484
rect 31500 29428 31556 29438
rect 31500 29334 31556 29372
rect 31836 29428 31892 29484
rect 33628 29446 33684 29484
rect 32060 29428 32116 29438
rect 33292 29428 33348 29438
rect 33964 29428 34020 30716
rect 31836 29426 32116 29428
rect 31836 29374 32062 29426
rect 32114 29374 32116 29426
rect 31836 29372 32116 29374
rect 31836 28868 31892 29372
rect 32060 29362 32116 29372
rect 33068 29372 33292 29428
rect 31276 27134 31278 27186
rect 31330 27134 31332 27186
rect 31276 27122 31332 27134
rect 31500 28812 31892 28868
rect 31500 26908 31556 28812
rect 33068 28754 33124 29372
rect 33292 29334 33348 29372
rect 33740 29426 34020 29428
rect 33740 29374 33966 29426
rect 34018 29374 34020 29426
rect 33740 29372 34020 29374
rect 33068 28702 33070 28754
rect 33122 28702 33124 28754
rect 33068 28690 33124 28702
rect 33628 28756 33684 28766
rect 33740 28756 33796 29372
rect 33964 29362 34020 29372
rect 33628 28754 33796 28756
rect 33628 28702 33630 28754
rect 33682 28702 33796 28754
rect 33628 28700 33796 28702
rect 33628 28690 33684 28700
rect 31836 27748 31892 27758
rect 31836 27300 31892 27692
rect 31836 27074 31892 27244
rect 31836 27022 31838 27074
rect 31890 27022 31892 27074
rect 31836 27010 31892 27022
rect 30604 26460 30996 26516
rect 31052 26852 31220 26908
rect 31276 26852 31556 26908
rect 31724 26962 31780 26974
rect 31724 26910 31726 26962
rect 31778 26910 31780 26962
rect 30492 26292 30548 26302
rect 30604 26292 30660 26460
rect 31052 26404 31108 26852
rect 30492 26290 30660 26292
rect 30492 26238 30494 26290
rect 30546 26238 30660 26290
rect 30492 26236 30660 26238
rect 30716 26348 31108 26404
rect 30716 26292 30772 26348
rect 30492 25396 30548 26236
rect 30716 26198 30772 26236
rect 31276 26292 31332 26852
rect 30828 25508 30884 25518
rect 31276 25508 31332 26236
rect 30828 25506 31332 25508
rect 30828 25454 30830 25506
rect 30882 25454 31332 25506
rect 30828 25452 31332 25454
rect 31612 26404 31668 26414
rect 30828 25442 30884 25452
rect 30716 25396 30772 25406
rect 30492 25394 30772 25396
rect 30492 25342 30718 25394
rect 30770 25342 30772 25394
rect 30492 25340 30772 25342
rect 30716 24836 30772 25340
rect 31276 25284 31332 25294
rect 31612 25284 31668 26348
rect 31276 25282 31612 25284
rect 31276 25230 31278 25282
rect 31330 25230 31612 25282
rect 31276 25228 31612 25230
rect 31276 25218 31332 25228
rect 31612 25190 31668 25228
rect 31388 24836 31444 24846
rect 30716 24834 31444 24836
rect 30716 24782 31390 24834
rect 31442 24782 31444 24834
rect 30716 24780 31444 24782
rect 30380 23090 30436 23100
rect 31388 23154 31444 24780
rect 31612 24724 31668 24734
rect 31724 24724 31780 26910
rect 34076 26964 34132 31612
rect 34412 27076 34468 31892
rect 34748 31220 34804 31892
rect 34860 31668 34916 32508
rect 34972 32498 35028 32508
rect 34860 31602 34916 31612
rect 34748 31126 34804 31164
rect 35084 31106 35140 34860
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35756 33124 35812 33134
rect 35980 33124 36036 33134
rect 35756 33122 36036 33124
rect 35756 33070 35758 33122
rect 35810 33070 35982 33122
rect 36034 33070 36036 33122
rect 35756 33068 36036 33070
rect 35756 32788 35812 33068
rect 35980 33058 36036 33068
rect 36316 33122 36372 33134
rect 36316 33070 36318 33122
rect 36370 33070 36372 33122
rect 35756 32722 35812 32732
rect 36316 32788 36372 33070
rect 36316 32722 36372 32732
rect 35756 32450 35812 32462
rect 35756 32398 35758 32450
rect 35810 32398 35812 32450
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35756 31948 35812 32398
rect 35756 31892 35924 31948
rect 35532 31220 35588 31230
rect 35532 31126 35588 31164
rect 35084 31054 35086 31106
rect 35138 31054 35140 31106
rect 34860 30996 34916 31006
rect 34860 30902 34916 30940
rect 35084 30884 35140 31054
rect 35084 30818 35140 30828
rect 35196 30994 35252 31006
rect 35196 30942 35198 30994
rect 35250 30942 35252 30994
rect 35196 30772 35252 30942
rect 35756 30996 35812 31006
rect 35756 30902 35812 30940
rect 35868 30882 35924 31892
rect 36876 31556 36932 31566
rect 36092 31554 36932 31556
rect 36092 31502 36878 31554
rect 36930 31502 36932 31554
rect 36092 31500 36932 31502
rect 36092 30994 36148 31500
rect 36876 31490 36932 31500
rect 36092 30942 36094 30994
rect 36146 30942 36148 30994
rect 36092 30930 36148 30942
rect 35868 30830 35870 30882
rect 35922 30830 35924 30882
rect 35868 30818 35924 30830
rect 35196 30716 35588 30772
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34860 27748 34916 27758
rect 34860 27654 34916 27692
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34412 26908 34468 27020
rect 34076 26898 34132 26908
rect 34188 26852 34468 26908
rect 31948 26292 32004 26302
rect 31948 26198 32004 26236
rect 32396 26178 32452 26190
rect 32396 26126 32398 26178
rect 32450 26126 32452 26178
rect 32396 25956 32452 26126
rect 32396 25890 32452 25900
rect 31612 24722 31780 24724
rect 31612 24670 31614 24722
rect 31666 24670 31780 24722
rect 31612 24668 31780 24670
rect 33852 24836 33908 24846
rect 31612 23380 31668 24668
rect 31724 23380 31780 23390
rect 31612 23324 31724 23380
rect 31724 23314 31780 23324
rect 32396 23380 32452 23390
rect 31388 23102 31390 23154
rect 31442 23102 31444 23154
rect 31388 23090 31444 23102
rect 30828 23044 30884 23054
rect 30492 23042 30884 23044
rect 30492 22990 30830 23042
rect 30882 22990 30884 23042
rect 30492 22988 30884 22990
rect 29596 21586 29652 21598
rect 29596 21534 29598 21586
rect 29650 21534 29652 21586
rect 28252 21422 28254 21474
rect 28306 21422 28308 21474
rect 28252 21410 28308 21422
rect 28700 21476 28756 21486
rect 28700 21382 28756 21420
rect 29596 21476 29652 21534
rect 29596 21410 29652 21420
rect 30268 21474 30324 21486
rect 30268 21422 30270 21474
rect 30322 21422 30324 21474
rect 27356 20974 27358 21026
rect 27410 20974 27412 21026
rect 27356 20962 27412 20974
rect 30268 20914 30324 21422
rect 30492 21026 30548 22988
rect 30828 22978 30884 22988
rect 31724 23042 31780 23054
rect 31724 22990 31726 23042
rect 31778 22990 31780 23042
rect 31724 22932 31780 22990
rect 31724 22866 31780 22876
rect 32284 23042 32340 23054
rect 32284 22990 32286 23042
rect 32338 22990 32340 23042
rect 32284 22932 32340 22990
rect 30492 20974 30494 21026
rect 30546 20974 30548 21026
rect 30492 20962 30548 20974
rect 30268 20862 30270 20914
rect 30322 20862 30324 20914
rect 30268 20850 30324 20862
rect 26684 20804 26740 20814
rect 27020 20804 27076 20814
rect 26740 20802 27076 20804
rect 26740 20750 27022 20802
rect 27074 20750 27076 20802
rect 26740 20748 27076 20750
rect 26684 20710 26740 20748
rect 27020 20738 27076 20748
rect 29820 20804 29876 20814
rect 30156 20804 30212 20814
rect 29876 20802 30212 20804
rect 29876 20750 30158 20802
rect 30210 20750 30212 20802
rect 29876 20748 30212 20750
rect 29820 20710 29876 20748
rect 30156 20738 30212 20748
rect 32172 20692 32228 20702
rect 32284 20692 32340 22876
rect 32396 21474 32452 23324
rect 33628 22372 33684 22382
rect 33628 22278 33684 22316
rect 32396 21422 32398 21474
rect 32450 21422 32452 21474
rect 32396 21410 32452 21422
rect 33180 21476 33236 21486
rect 32172 20690 32340 20692
rect 32172 20638 32174 20690
rect 32226 20638 32340 20690
rect 32172 20636 32340 20638
rect 32396 20802 32452 20814
rect 32396 20750 32398 20802
rect 32450 20750 32452 20802
rect 32172 20626 32228 20636
rect 31948 20578 32004 20590
rect 31948 20526 31950 20578
rect 32002 20526 32004 20578
rect 31948 20468 32004 20526
rect 32396 20468 32452 20750
rect 31948 20412 32452 20468
rect 31948 19124 32004 20412
rect 29820 18452 29876 18462
rect 28700 18450 29876 18452
rect 28700 18398 29822 18450
rect 29874 18398 29876 18450
rect 28700 18396 29876 18398
rect 25900 17714 25956 17724
rect 27356 17778 27412 17790
rect 27356 17726 27358 17778
rect 27410 17726 27412 17778
rect 26572 16884 26628 16894
rect 26124 15986 26180 15998
rect 26124 15934 26126 15986
rect 26178 15934 26180 15986
rect 26012 15092 26068 15102
rect 26124 15092 26180 15934
rect 26572 15874 26628 16828
rect 27356 16772 27412 17726
rect 27804 17444 27860 17454
rect 28588 17444 28644 17454
rect 27860 17388 28084 17444
rect 27804 17350 27860 17388
rect 27692 16996 27748 17006
rect 27692 16902 27748 16940
rect 27356 16706 27412 16716
rect 26908 16100 26964 16110
rect 26572 15822 26574 15874
rect 26626 15822 26628 15874
rect 26572 15810 26628 15822
rect 26796 15986 26852 15998
rect 26796 15934 26798 15986
rect 26850 15934 26852 15986
rect 26796 15876 26852 15934
rect 26796 15810 26852 15820
rect 26908 15148 26964 16044
rect 26908 15092 27076 15148
rect 26068 15036 26180 15092
rect 26012 15026 26068 15036
rect 25788 14642 26404 14644
rect 25788 14590 25790 14642
rect 25842 14590 26404 14642
rect 25788 14588 26404 14590
rect 25788 14578 25844 14588
rect 26124 13858 26180 13870
rect 26124 13806 26126 13858
rect 26178 13806 26180 13858
rect 25564 13430 25620 13468
rect 25676 13522 25732 13534
rect 25676 13470 25678 13522
rect 25730 13470 25732 13522
rect 25452 12126 25454 12178
rect 25506 12126 25508 12178
rect 25452 12114 25508 12126
rect 25676 11956 25732 13470
rect 26124 13412 26180 13806
rect 26348 13746 26404 14588
rect 26348 13694 26350 13746
rect 26402 13694 26404 13746
rect 26348 13682 26404 13694
rect 27020 13524 27076 15092
rect 27020 13468 27300 13524
rect 26124 13346 26180 13356
rect 25788 12962 25844 12974
rect 25788 12910 25790 12962
rect 25842 12910 25844 12962
rect 25788 12740 25844 12910
rect 26236 12740 26292 12750
rect 25788 12738 26292 12740
rect 25788 12686 26238 12738
rect 26290 12686 26292 12738
rect 25788 12684 26292 12686
rect 26236 12180 26292 12684
rect 26236 12114 26292 12124
rect 26908 12180 26964 12190
rect 25788 11956 25844 11966
rect 25676 11954 25844 11956
rect 25676 11902 25790 11954
rect 25842 11902 25844 11954
rect 25676 11900 25844 11902
rect 25340 11330 25396 11340
rect 25788 11284 25844 11900
rect 25788 11218 25844 11228
rect 24108 9846 24164 9884
rect 23212 9436 23380 9492
rect 23436 9602 23492 9614
rect 23436 9550 23438 9602
rect 23490 9550 23492 9602
rect 22540 8932 22596 8942
rect 22540 8930 23156 8932
rect 22540 8878 22542 8930
rect 22594 8878 23156 8930
rect 22540 8876 23156 8878
rect 22540 8866 22596 8876
rect 22988 8708 23044 8718
rect 22652 8260 22708 8270
rect 22988 8260 23044 8652
rect 23100 8370 23156 8876
rect 23100 8318 23102 8370
rect 23154 8318 23156 8370
rect 23100 8306 23156 8318
rect 22652 8258 23044 8260
rect 22652 8206 22654 8258
rect 22706 8206 22990 8258
rect 23042 8206 23044 8258
rect 22652 8204 23044 8206
rect 22652 8194 22708 8204
rect 22988 8194 23044 8204
rect 23212 8260 23268 9436
rect 23436 9156 23492 9550
rect 23436 8428 23492 9100
rect 23660 9602 23716 9614
rect 23660 9550 23662 9602
rect 23714 9550 23716 9602
rect 23660 8708 23716 9550
rect 26348 9380 26404 9390
rect 25340 9156 25396 9166
rect 25340 9062 25396 9100
rect 24668 9044 24724 9054
rect 24668 8930 24724 8988
rect 25676 9044 25732 9054
rect 25676 8950 25732 8988
rect 24668 8878 24670 8930
rect 24722 8878 24724 8930
rect 24668 8866 24724 8878
rect 23660 8642 23716 8652
rect 23212 8194 23268 8204
rect 23324 8372 23492 8428
rect 26348 8484 26404 9324
rect 23324 8258 23380 8372
rect 23324 8206 23326 8258
rect 23378 8206 23380 8258
rect 23324 8194 23380 8206
rect 23548 8260 23604 8270
rect 23548 8166 23604 8204
rect 22428 7982 22430 8034
rect 22482 7982 22484 8034
rect 22428 7700 22484 7982
rect 22540 8036 22596 8046
rect 22540 8034 23156 8036
rect 22540 7982 22542 8034
rect 22594 7982 23156 8034
rect 22540 7980 23156 7982
rect 22540 7970 22596 7980
rect 22988 7700 23044 7710
rect 22428 7698 23044 7700
rect 22428 7646 22990 7698
rect 23042 7646 23044 7698
rect 22428 7644 23044 7646
rect 22988 7634 23044 7644
rect 20300 7362 20916 7364
rect 20300 7310 20750 7362
rect 20802 7310 20916 7362
rect 20300 7308 20916 7310
rect 20748 7298 20804 7308
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 15372 6132 15428 6142
rect 15372 6038 15428 6076
rect 14924 5796 14980 5806
rect 14588 5794 14980 5796
rect 14588 5742 14926 5794
rect 14978 5742 14980 5794
rect 14588 5740 14980 5742
rect 14924 5730 14980 5740
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 20860 5124 20916 7308
rect 23100 5906 23156 7980
rect 26348 6804 26404 8428
rect 26684 7588 26740 7598
rect 25900 6748 26404 6804
rect 25900 6690 25956 6748
rect 25900 6638 25902 6690
rect 25954 6638 25956 6690
rect 25900 6626 25956 6638
rect 25788 6580 25844 6590
rect 23100 5854 23102 5906
rect 23154 5854 23156 5906
rect 23100 5842 23156 5854
rect 24556 6020 24612 6030
rect 23324 5796 23380 5806
rect 23324 5702 23380 5740
rect 22764 5682 22820 5694
rect 22764 5630 22766 5682
rect 22818 5630 22820 5682
rect 21644 5124 21700 5134
rect 20860 5122 21700 5124
rect 20860 5070 20862 5122
rect 20914 5070 21646 5122
rect 21698 5070 21700 5122
rect 20860 5068 21700 5070
rect 20860 5058 20916 5068
rect 21644 5058 21700 5068
rect 22428 5010 22484 5022
rect 22428 4958 22430 5010
rect 22482 4958 22484 5010
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 22428 4562 22484 4958
rect 22428 4510 22430 4562
rect 22482 4510 22484 4562
rect 22428 4498 22484 4510
rect 22764 4450 22820 5630
rect 24556 5234 24612 5964
rect 25676 5906 25732 5918
rect 25676 5854 25678 5906
rect 25730 5854 25732 5906
rect 25676 5796 25732 5854
rect 25788 5908 25844 6524
rect 26236 6580 26292 6590
rect 26236 6486 26292 6524
rect 26348 6578 26404 6748
rect 26348 6526 26350 6578
rect 26402 6526 26404 6578
rect 26348 6514 26404 6526
rect 26460 7586 26740 7588
rect 26460 7534 26686 7586
rect 26738 7534 26740 7586
rect 26460 7532 26740 7534
rect 25900 6132 25956 6142
rect 25900 6130 26180 6132
rect 25900 6078 25902 6130
rect 25954 6078 26180 6130
rect 25900 6076 26180 6078
rect 25900 6066 25956 6076
rect 26012 5908 26068 5918
rect 25788 5906 26068 5908
rect 25788 5854 26014 5906
rect 26066 5854 26068 5906
rect 25788 5852 26068 5854
rect 26012 5842 26068 5852
rect 25676 5730 25732 5740
rect 26124 5684 26180 6076
rect 26460 6020 26516 7532
rect 26684 7522 26740 7532
rect 26796 6916 26852 6954
rect 26796 6850 26852 6860
rect 26796 6692 26852 6702
rect 26684 6690 26852 6692
rect 26684 6638 26798 6690
rect 26850 6638 26852 6690
rect 26684 6636 26852 6638
rect 26908 6692 26964 12124
rect 27020 11284 27076 11294
rect 27020 8484 27076 11228
rect 27132 9042 27188 9054
rect 27132 8990 27134 9042
rect 27186 8990 27188 9042
rect 27132 8708 27188 8990
rect 27244 8932 27300 13468
rect 28028 12180 28084 17388
rect 28588 17350 28644 17388
rect 28364 16882 28420 16894
rect 28364 16830 28366 16882
rect 28418 16830 28420 16882
rect 28364 16772 28420 16830
rect 28364 16100 28420 16716
rect 28588 16772 28644 16782
rect 28700 16772 28756 18396
rect 29820 18386 29876 18396
rect 30044 18340 30100 18350
rect 30044 18246 30100 18284
rect 31276 18340 31332 18350
rect 30156 18226 30212 18238
rect 30156 18174 30158 18226
rect 30210 18174 30212 18226
rect 30156 17892 30212 18174
rect 30044 17836 30212 17892
rect 29484 17780 29540 17790
rect 28588 16770 28756 16772
rect 28588 16718 28590 16770
rect 28642 16718 28756 16770
rect 28588 16716 28756 16718
rect 28588 16706 28644 16716
rect 28364 16034 28420 16044
rect 28700 15148 28756 16716
rect 29148 16772 29204 16782
rect 29148 16770 29316 16772
rect 29148 16718 29150 16770
rect 29202 16718 29316 16770
rect 29148 16716 29316 16718
rect 29148 16706 29204 16716
rect 29148 16100 29204 16110
rect 29148 16006 29204 16044
rect 29260 15986 29316 16716
rect 29260 15934 29262 15986
rect 29314 15934 29316 15986
rect 29260 15316 29316 15934
rect 29372 15876 29428 15886
rect 29372 15782 29428 15820
rect 29260 15250 29316 15260
rect 29484 15540 29540 17724
rect 30044 16660 30100 17836
rect 30156 17666 30212 17678
rect 30156 17614 30158 17666
rect 30210 17614 30212 17666
rect 30156 17444 30212 17614
rect 30156 16884 30212 17388
rect 31276 16994 31332 18284
rect 31948 17108 32004 19068
rect 33180 17778 33236 21420
rect 33180 17726 33182 17778
rect 33234 17726 33236 17778
rect 33180 17714 33236 17726
rect 33852 17668 33908 24780
rect 33852 17602 33908 17612
rect 31948 17042 32004 17052
rect 31276 16942 31278 16994
rect 31330 16942 31332 16994
rect 31276 16930 31332 16942
rect 32060 16996 32116 17006
rect 30156 16818 30212 16828
rect 32060 16882 32116 16940
rect 32508 16996 32564 17006
rect 32508 16902 32564 16940
rect 33628 16996 33684 17006
rect 32060 16830 32062 16882
rect 32114 16830 32116 16882
rect 32060 16818 32116 16830
rect 33292 16884 33348 16894
rect 30044 16604 30324 16660
rect 28700 15092 29204 15148
rect 29260 15092 29316 15102
rect 29148 15090 29316 15092
rect 29148 15038 29262 15090
rect 29314 15038 29316 15090
rect 29148 15036 29316 15038
rect 29260 15026 29316 15036
rect 29484 14754 29540 15484
rect 30268 15538 30324 16604
rect 32956 16098 33012 16110
rect 32956 16046 32958 16098
rect 33010 16046 33012 16098
rect 32284 15986 32340 15998
rect 32284 15934 32286 15986
rect 32338 15934 32340 15986
rect 30268 15486 30270 15538
rect 30322 15486 30324 15538
rect 30268 15474 30324 15486
rect 30604 15540 30660 15550
rect 30604 15446 30660 15484
rect 30156 15428 30212 15438
rect 29484 14702 29486 14754
rect 29538 14702 29540 14754
rect 29484 14690 29540 14702
rect 29596 15426 30212 15428
rect 29596 15374 30158 15426
rect 30210 15374 30212 15426
rect 29596 15372 30212 15374
rect 29596 15202 29652 15372
rect 30156 15362 30212 15372
rect 30380 15316 30436 15326
rect 29596 15150 29598 15202
rect 29650 15150 29652 15202
rect 29596 13636 29652 15150
rect 29820 15204 29876 15242
rect 30380 15222 30436 15260
rect 29820 15138 29876 15148
rect 29932 14754 29988 14766
rect 29932 14702 29934 14754
rect 29986 14702 29988 14754
rect 29932 14642 29988 14702
rect 29932 14590 29934 14642
rect 29986 14590 29988 14642
rect 29932 14578 29988 14590
rect 29596 13580 29876 13636
rect 29484 13412 29540 13422
rect 29484 13188 29540 13356
rect 29484 13186 29652 13188
rect 29484 13134 29486 13186
rect 29538 13134 29652 13186
rect 29484 13132 29652 13134
rect 29484 13122 29540 13132
rect 29372 12852 29428 12862
rect 28812 12850 29428 12852
rect 28812 12798 29374 12850
rect 29426 12798 29428 12850
rect 28812 12796 29428 12798
rect 28812 12290 28868 12796
rect 29372 12786 29428 12796
rect 28812 12238 28814 12290
rect 28866 12238 28868 12290
rect 28812 12226 28868 12238
rect 29596 12292 29652 13132
rect 29708 12964 29764 12974
rect 29820 12964 29876 13580
rect 30828 13524 30884 13534
rect 29932 12964 29988 12974
rect 29820 12962 29988 12964
rect 29820 12910 29934 12962
rect 29986 12910 29988 12962
rect 29820 12908 29988 12910
rect 29708 12870 29764 12908
rect 29596 12236 29876 12292
rect 28140 12180 28196 12190
rect 28028 12124 28140 12180
rect 28140 12086 28196 12124
rect 29596 10724 29652 10734
rect 28924 10612 28980 10622
rect 27468 9828 27524 9838
rect 27468 9266 27524 9772
rect 27468 9214 27470 9266
rect 27522 9214 27524 9266
rect 27468 9202 27524 9214
rect 28924 9266 28980 10556
rect 29596 10050 29652 10668
rect 29596 9998 29598 10050
rect 29650 9998 29652 10050
rect 29596 9986 29652 9998
rect 29820 10050 29876 12236
rect 29932 11618 29988 12908
rect 30380 12964 30436 12974
rect 30380 12870 30436 12908
rect 30828 12964 30884 13468
rect 32284 13524 32340 15934
rect 32284 13458 32340 13468
rect 32956 12964 33012 16046
rect 33292 15538 33348 16828
rect 33628 16098 33684 16940
rect 33628 16046 33630 16098
rect 33682 16046 33684 16098
rect 33628 16034 33684 16046
rect 33292 15486 33294 15538
rect 33346 15486 33348 15538
rect 33292 15474 33348 15486
rect 34188 14084 34244 26852
rect 35532 26516 35588 30716
rect 36988 30212 37044 36316
rect 37100 36306 37156 36316
rect 37212 36260 37268 36270
rect 37324 36260 37380 38892
rect 37548 38834 37604 38846
rect 37772 38836 37828 38846
rect 37548 38782 37550 38834
rect 37602 38782 37604 38834
rect 37548 38724 37604 38782
rect 37548 38658 37604 38668
rect 37660 38834 37828 38836
rect 37660 38782 37774 38834
rect 37826 38782 37828 38834
rect 37660 38780 37828 38782
rect 37660 38388 37716 38780
rect 37772 38770 37828 38780
rect 38108 38836 38164 38846
rect 38108 38834 38276 38836
rect 38108 38782 38110 38834
rect 38162 38782 38276 38834
rect 38108 38780 38276 38782
rect 38108 38770 38164 38780
rect 37996 38612 38052 38622
rect 37996 38518 38052 38556
rect 37436 38332 37716 38388
rect 37436 38050 37492 38332
rect 37436 37998 37438 38050
rect 37490 37998 37492 38050
rect 37436 37986 37492 37998
rect 37772 37940 37828 37950
rect 37660 36484 37716 36494
rect 37660 36390 37716 36428
rect 37772 36370 37828 37884
rect 37772 36318 37774 36370
rect 37826 36318 37828 36370
rect 37772 36306 37828 36318
rect 37212 36258 37380 36260
rect 37212 36206 37214 36258
rect 37266 36206 37380 36258
rect 37212 36204 37380 36206
rect 37436 36258 37492 36270
rect 37436 36206 37438 36258
rect 37490 36206 37492 36258
rect 37212 36194 37268 36204
rect 37436 35810 37492 36206
rect 37996 36260 38052 36270
rect 37996 36166 38052 36204
rect 37436 35758 37438 35810
rect 37490 35758 37492 35810
rect 37436 35746 37492 35758
rect 37100 35698 37156 35710
rect 37100 35646 37102 35698
rect 37154 35646 37156 35698
rect 37100 35138 37156 35646
rect 37548 35698 37604 35710
rect 37548 35646 37550 35698
rect 37602 35646 37604 35698
rect 37212 35588 37268 35598
rect 37212 35494 37268 35532
rect 37548 35588 37604 35646
rect 38108 35700 38164 35710
rect 38108 35606 38164 35644
rect 37100 35086 37102 35138
rect 37154 35086 37156 35138
rect 37100 35074 37156 35086
rect 37100 34916 37156 34926
rect 37100 34802 37156 34860
rect 37100 34750 37102 34802
rect 37154 34750 37156 34802
rect 37100 34738 37156 34750
rect 37212 34802 37268 34814
rect 37212 34750 37214 34802
rect 37266 34750 37268 34802
rect 37212 32004 37268 34750
rect 37212 31938 37268 31948
rect 37212 31668 37268 31678
rect 37212 31574 37268 31612
rect 36988 30118 37044 30156
rect 37100 31554 37156 31566
rect 37100 31502 37102 31554
rect 37154 31502 37156 31554
rect 37100 30100 37156 31502
rect 37100 30006 37156 30044
rect 37324 29986 37380 29998
rect 37324 29934 37326 29986
rect 37378 29934 37380 29986
rect 37100 28644 37156 28654
rect 36988 28588 37100 28644
rect 36988 28530 37044 28588
rect 37100 28578 37156 28588
rect 37324 28642 37380 29934
rect 37324 28590 37326 28642
rect 37378 28590 37380 28642
rect 37324 28578 37380 28590
rect 37548 28756 37604 35532
rect 38220 34692 38276 38780
rect 38780 38724 38836 38734
rect 38892 38724 38948 39340
rect 38836 38668 38948 38724
rect 38780 35700 38836 38668
rect 39228 37940 39284 39678
rect 39900 38948 39956 38958
rect 39900 38854 39956 38892
rect 39788 38834 39844 38846
rect 39788 38782 39790 38834
rect 39842 38782 39844 38834
rect 39788 37940 39844 38782
rect 40124 38836 40180 38846
rect 40124 38742 40180 38780
rect 40348 38164 40404 41918
rect 41132 41860 41188 41870
rect 41132 41766 41188 41804
rect 43596 41300 43652 41310
rect 43708 41300 43764 45200
rect 43596 41298 43764 41300
rect 43596 41246 43598 41298
rect 43650 41246 43764 41298
rect 43596 41244 43764 41246
rect 43596 41234 43652 41244
rect 41580 41186 41636 41198
rect 41580 41134 41582 41186
rect 41634 41134 41636 41186
rect 40460 40404 40516 40414
rect 41020 40404 41076 40414
rect 40460 40402 41076 40404
rect 40460 40350 40462 40402
rect 40514 40350 41022 40402
rect 41074 40350 41076 40402
rect 40460 40348 41076 40350
rect 40460 39396 40516 40348
rect 41020 40338 41076 40348
rect 41580 40292 41636 41134
rect 41356 39508 41412 39518
rect 41356 39506 41524 39508
rect 41356 39454 41358 39506
rect 41410 39454 41524 39506
rect 41356 39452 41524 39454
rect 41356 39442 41412 39452
rect 40460 39330 40516 39340
rect 40908 39060 40964 39070
rect 40796 38836 40852 38846
rect 40572 38834 40852 38836
rect 40572 38782 40798 38834
rect 40850 38782 40852 38834
rect 40572 38780 40852 38782
rect 40348 38108 40516 38164
rect 40236 37940 40292 37950
rect 39788 37938 40292 37940
rect 39788 37886 40238 37938
rect 40290 37886 40292 37938
rect 39788 37884 40292 37886
rect 39228 37874 39284 37884
rect 38780 35634 38836 35644
rect 39340 37044 39396 37054
rect 38220 34626 38276 34636
rect 37884 32450 37940 32462
rect 37884 32398 37886 32450
rect 37938 32398 37940 32450
rect 37884 30100 37940 32398
rect 37884 30034 37940 30044
rect 38108 31892 38164 31902
rect 37548 28642 37604 28700
rect 37548 28590 37550 28642
rect 37602 28590 37604 28642
rect 37548 28578 37604 28590
rect 37772 28644 37828 28654
rect 37772 28550 37828 28588
rect 36988 28478 36990 28530
rect 37042 28478 37044 28530
rect 36988 28466 37044 28478
rect 38108 28530 38164 31836
rect 39340 31668 39396 36988
rect 40236 37044 40292 37884
rect 40348 37940 40404 37950
rect 40348 37846 40404 37884
rect 40236 36978 40292 36988
rect 40460 36820 40516 38108
rect 40572 38050 40628 38780
rect 40796 38770 40852 38780
rect 40572 37998 40574 38050
rect 40626 37998 40628 38050
rect 40572 37986 40628 37998
rect 40348 36764 40516 36820
rect 40012 36260 40068 36270
rect 40012 35810 40068 36204
rect 40012 35758 40014 35810
rect 40066 35758 40068 35810
rect 40012 35746 40068 35758
rect 39452 35700 39508 35710
rect 39452 35606 39508 35644
rect 39788 35698 39844 35710
rect 39788 35646 39790 35698
rect 39842 35646 39844 35698
rect 39788 35588 39844 35646
rect 39788 35522 39844 35532
rect 40236 35588 40292 35598
rect 40236 35494 40292 35532
rect 40348 35140 40404 36764
rect 40796 36708 40852 36718
rect 40460 36706 40852 36708
rect 40460 36654 40798 36706
rect 40850 36654 40852 36706
rect 40460 36652 40852 36654
rect 40460 35698 40516 36652
rect 40796 36642 40852 36652
rect 40684 36372 40740 36382
rect 40460 35646 40462 35698
rect 40514 35646 40516 35698
rect 40460 35634 40516 35646
rect 40572 36370 40740 36372
rect 40572 36318 40686 36370
rect 40738 36318 40740 36370
rect 40572 36316 40740 36318
rect 40348 35074 40404 35084
rect 40572 34916 40628 36316
rect 40684 36306 40740 36316
rect 40796 36260 40852 36270
rect 40796 36166 40852 36204
rect 40236 34860 40628 34916
rect 40684 36148 40740 36158
rect 40236 34468 40292 34860
rect 40684 34802 40740 36092
rect 40908 35924 40964 39004
rect 41356 39060 41412 39070
rect 41356 38966 41412 39004
rect 41468 39058 41524 39452
rect 41468 39006 41470 39058
rect 41522 39006 41524 39058
rect 41468 38994 41524 39006
rect 41580 38948 41636 40236
rect 41804 40290 41860 40302
rect 41804 40238 41806 40290
rect 41858 40238 41860 40290
rect 41692 39060 41748 39070
rect 41692 38966 41748 39004
rect 41580 38882 41636 38892
rect 41132 38836 41188 38846
rect 41132 38834 41300 38836
rect 41132 38782 41134 38834
rect 41186 38782 41300 38834
rect 41132 38780 41300 38782
rect 41132 38770 41188 38780
rect 41020 37938 41076 37950
rect 41020 37886 41022 37938
rect 41074 37886 41076 37938
rect 41020 37266 41076 37886
rect 41132 37940 41188 37950
rect 41132 37846 41188 37884
rect 41244 37492 41300 38780
rect 41804 38722 41860 40238
rect 43932 40292 43988 40302
rect 43932 40198 43988 40236
rect 42028 39618 42084 39630
rect 42028 39566 42030 39618
rect 42082 39566 42084 39618
rect 42028 39396 42084 39566
rect 42028 39330 42084 39340
rect 41804 38670 41806 38722
rect 41858 38670 41860 38722
rect 41804 38658 41860 38670
rect 41916 38834 41972 38846
rect 41916 38782 41918 38834
rect 41970 38782 41972 38834
rect 41916 38388 41972 38782
rect 42140 38836 42196 38846
rect 42140 38742 42196 38780
rect 41692 38332 41972 38388
rect 41356 37940 41412 37950
rect 41692 37940 41748 38332
rect 41356 37938 41748 37940
rect 41356 37886 41358 37938
rect 41410 37886 41748 37938
rect 41356 37884 41748 37886
rect 41356 37874 41412 37884
rect 41356 37492 41412 37502
rect 41244 37490 41412 37492
rect 41244 37438 41358 37490
rect 41410 37438 41412 37490
rect 41244 37436 41412 37438
rect 41356 37426 41412 37436
rect 41020 37214 41022 37266
rect 41074 37214 41076 37266
rect 41020 36148 41076 37214
rect 41132 37378 41188 37390
rect 41132 37326 41134 37378
rect 41186 37326 41188 37378
rect 41132 36260 41188 37326
rect 41132 36194 41188 36204
rect 43820 36260 43876 36270
rect 41020 36082 41076 36092
rect 40908 35868 41076 35924
rect 40684 34750 40686 34802
rect 40738 34750 40740 34802
rect 40348 34692 40404 34702
rect 40572 34692 40628 34702
rect 40348 34598 40404 34636
rect 40460 34690 40628 34692
rect 40460 34638 40574 34690
rect 40626 34638 40628 34690
rect 40460 34636 40628 34638
rect 40236 34412 40404 34468
rect 40012 33348 40068 33358
rect 40012 33254 40068 33292
rect 40348 33346 40404 34412
rect 40348 33294 40350 33346
rect 40402 33294 40404 33346
rect 39340 31218 39396 31612
rect 39340 31166 39342 31218
rect 39394 31166 39396 31218
rect 39340 31154 39396 31166
rect 39564 31892 39620 31902
rect 39004 30994 39060 31006
rect 39004 30942 39006 30994
rect 39058 30942 39060 30994
rect 38668 30882 38724 30894
rect 38668 30830 38670 30882
rect 38722 30830 38724 30882
rect 38668 29988 38724 30830
rect 38892 29988 38948 29998
rect 39004 29988 39060 30942
rect 39564 30098 39620 31836
rect 40348 31892 40404 33294
rect 40460 33460 40516 34636
rect 40572 34626 40628 34636
rect 40684 34468 40740 34750
rect 40460 33234 40516 33404
rect 40460 33182 40462 33234
rect 40514 33182 40516 33234
rect 40460 33170 40516 33182
rect 40572 34412 40740 34468
rect 40908 35700 40964 35710
rect 40348 31826 40404 31836
rect 40572 31668 40628 34412
rect 40908 33348 40964 35644
rect 40684 33124 40740 33134
rect 40684 33122 40852 33124
rect 40684 33070 40686 33122
rect 40738 33070 40852 33122
rect 40684 33068 40852 33070
rect 40684 33058 40740 33068
rect 40796 32674 40852 33068
rect 40796 32622 40798 32674
rect 40850 32622 40852 32674
rect 40796 32610 40852 32622
rect 40348 31612 40572 31668
rect 40348 31218 40404 31612
rect 40572 31602 40628 31612
rect 40348 31166 40350 31218
rect 40402 31166 40404 31218
rect 40348 31154 40404 31166
rect 40012 30996 40068 31006
rect 39564 30046 39566 30098
rect 39618 30046 39620 30098
rect 39564 30034 39620 30046
rect 39788 30994 40068 30996
rect 39788 30942 40014 30994
rect 40066 30942 40068 30994
rect 39788 30940 40068 30942
rect 39228 29988 39284 29998
rect 38668 29986 39284 29988
rect 38668 29934 38894 29986
rect 38946 29934 39230 29986
rect 39282 29934 39284 29986
rect 38668 29932 39284 29934
rect 38556 29428 38612 29438
rect 38556 29316 38612 29372
rect 38108 28478 38110 28530
rect 38162 28478 38164 28530
rect 38108 28466 38164 28478
rect 38220 29314 38612 29316
rect 38220 29262 38558 29314
rect 38610 29262 38612 29314
rect 38220 29260 38612 29262
rect 36092 28420 36148 28430
rect 35756 27748 35812 27758
rect 35756 27076 35812 27692
rect 35756 26982 35812 27020
rect 36092 26962 36148 28364
rect 37100 28418 37156 28430
rect 37100 28366 37102 28418
rect 37154 28366 37156 28418
rect 36988 27972 37044 27982
rect 37100 27972 37156 28366
rect 37996 28420 38052 28430
rect 37996 28326 38052 28364
rect 38220 28084 38276 29260
rect 38556 29250 38612 29260
rect 36988 27970 37156 27972
rect 36988 27918 36990 27970
rect 37042 27918 37156 27970
rect 36988 27916 37156 27918
rect 37772 28082 38276 28084
rect 37772 28030 38222 28082
rect 38274 28030 38276 28082
rect 37772 28028 38276 28030
rect 36988 27906 37044 27916
rect 37772 27858 37828 28028
rect 37772 27806 37774 27858
rect 37826 27806 37828 27858
rect 37772 27794 37828 27806
rect 36092 26910 36094 26962
rect 36146 26910 36148 26962
rect 35644 26516 35700 26526
rect 35532 26460 35644 26516
rect 35644 26422 35700 26460
rect 35420 26292 35476 26302
rect 35420 26290 35588 26292
rect 35420 26238 35422 26290
rect 35474 26238 35588 26290
rect 35420 26236 35588 26238
rect 35420 26226 35476 26236
rect 34860 25956 34916 25966
rect 34300 22258 34356 22270
rect 34300 22206 34302 22258
rect 34354 22206 34356 22258
rect 34300 21812 34356 22206
rect 34300 21746 34356 21756
rect 34860 18676 34916 25900
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 24948 35588 26236
rect 35532 24882 35588 24892
rect 35644 25284 35700 25294
rect 35644 24948 35700 25228
rect 35644 24946 35924 24948
rect 35644 24894 35646 24946
rect 35698 24894 35924 24946
rect 35644 24892 35924 24894
rect 35644 24882 35700 24892
rect 35868 24834 35924 24892
rect 35868 24782 35870 24834
rect 35922 24782 35924 24834
rect 35868 24770 35924 24782
rect 35980 24836 36036 24846
rect 36092 24836 36148 26910
rect 37436 27076 37492 27086
rect 35980 24834 36148 24836
rect 35980 24782 35982 24834
rect 36034 24782 36148 24834
rect 35980 24780 36148 24782
rect 35980 24770 36036 24780
rect 36092 24500 36148 24780
rect 36428 26516 36484 26526
rect 35980 24444 36148 24500
rect 36204 24722 36260 24734
rect 36204 24670 36206 24722
rect 36258 24670 36260 24722
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35980 23548 36036 24444
rect 35868 23492 36036 23548
rect 36092 23716 36148 23726
rect 35308 23268 35364 23278
rect 35308 23156 35364 23212
rect 35644 23156 35700 23166
rect 35308 23100 35644 23156
rect 35644 23062 35700 23100
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35420 22596 35476 22606
rect 35308 21812 35364 21822
rect 35308 21718 35364 21756
rect 35420 21698 35476 22540
rect 35868 22260 35924 23492
rect 36092 23266 36148 23660
rect 36204 23492 36260 24670
rect 36204 23426 36260 23436
rect 36092 23214 36094 23266
rect 36146 23214 36148 23266
rect 36092 23202 36148 23214
rect 36204 23266 36260 23278
rect 36204 23214 36206 23266
rect 36258 23214 36260 23266
rect 36092 23042 36148 23054
rect 36092 22990 36094 23042
rect 36146 22990 36148 23042
rect 36092 22596 36148 22990
rect 36092 22530 36148 22540
rect 36204 22484 36260 23214
rect 36428 23156 36484 26460
rect 37436 25506 37492 27020
rect 37884 25620 37940 25630
rect 37884 25526 37940 25564
rect 38220 25620 38276 28028
rect 38668 27748 38724 27758
rect 38668 27654 38724 27692
rect 38220 25554 38276 25564
rect 38668 25620 38724 25630
rect 37436 25454 37438 25506
rect 37490 25454 37492 25506
rect 37436 25442 37492 25454
rect 36988 25396 37044 25406
rect 36652 25394 37044 25396
rect 36652 25342 36990 25394
rect 37042 25342 37044 25394
rect 36652 25340 37044 25342
rect 36540 24948 36596 24958
rect 36540 24854 36596 24892
rect 36652 24834 36708 25340
rect 36988 25330 37044 25340
rect 36652 24782 36654 24834
rect 36706 24782 36708 24834
rect 36652 24770 36708 24782
rect 36540 24498 36596 24510
rect 36540 24446 36542 24498
rect 36594 24446 36596 24498
rect 36540 23716 36596 24446
rect 38668 24052 38724 25564
rect 38780 24612 38836 29932
rect 38892 29922 38948 29932
rect 39228 29922 39284 29932
rect 39788 29540 39844 30940
rect 40012 30930 40068 30940
rect 39004 28756 39060 28766
rect 39004 28082 39060 28700
rect 39004 28030 39006 28082
rect 39058 28030 39060 28082
rect 39004 28018 39060 28030
rect 39340 27858 39396 27870
rect 39340 27806 39342 27858
rect 39394 27806 39396 27858
rect 39340 27748 39396 27806
rect 39228 24834 39284 24846
rect 39228 24782 39230 24834
rect 39282 24782 39284 24834
rect 39116 24722 39172 24734
rect 39116 24670 39118 24722
rect 39170 24670 39172 24722
rect 39116 24612 39172 24670
rect 39228 24724 39284 24782
rect 39228 24658 39284 24668
rect 38780 24610 39172 24612
rect 38780 24558 38782 24610
rect 38834 24558 39172 24610
rect 38780 24556 39172 24558
rect 38780 24546 38836 24556
rect 38668 24050 38948 24052
rect 38668 23998 38670 24050
rect 38722 23998 38948 24050
rect 38668 23996 38948 23998
rect 38668 23986 38724 23996
rect 38892 23938 38948 23996
rect 38892 23886 38894 23938
rect 38946 23886 38948 23938
rect 38892 23874 38948 23886
rect 36540 23650 36596 23660
rect 37212 23156 37268 23166
rect 36428 23154 36596 23156
rect 36428 23102 36430 23154
rect 36482 23102 36596 23154
rect 36428 23100 36596 23102
rect 36428 23090 36484 23100
rect 36428 22484 36484 22494
rect 36204 22482 36484 22484
rect 36204 22430 36430 22482
rect 36482 22430 36484 22482
rect 36204 22428 36484 22430
rect 35868 22204 36036 22260
rect 35420 21646 35422 21698
rect 35474 21646 35476 21698
rect 35420 21634 35476 21646
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35980 20802 36036 22204
rect 36204 20914 36260 22428
rect 36428 22418 36484 22428
rect 36204 20862 36206 20914
rect 36258 20862 36260 20914
rect 36204 20850 36260 20862
rect 36316 20914 36372 20926
rect 36316 20862 36318 20914
rect 36370 20862 36372 20914
rect 35980 20750 35982 20802
rect 36034 20750 36036 20802
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35644 19012 35700 19022
rect 35196 18676 35252 18686
rect 35644 18676 35700 18956
rect 34860 18674 35700 18676
rect 34860 18622 34862 18674
rect 34914 18622 35198 18674
rect 35250 18622 35700 18674
rect 34860 18620 35700 18622
rect 35868 19010 35924 19022
rect 35868 18958 35870 19010
rect 35922 18958 35924 19010
rect 34860 18610 34916 18620
rect 35196 18610 35252 18620
rect 35756 18564 35812 18574
rect 35308 18452 35364 18462
rect 35644 18452 35700 18462
rect 35308 18450 35700 18452
rect 35308 18398 35310 18450
rect 35362 18398 35646 18450
rect 35698 18398 35700 18450
rect 35308 18396 35700 18398
rect 35308 18386 35364 18396
rect 35644 18386 35700 18396
rect 35196 18228 35252 18238
rect 35196 18226 35588 18228
rect 35196 18174 35198 18226
rect 35250 18174 35588 18226
rect 35196 18172 35588 18174
rect 35196 18162 35252 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 34860 17780 34916 17790
rect 35196 17780 35252 17790
rect 34860 17778 35252 17780
rect 34860 17726 34862 17778
rect 34914 17726 35198 17778
rect 35250 17726 35252 17778
rect 34860 17724 35252 17726
rect 34860 17714 34916 17724
rect 35196 17714 35252 17724
rect 35308 17668 35364 17678
rect 35308 17556 35364 17612
rect 35532 17666 35588 18172
rect 35532 17614 35534 17666
rect 35586 17614 35588 17666
rect 35532 17602 35588 17614
rect 35084 17500 35364 17556
rect 35756 17554 35812 18508
rect 35868 17668 35924 18958
rect 35980 18452 36036 20750
rect 36204 19236 36260 19246
rect 36316 19236 36372 20862
rect 36204 19234 36372 19236
rect 36204 19182 36206 19234
rect 36258 19182 36372 19234
rect 36204 19180 36372 19182
rect 36204 19170 36260 19180
rect 36092 19012 36148 19022
rect 36092 18918 36148 18956
rect 36092 18452 36148 18462
rect 35980 18450 36148 18452
rect 35980 18398 36094 18450
rect 36146 18398 36148 18450
rect 35980 18396 36148 18398
rect 36092 18386 36148 18396
rect 36428 18452 36484 18462
rect 36428 18338 36484 18396
rect 36428 18286 36430 18338
rect 36482 18286 36484 18338
rect 36428 18274 36484 18286
rect 36428 17780 36484 17790
rect 36428 17686 36484 17724
rect 35868 17602 35924 17612
rect 35756 17502 35758 17554
rect 35810 17502 35812 17554
rect 34748 17444 34804 17454
rect 34300 17442 34804 17444
rect 34300 17390 34750 17442
rect 34802 17390 34804 17442
rect 34300 17388 34804 17390
rect 34300 16210 34356 17388
rect 34748 17378 34804 17388
rect 34300 16158 34302 16210
rect 34354 16158 34356 16210
rect 34300 16146 34356 16158
rect 34188 14028 34468 14084
rect 34412 13972 34468 14028
rect 34412 13970 34804 13972
rect 34412 13918 34414 13970
rect 34466 13918 34804 13970
rect 34412 13916 34804 13918
rect 34412 13906 34468 13916
rect 30828 12962 30996 12964
rect 30828 12910 30830 12962
rect 30882 12910 30996 12962
rect 30828 12908 30996 12910
rect 30828 12898 30884 12908
rect 30268 12852 30324 12862
rect 30268 12758 30324 12796
rect 30604 12850 30660 12862
rect 30604 12798 30606 12850
rect 30658 12798 30660 12850
rect 30604 12404 30660 12798
rect 30604 12338 30660 12348
rect 30940 12068 30996 12908
rect 31948 12852 32004 12862
rect 31388 12180 31444 12190
rect 31388 12086 31444 12124
rect 29932 11566 29934 11618
rect 29986 11566 29988 11618
rect 29932 11554 29988 11566
rect 30716 12066 30996 12068
rect 30716 12014 30942 12066
rect 30994 12014 30996 12066
rect 30716 12012 30996 12014
rect 30716 11394 30772 12012
rect 30940 12002 30996 12012
rect 30716 11342 30718 11394
rect 30770 11342 30772 11394
rect 30716 11330 30772 11342
rect 30380 11284 30436 11294
rect 30268 11282 30436 11284
rect 30268 11230 30382 11282
rect 30434 11230 30436 11282
rect 30268 11228 30436 11230
rect 30044 10612 30100 10622
rect 30268 10612 30324 11228
rect 30380 11218 30436 11228
rect 30492 11284 30548 11294
rect 30492 11190 30548 11228
rect 30380 10724 30436 10734
rect 30380 10630 30436 10668
rect 31948 10724 32004 12796
rect 32844 12852 32900 12862
rect 32060 12404 32116 12414
rect 32060 11284 32116 12348
rect 32060 11218 32116 11228
rect 32396 12068 32452 12078
rect 31948 10658 32004 10668
rect 30100 10556 30324 10612
rect 30044 10518 30100 10556
rect 29820 9998 29822 10050
rect 29874 9998 29876 10050
rect 29820 9986 29876 9998
rect 29372 9828 29428 9838
rect 29372 9734 29428 9772
rect 28924 9214 28926 9266
rect 28978 9214 28980 9266
rect 28924 9202 28980 9214
rect 29932 9714 29988 9726
rect 29932 9662 29934 9714
rect 29986 9662 29988 9714
rect 27580 9156 27636 9166
rect 27580 9062 27636 9100
rect 28364 9156 28420 9166
rect 28364 9062 28420 9100
rect 27804 9044 27860 9054
rect 28252 9044 28308 9054
rect 27804 9042 28308 9044
rect 27804 8990 27806 9042
rect 27858 8990 28254 9042
rect 28306 8990 28308 9042
rect 27804 8988 28308 8990
rect 27804 8978 27860 8988
rect 27244 8876 27524 8932
rect 27132 8642 27188 8652
rect 27020 8428 27412 8484
rect 27356 6692 27412 8428
rect 27468 7700 27524 8876
rect 27580 8708 27636 8718
rect 27580 8146 27636 8652
rect 28252 8372 28308 8988
rect 27580 8094 27582 8146
rect 27634 8094 27636 8146
rect 27580 8082 27636 8094
rect 27804 8260 27860 8270
rect 27580 7700 27636 7710
rect 27468 7698 27636 7700
rect 27468 7646 27582 7698
rect 27634 7646 27636 7698
rect 27468 7644 27636 7646
rect 27580 7634 27636 7644
rect 27692 7474 27748 7486
rect 27692 7422 27694 7474
rect 27746 7422 27748 7474
rect 27468 6692 27524 6702
rect 26908 6636 27076 6692
rect 26572 6466 26628 6478
rect 26572 6414 26574 6466
rect 26626 6414 26628 6466
rect 26572 6356 26628 6414
rect 26684 6356 26740 6636
rect 26796 6626 26852 6636
rect 26908 6356 26964 6366
rect 26684 6300 26852 6356
rect 26572 6290 26628 6300
rect 26460 5926 26516 5964
rect 26348 5684 26404 5694
rect 26124 5682 26404 5684
rect 26124 5630 26350 5682
rect 26402 5630 26404 5682
rect 26124 5628 26404 5630
rect 26348 5460 26404 5628
rect 26796 5460 26852 6300
rect 26908 5684 26964 6300
rect 26908 5618 26964 5628
rect 26348 5404 26852 5460
rect 24556 5182 24558 5234
rect 24610 5182 24612 5234
rect 24556 5170 24612 5182
rect 22764 4398 22766 4450
rect 22818 4398 22820 4450
rect 22764 4386 22820 4398
rect 27020 4564 27076 6636
rect 27244 6690 27524 6692
rect 27244 6638 27470 6690
rect 27522 6638 27524 6690
rect 27244 6636 27524 6638
rect 27132 6580 27188 6590
rect 27132 6486 27188 6524
rect 27132 6020 27188 6030
rect 27244 6020 27300 6636
rect 27468 6626 27524 6636
rect 27580 6468 27636 6478
rect 27692 6468 27748 7422
rect 27804 6916 27860 8204
rect 28252 7474 28308 8316
rect 28476 9042 28532 9054
rect 28476 8990 28478 9042
rect 28530 8990 28532 9042
rect 28476 8260 28532 8990
rect 28476 8194 28532 8204
rect 28700 9044 28756 9054
rect 28700 7586 28756 8988
rect 29484 8372 29540 8382
rect 29484 8278 29540 8316
rect 29932 8372 29988 9662
rect 29932 8306 29988 8316
rect 31612 8372 31668 8382
rect 31612 8278 31668 8316
rect 32396 8260 32452 12012
rect 32508 11396 32564 11406
rect 32508 11302 32564 11340
rect 32844 11394 32900 12796
rect 32956 12068 33012 12908
rect 33292 12962 33348 12974
rect 33292 12910 33294 12962
rect 33346 12910 33348 12962
rect 33180 12850 33236 12862
rect 33180 12798 33182 12850
rect 33234 12798 33236 12850
rect 33068 12740 33124 12750
rect 33068 12646 33124 12684
rect 33068 12404 33124 12414
rect 33180 12404 33236 12798
rect 33124 12348 33236 12404
rect 33068 12338 33124 12348
rect 33068 12068 33124 12078
rect 32956 12066 33124 12068
rect 32956 12014 33070 12066
rect 33122 12014 33124 12066
rect 32956 12012 33124 12014
rect 33068 12002 33124 12012
rect 33292 11732 33348 12910
rect 33964 12964 34020 12974
rect 33964 12870 34020 12908
rect 34748 12962 34804 13916
rect 34748 12910 34750 12962
rect 34802 12910 34804 12962
rect 33740 12738 33796 12750
rect 33740 12686 33742 12738
rect 33794 12686 33796 12738
rect 33740 12404 33796 12686
rect 33740 12338 33796 12348
rect 32956 11676 33348 11732
rect 32956 11506 33012 11676
rect 32956 11454 32958 11506
rect 33010 11454 33012 11506
rect 32956 11442 33012 11454
rect 32844 11342 32846 11394
rect 32898 11342 32900 11394
rect 32844 11330 32900 11342
rect 33516 11396 33572 11406
rect 33516 11302 33572 11340
rect 34748 11396 34804 12910
rect 34748 11330 34804 11340
rect 35084 13076 35140 17500
rect 35756 17220 35812 17502
rect 35980 17556 36036 17566
rect 35980 17462 36036 17500
rect 36540 17556 36596 23100
rect 36540 17490 36596 17500
rect 36764 22372 36820 22382
rect 35756 17164 36484 17220
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 36428 16210 36484 17164
rect 36764 16996 36820 22316
rect 37100 22372 37156 22382
rect 37100 22278 37156 22316
rect 37212 18452 37268 23100
rect 39004 22932 39060 24556
rect 39228 24498 39284 24510
rect 39228 24446 39230 24498
rect 39282 24446 39284 24498
rect 39228 23154 39284 24446
rect 39228 23102 39230 23154
rect 39282 23102 39284 23154
rect 39228 23090 39284 23102
rect 39004 22866 39060 22876
rect 39116 20468 39172 20478
rect 39340 20468 39396 27692
rect 39788 24948 39844 29484
rect 40348 29428 40404 29438
rect 40908 29428 40964 33292
rect 41020 32900 41076 35868
rect 41692 35588 41748 35598
rect 41692 35494 41748 35532
rect 43820 35586 43876 36204
rect 43820 35534 43822 35586
rect 43874 35534 43876 35586
rect 43820 35522 43876 35534
rect 43820 33460 43876 33470
rect 43820 33366 43876 33404
rect 41692 33236 41748 33246
rect 41692 33234 41860 33236
rect 41692 33182 41694 33234
rect 41746 33182 41860 33234
rect 41692 33180 41860 33182
rect 41692 33170 41748 33180
rect 41020 32834 41076 32844
rect 41692 32788 41748 32798
rect 41692 32694 41748 32732
rect 41804 32786 41860 33180
rect 41804 32734 41806 32786
rect 41858 32734 41860 32786
rect 41804 32722 41860 32734
rect 41020 32676 41076 32686
rect 41020 32674 41188 32676
rect 41020 32622 41022 32674
rect 41074 32622 41188 32674
rect 41020 32620 41188 32622
rect 41020 32610 41076 32620
rect 41132 32562 41188 32620
rect 41132 32510 41134 32562
rect 41186 32510 41188 32562
rect 41132 32498 41188 32510
rect 41468 32564 41524 32574
rect 41468 32562 41636 32564
rect 41468 32510 41470 32562
rect 41522 32510 41636 32562
rect 41468 32508 41636 32510
rect 41468 32498 41524 32508
rect 41580 32004 41636 32508
rect 41692 32004 41748 32014
rect 41580 32002 41748 32004
rect 41580 31950 41694 32002
rect 41746 31950 41748 32002
rect 41580 31948 41748 31950
rect 41692 31938 41748 31948
rect 41580 31668 41636 31678
rect 41580 31574 41636 31612
rect 41692 31554 41748 31566
rect 41692 31502 41694 31554
rect 41746 31502 41748 31554
rect 41692 29764 41748 31502
rect 41692 29698 41748 29708
rect 42476 29764 42532 29774
rect 42532 29708 42644 29764
rect 42476 29698 42532 29708
rect 40404 29426 40964 29428
rect 40404 29374 40910 29426
rect 40962 29374 40964 29426
rect 40404 29372 40964 29374
rect 40348 29334 40404 29372
rect 40908 29362 40964 29372
rect 41692 29316 41748 29326
rect 42588 29316 42644 29708
rect 41692 29314 41972 29316
rect 41692 29262 41694 29314
rect 41746 29262 41972 29314
rect 41692 29260 41972 29262
rect 41692 29250 41748 29260
rect 41468 28756 41524 28766
rect 41468 28642 41524 28700
rect 41916 28754 41972 29260
rect 42476 28866 42532 28878
rect 42476 28814 42478 28866
rect 42530 28814 42532 28866
rect 42476 28756 42532 28814
rect 41916 28702 41918 28754
rect 41970 28702 41972 28754
rect 41916 28690 41972 28702
rect 42252 28700 42532 28756
rect 41468 28590 41470 28642
rect 41522 28590 41524 28642
rect 41468 28578 41524 28590
rect 42140 28644 42196 28654
rect 42252 28644 42308 28700
rect 42140 28642 42308 28644
rect 42140 28590 42142 28642
rect 42194 28590 42308 28642
rect 42140 28588 42308 28590
rect 42140 28578 42196 28588
rect 40572 28532 40628 28542
rect 40236 25620 40292 25630
rect 40236 25526 40292 25564
rect 39788 24722 39844 24892
rect 40572 25506 40628 28476
rect 41692 28530 41748 28542
rect 41692 28478 41694 28530
rect 41746 28478 41748 28530
rect 41132 25620 41188 25630
rect 40572 25454 40574 25506
rect 40626 25454 40628 25506
rect 40012 24836 40068 24846
rect 40012 24742 40068 24780
rect 39788 24670 39790 24722
rect 39842 24670 39844 24722
rect 39788 24658 39844 24670
rect 39900 24164 39956 24174
rect 39676 23826 39732 23838
rect 39676 23774 39678 23826
rect 39730 23774 39732 23826
rect 39564 23380 39620 23390
rect 39676 23380 39732 23774
rect 39564 23378 39732 23380
rect 39564 23326 39566 23378
rect 39618 23326 39732 23378
rect 39564 23324 39732 23326
rect 39564 23314 39620 23324
rect 39900 23266 39956 24108
rect 39900 23214 39902 23266
rect 39954 23214 39956 23266
rect 39676 23156 39732 23166
rect 39676 23062 39732 23100
rect 39172 20412 39396 20468
rect 39116 20132 39172 20412
rect 39452 20132 39508 20142
rect 39116 20130 39508 20132
rect 39116 20078 39118 20130
rect 39170 20078 39454 20130
rect 39506 20078 39508 20130
rect 39116 20076 39508 20078
rect 39116 20066 39172 20076
rect 39452 20066 39508 20076
rect 39564 20132 39620 20142
rect 38892 19124 38948 19134
rect 39228 19124 39284 19134
rect 38948 19122 39284 19124
rect 38948 19070 39230 19122
rect 39282 19070 39284 19122
rect 38948 19068 39284 19070
rect 38892 19030 38948 19068
rect 39228 19058 39284 19068
rect 39564 19122 39620 20076
rect 39788 20132 39844 20142
rect 39900 20132 39956 23214
rect 39788 20130 39956 20132
rect 39788 20078 39790 20130
rect 39842 20078 39956 20130
rect 39788 20076 39956 20078
rect 39788 20066 39844 20076
rect 39564 19070 39566 19122
rect 39618 19070 39620 19122
rect 39564 19058 39620 19070
rect 39900 19124 39956 20076
rect 40572 20132 40628 25454
rect 40684 25508 40740 25518
rect 40684 25394 40740 25452
rect 41132 25506 41188 25564
rect 41132 25454 41134 25506
rect 41186 25454 41188 25506
rect 41132 25442 41188 25454
rect 40684 25342 40686 25394
rect 40738 25342 40740 25394
rect 40684 25330 40740 25342
rect 40908 25282 40964 25294
rect 40908 25230 40910 25282
rect 40962 25230 40964 25282
rect 40908 24724 40964 25230
rect 41468 24724 41524 24734
rect 40908 24722 41524 24724
rect 40908 24670 41470 24722
rect 41522 24670 41524 24722
rect 40908 24668 41524 24670
rect 41468 24658 41524 24668
rect 41692 21028 41748 28478
rect 42364 28532 42420 28542
rect 42364 28438 42420 28476
rect 42476 28532 42532 28542
rect 42588 28532 42644 29260
rect 43820 29316 43876 29326
rect 43820 29222 43876 29260
rect 42476 28530 42644 28532
rect 42476 28478 42478 28530
rect 42530 28478 42644 28530
rect 42476 28476 42644 28478
rect 42476 28466 42532 28476
rect 44044 25620 44100 25630
rect 44044 25526 44100 25564
rect 41916 25394 41972 25406
rect 41916 25342 41918 25394
rect 41970 25342 41972 25394
rect 41804 24948 41860 24958
rect 41916 24948 41972 25342
rect 41804 24946 41972 24948
rect 41804 24894 41806 24946
rect 41858 24894 41972 24946
rect 41804 24892 41972 24894
rect 41804 24882 41860 24892
rect 42364 24836 42420 24846
rect 41804 24724 41860 24734
rect 41804 24050 41860 24668
rect 41804 23998 41806 24050
rect 41858 23998 41860 24050
rect 41804 23716 41860 23998
rect 41916 24722 41972 24734
rect 41916 24670 41918 24722
rect 41970 24670 41972 24722
rect 41916 23940 41972 24670
rect 42028 24722 42084 24734
rect 42028 24670 42030 24722
rect 42082 24670 42084 24722
rect 42028 24164 42084 24670
rect 42028 24098 42084 24108
rect 42028 23940 42084 23950
rect 41916 23938 42084 23940
rect 41916 23886 42030 23938
rect 42082 23886 42084 23938
rect 41916 23884 42084 23886
rect 42028 23874 42084 23884
rect 42364 23938 42420 24780
rect 42364 23886 42366 23938
rect 42418 23886 42420 23938
rect 42252 23716 42308 23726
rect 41804 23714 42308 23716
rect 41804 23662 42254 23714
rect 42306 23662 42308 23714
rect 41804 23660 42308 23662
rect 42252 23650 42308 23660
rect 42364 23548 42420 23886
rect 41916 23492 42420 23548
rect 41804 21028 41860 21038
rect 41692 21026 41860 21028
rect 41692 20974 41806 21026
rect 41858 20974 41860 21026
rect 41692 20972 41860 20974
rect 41804 20962 41860 20972
rect 41916 20804 41972 23492
rect 41692 20802 41972 20804
rect 41692 20750 41918 20802
rect 41970 20750 41972 20802
rect 41692 20748 41972 20750
rect 41692 20188 41748 20748
rect 41916 20738 41972 20748
rect 40572 20066 40628 20076
rect 41244 20132 41748 20188
rect 41804 20578 41860 20590
rect 41804 20526 41806 20578
rect 41858 20526 41860 20578
rect 41132 20018 41188 20030
rect 41132 19966 41134 20018
rect 41186 19966 41188 20018
rect 39900 19058 39956 19068
rect 40348 19908 40404 19918
rect 41132 19908 41188 19966
rect 40348 19906 41188 19908
rect 40348 19854 40350 19906
rect 40402 19854 41188 19906
rect 40348 19852 41188 19854
rect 40348 18676 40404 19852
rect 41244 19348 41300 20132
rect 40236 18620 40404 18676
rect 40908 19292 41300 19348
rect 41692 20020 41748 20030
rect 37212 18450 37492 18452
rect 37212 18398 37214 18450
rect 37266 18398 37492 18450
rect 37212 18396 37492 18398
rect 37212 18386 37268 18396
rect 37324 17668 37380 17678
rect 36988 17556 37044 17566
rect 36988 17462 37044 17500
rect 37324 17554 37380 17612
rect 37324 17502 37326 17554
rect 37378 17502 37380 17554
rect 37324 17490 37380 17502
rect 37436 17554 37492 18396
rect 40236 17556 40292 18620
rect 40908 18564 40964 19292
rect 41692 19236 41748 19964
rect 41804 19908 41860 20526
rect 41804 19842 41860 19852
rect 41916 19906 41972 19918
rect 41916 19854 41918 19906
rect 41970 19854 41972 19906
rect 41804 19348 41860 19358
rect 41916 19348 41972 19854
rect 41804 19346 41972 19348
rect 41804 19294 41806 19346
rect 41858 19294 41972 19346
rect 41804 19292 41972 19294
rect 42364 19908 42420 19918
rect 41804 19282 41860 19292
rect 41132 19124 41188 19134
rect 41356 19124 41412 19134
rect 41580 19124 41636 19134
rect 41188 19122 41412 19124
rect 41188 19070 41358 19122
rect 41410 19070 41412 19122
rect 41188 19068 41412 19070
rect 40348 18562 40964 18564
rect 40348 18510 40910 18562
rect 40962 18510 40964 18562
rect 40348 18508 40964 18510
rect 40348 17666 40404 18508
rect 40908 18498 40964 18508
rect 41020 18564 41076 18574
rect 41020 18470 41076 18508
rect 41132 18340 41188 19068
rect 41356 19058 41412 19068
rect 41468 19122 41636 19124
rect 41468 19070 41582 19122
rect 41634 19070 41636 19122
rect 41468 19068 41636 19070
rect 41244 18676 41300 18686
rect 41468 18676 41524 19068
rect 41580 19058 41636 19068
rect 41244 18674 41524 18676
rect 41244 18622 41246 18674
rect 41298 18622 41524 18674
rect 41244 18620 41524 18622
rect 41244 18610 41300 18620
rect 41580 18562 41636 18574
rect 41580 18510 41582 18562
rect 41634 18510 41636 18562
rect 41580 18452 41636 18510
rect 41692 18562 41748 19180
rect 41916 19124 41972 19134
rect 42140 19124 42196 19134
rect 41916 19122 42196 19124
rect 41916 19070 41918 19122
rect 41970 19070 42142 19122
rect 42194 19070 42196 19122
rect 41916 19068 42196 19070
rect 41916 19058 41972 19068
rect 42140 19058 42196 19068
rect 42364 19122 42420 19852
rect 44044 19908 44100 19918
rect 44044 19814 44100 19852
rect 42476 19236 42532 19246
rect 42476 19142 42532 19180
rect 42364 19070 42366 19122
rect 42418 19070 42420 19122
rect 42364 19058 42420 19070
rect 41692 18510 41694 18562
rect 41746 18510 41748 18562
rect 41692 18498 41748 18510
rect 41580 18386 41636 18396
rect 43372 18452 43428 18462
rect 40348 17614 40350 17666
rect 40402 17614 40404 17666
rect 40348 17602 40404 17614
rect 41020 18284 41188 18340
rect 37436 17502 37438 17554
rect 37490 17502 37492 17554
rect 37436 17490 37492 17502
rect 40124 17500 40292 17556
rect 40908 17556 40964 17566
rect 41020 17556 41076 18284
rect 41580 18226 41636 18238
rect 41580 18174 41582 18226
rect 41634 18174 41636 18226
rect 41580 17666 41636 18174
rect 41580 17614 41582 17666
rect 41634 17614 41636 17666
rect 41580 17602 41636 17614
rect 40908 17554 41076 17556
rect 40908 17502 40910 17554
rect 40962 17502 41076 17554
rect 40908 17500 41076 17502
rect 41132 17554 41188 17566
rect 41132 17502 41134 17554
rect 41186 17502 41188 17554
rect 37100 17442 37156 17454
rect 37100 17390 37102 17442
rect 37154 17390 37156 17442
rect 36820 16940 36932 16996
rect 36764 16902 36820 16940
rect 36876 16772 36932 16940
rect 37100 16884 37156 17390
rect 37212 17444 37268 17454
rect 37212 17350 37268 17388
rect 37100 16828 37492 16884
rect 36876 16716 37156 16772
rect 36428 16158 36430 16210
rect 36482 16158 36484 16210
rect 36428 16146 36484 16158
rect 37100 16210 37156 16716
rect 37100 16158 37102 16210
rect 37154 16158 37156 16210
rect 37100 15876 37156 16158
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 37100 14532 37156 15820
rect 37436 15426 37492 16828
rect 40124 15876 40180 17500
rect 40908 17490 40964 17500
rect 40460 17444 40516 17454
rect 40460 16884 40516 17388
rect 40684 17442 40740 17454
rect 40684 17390 40686 17442
rect 40738 17390 40740 17442
rect 40684 17332 40740 17390
rect 41132 17332 41188 17502
rect 40684 17276 41188 17332
rect 41244 17442 41300 17454
rect 41244 17390 41246 17442
rect 41298 17390 41300 17442
rect 40124 15782 40180 15820
rect 40236 16828 40516 16884
rect 37436 15374 37438 15426
rect 37490 15374 37492 15426
rect 37436 15362 37492 15374
rect 37548 15092 37604 15102
rect 37548 15090 38164 15092
rect 37548 15038 37550 15090
rect 37602 15038 38164 15090
rect 37548 15036 38164 15038
rect 37548 15026 37604 15036
rect 38108 14642 38164 15036
rect 38108 14590 38110 14642
rect 38162 14590 38164 14642
rect 38108 14578 38164 14590
rect 40236 14642 40292 16828
rect 41244 16210 41300 17390
rect 41244 16158 41246 16210
rect 41298 16158 41300 16210
rect 41244 16146 41300 16158
rect 43372 16210 43428 18396
rect 43372 16158 43374 16210
rect 43426 16158 43428 16210
rect 43372 16146 43428 16158
rect 40460 16098 40516 16110
rect 40460 16046 40462 16098
rect 40514 16046 40516 16098
rect 40460 15876 40516 16046
rect 40460 15810 40516 15820
rect 40236 14590 40238 14642
rect 40290 14590 40292 14642
rect 40236 14578 40292 14590
rect 37324 14532 37380 14542
rect 37100 14530 37380 14532
rect 37100 14478 37326 14530
rect 37378 14478 37380 14530
rect 37100 14476 37380 14478
rect 36428 14308 36484 14318
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 13076 35252 13086
rect 35084 13074 35252 13076
rect 35084 13022 35198 13074
rect 35250 13022 35252 13074
rect 35084 13020 35252 13022
rect 33068 11284 33124 11294
rect 33068 11190 33124 11228
rect 34972 8484 35028 8494
rect 35084 8484 35140 13020
rect 35196 13010 35252 13020
rect 35196 12740 35252 12750
rect 35196 12290 35252 12684
rect 35196 12238 35198 12290
rect 35250 12238 35252 12290
rect 35196 12226 35252 12238
rect 35868 12178 35924 12190
rect 35868 12126 35870 12178
rect 35922 12126 35924 12178
rect 35868 12068 35924 12126
rect 35868 12002 35924 12012
rect 36428 12068 36484 14252
rect 37324 14308 37380 14476
rect 37324 14242 37380 14252
rect 36428 11974 36484 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35028 8428 35140 8484
rect 34972 8418 35028 8428
rect 32956 8260 33012 8270
rect 32396 8258 33012 8260
rect 32396 8206 32398 8258
rect 32450 8206 32958 8258
rect 33010 8206 33012 8258
rect 32396 8204 33012 8206
rect 32396 8194 32452 8204
rect 32956 8194 33012 8204
rect 28700 7534 28702 7586
rect 28754 7534 28756 7586
rect 28700 7522 28756 7534
rect 28252 7422 28254 7474
rect 28306 7422 28308 7474
rect 28252 7410 28308 7422
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 27804 6850 27860 6860
rect 27804 6580 27860 6590
rect 27804 6486 27860 6524
rect 27580 6466 27748 6468
rect 27580 6414 27582 6466
rect 27634 6414 27748 6466
rect 27580 6412 27748 6414
rect 27132 6018 27300 6020
rect 27132 5966 27134 6018
rect 27186 5966 27300 6018
rect 27132 5964 27300 5966
rect 27356 6020 27412 6030
rect 27580 6020 27636 6412
rect 27356 6018 27636 6020
rect 27356 5966 27358 6018
rect 27410 5966 27636 6018
rect 27356 5964 27636 5966
rect 28028 6018 28084 6030
rect 28028 5966 28030 6018
rect 28082 5966 28084 6018
rect 27132 5954 27188 5964
rect 27020 4338 27076 4508
rect 27020 4286 27022 4338
rect 27074 4286 27076 4338
rect 27020 4274 27076 4286
rect 27356 4228 27412 5964
rect 28028 5908 28084 5966
rect 27692 5852 28084 5908
rect 27468 5796 27524 5806
rect 27692 5796 27748 5852
rect 27468 5794 27748 5796
rect 27468 5742 27470 5794
rect 27522 5742 27748 5794
rect 27468 5740 27748 5742
rect 27468 5730 27524 5740
rect 27804 5684 27860 5694
rect 28140 5684 28196 5694
rect 27804 5590 27860 5628
rect 27916 5682 28196 5684
rect 27916 5630 28142 5682
rect 28194 5630 28196 5682
rect 27916 5628 28196 5630
rect 27692 4452 27748 4462
rect 27916 4452 27972 5628
rect 28140 5618 28196 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 30268 4564 30324 4574
rect 30268 4470 30324 4508
rect 27692 4450 27972 4452
rect 27692 4398 27694 4450
rect 27746 4398 27972 4450
rect 27692 4396 27972 4398
rect 27692 4386 27748 4396
rect 27468 4228 27524 4238
rect 27356 4172 27468 4228
rect 27468 4162 27524 4172
rect 29820 4228 29876 4238
rect 29820 4134 29876 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
<< via2 >>
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5628 40514 5684 40516
rect 5628 40462 5630 40514
rect 5630 40462 5682 40514
rect 5682 40462 5684 40514
rect 5628 40460 5684 40462
rect 4956 40402 5012 40404
rect 4956 40350 4958 40402
rect 4958 40350 5010 40402
rect 5010 40350 5012 40402
rect 4956 40348 5012 40350
rect 5740 40348 5796 40404
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4732 39730 4788 39732
rect 4732 39678 4734 39730
rect 4734 39678 4786 39730
rect 4786 39678 4788 39730
rect 4732 39676 4788 39678
rect 1820 38108 1876 38164
rect 2268 38108 2324 38164
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 2940 37938 2996 37940
rect 2940 37886 2942 37938
rect 2942 37886 2994 37938
rect 2994 37886 2996 37938
rect 2940 37884 2996 37886
rect 5068 37884 5124 37940
rect 2604 37436 2660 37492
rect 4620 37490 4676 37492
rect 4620 37438 4622 37490
rect 4622 37438 4674 37490
rect 4674 37438 4676 37490
rect 4620 37436 4676 37438
rect 4396 37266 4452 37268
rect 4396 37214 4398 37266
rect 4398 37214 4450 37266
rect 4450 37214 4452 37266
rect 4396 37212 4452 37214
rect 2940 33852 2996 33908
rect 3052 32450 3108 32452
rect 3052 32398 3054 32450
rect 3054 32398 3106 32450
rect 3106 32398 3108 32450
rect 3052 32396 3108 32398
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4844 36652 4900 36708
rect 5740 38162 5796 38164
rect 5740 38110 5742 38162
rect 5742 38110 5794 38162
rect 5794 38110 5796 38162
rect 5740 38108 5796 38110
rect 5628 37266 5684 37268
rect 5628 37214 5630 37266
rect 5630 37214 5682 37266
rect 5682 37214 5684 37266
rect 5628 37212 5684 37214
rect 5292 35420 5348 35476
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 5180 35308 5236 35364
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 8764 40514 8820 40516
rect 8764 40462 8766 40514
rect 8766 40462 8818 40514
rect 8818 40462 8820 40514
rect 8764 40460 8820 40462
rect 8316 40402 8372 40404
rect 8316 40350 8318 40402
rect 8318 40350 8370 40402
rect 8370 40350 8372 40402
rect 8316 40348 8372 40350
rect 9772 40402 9828 40404
rect 9772 40350 9774 40402
rect 9774 40350 9826 40402
rect 9826 40350 9828 40402
rect 9772 40348 9828 40350
rect 12684 41916 12740 41972
rect 6188 36428 6244 36484
rect 6972 39676 7028 39732
rect 7756 39676 7812 39732
rect 8764 39730 8820 39732
rect 8764 39678 8766 39730
rect 8766 39678 8818 39730
rect 8818 39678 8820 39730
rect 8764 39676 8820 39678
rect 7420 36706 7476 36708
rect 7420 36654 7422 36706
rect 7422 36654 7474 36706
rect 7474 36654 7476 36706
rect 7420 36652 7476 36654
rect 7756 36652 7812 36708
rect 6972 36316 7028 36372
rect 6972 35420 7028 35476
rect 5068 32956 5124 33012
rect 5740 33516 5796 33572
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 2604 26908 2660 26964
rect 3724 26908 3780 26964
rect 2604 26178 2660 26180
rect 2604 26126 2606 26178
rect 2606 26126 2658 26178
rect 2658 26126 2660 26178
rect 2604 26124 2660 26126
rect 4060 26124 4116 26180
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 6636 33068 6692 33124
rect 7980 36370 8036 36372
rect 7980 36318 7982 36370
rect 7982 36318 8034 36370
rect 8034 36318 8036 36370
rect 7980 36316 8036 36318
rect 7756 34860 7812 34916
rect 8428 35532 8484 35588
rect 8540 35308 8596 35364
rect 7644 34300 7700 34356
rect 6972 33852 7028 33908
rect 7308 33292 7364 33348
rect 6748 32060 6804 32116
rect 6188 31890 6244 31892
rect 6188 31838 6190 31890
rect 6190 31838 6242 31890
rect 6242 31838 6244 31890
rect 6188 31836 6244 31838
rect 4732 29372 4788 29428
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 6972 32450 7028 32452
rect 6972 32398 6974 32450
rect 6974 32398 7026 32450
rect 7026 32398 7028 32450
rect 6972 32396 7028 32398
rect 6860 31836 6916 31892
rect 6860 30604 6916 30660
rect 6636 30210 6692 30212
rect 6636 30158 6638 30210
rect 6638 30158 6690 30210
rect 6690 30158 6692 30210
rect 6636 30156 6692 30158
rect 5964 29426 6020 29428
rect 5964 29374 5966 29426
rect 5966 29374 6018 29426
rect 6018 29374 6020 29426
rect 5964 29372 6020 29374
rect 6636 29372 6692 29428
rect 6412 29314 6468 29316
rect 6412 29262 6414 29314
rect 6414 29262 6466 29314
rect 6466 29262 6468 29314
rect 6412 29260 6468 29262
rect 4732 26178 4788 26180
rect 4732 26126 4734 26178
rect 4734 26126 4786 26178
rect 4786 26126 4788 26178
rect 4732 26124 4788 26126
rect 5964 26124 6020 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4396 25618 4452 25620
rect 4396 25566 4398 25618
rect 4398 25566 4450 25618
rect 4450 25566 4452 25618
rect 4396 25564 4452 25566
rect 5852 25618 5908 25620
rect 5852 25566 5854 25618
rect 5854 25566 5906 25618
rect 5906 25566 5908 25618
rect 5852 25564 5908 25566
rect 4060 24556 4116 24612
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 1708 22316 1764 22372
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 22482 4228 22484
rect 4172 22430 4174 22482
rect 4174 22430 4226 22482
rect 4226 22430 4228 22482
rect 4172 22428 4228 22430
rect 2604 22092 2660 22148
rect 4060 22146 4116 22148
rect 4060 22094 4062 22146
rect 4062 22094 4114 22146
rect 4114 22094 4116 22146
rect 4060 22092 4116 22094
rect 4844 22092 4900 22148
rect 5404 24668 5460 24724
rect 6076 24722 6132 24724
rect 6076 24670 6078 24722
rect 6078 24670 6130 24722
rect 6130 24670 6132 24722
rect 6076 24668 6132 24670
rect 6748 28866 6804 28868
rect 6748 28814 6750 28866
rect 6750 28814 6802 28866
rect 6802 28814 6804 28866
rect 6748 28812 6804 28814
rect 8204 33346 8260 33348
rect 8204 33294 8206 33346
rect 8206 33294 8258 33346
rect 8258 33294 8260 33346
rect 8204 33292 8260 33294
rect 7756 33122 7812 33124
rect 7756 33070 7758 33122
rect 7758 33070 7810 33122
rect 7810 33070 7812 33122
rect 7756 33068 7812 33070
rect 7756 32674 7812 32676
rect 7756 32622 7758 32674
rect 7758 32622 7810 32674
rect 7810 32622 7812 32674
rect 7756 32620 7812 32622
rect 8092 31724 8148 31780
rect 7420 30604 7476 30660
rect 7084 30098 7140 30100
rect 7084 30046 7086 30098
rect 7086 30046 7138 30098
rect 7138 30046 7140 30098
rect 7084 30044 7140 30046
rect 7420 29260 7476 29316
rect 6748 26290 6804 26292
rect 6748 26238 6750 26290
rect 6750 26238 6802 26290
rect 6802 26238 6804 26290
rect 6748 26236 6804 26238
rect 6636 26124 6692 26180
rect 6524 25340 6580 25396
rect 6300 24610 6356 24612
rect 6300 24558 6302 24610
rect 6302 24558 6354 24610
rect 6354 24558 6356 24610
rect 6300 24556 6356 24558
rect 6188 23660 6244 23716
rect 6076 23324 6132 23380
rect 5740 22482 5796 22484
rect 5740 22430 5742 22482
rect 5742 22430 5794 22482
rect 5794 22430 5796 22482
rect 5740 22428 5796 22430
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3836 20524 3892 20580
rect 1932 19964 1988 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 2604 18172 2660 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4732 17612 4788 17668
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 2716 15820 2772 15876
rect 5292 19852 5348 19908
rect 4956 18450 5012 18452
rect 4956 18398 4958 18450
rect 4958 18398 5010 18450
rect 5010 18398 5012 18450
rect 4956 18396 5012 18398
rect 5852 22146 5908 22148
rect 5852 22094 5854 22146
rect 5854 22094 5906 22146
rect 5906 22094 5908 22146
rect 5852 22092 5908 22094
rect 6748 25340 6804 25396
rect 7084 26236 7140 26292
rect 7756 28812 7812 28868
rect 7308 26178 7364 26180
rect 7308 26126 7310 26178
rect 7310 26126 7362 26178
rect 7362 26126 7364 26178
rect 7308 26124 7364 26126
rect 7308 25282 7364 25284
rect 7308 25230 7310 25282
rect 7310 25230 7362 25282
rect 7362 25230 7364 25282
rect 7308 25228 7364 25230
rect 7756 25282 7812 25284
rect 7756 25230 7758 25282
rect 7758 25230 7810 25282
rect 7810 25230 7812 25282
rect 7756 25228 7812 25230
rect 8876 35084 8932 35140
rect 9548 36652 9604 36708
rect 9884 35868 9940 35924
rect 9660 35532 9716 35588
rect 9324 34972 9380 35028
rect 8764 34524 8820 34580
rect 8540 34354 8596 34356
rect 8540 34302 8542 34354
rect 8542 34302 8594 34354
rect 8594 34302 8596 34354
rect 8540 34300 8596 34302
rect 9548 34524 9604 34580
rect 9772 34914 9828 34916
rect 9772 34862 9774 34914
rect 9774 34862 9826 34914
rect 9826 34862 9828 34914
rect 9772 34860 9828 34862
rect 10108 34802 10164 34804
rect 10108 34750 10110 34802
rect 10110 34750 10162 34802
rect 10162 34750 10164 34802
rect 10108 34748 10164 34750
rect 9996 34690 10052 34692
rect 9996 34638 9998 34690
rect 9998 34638 10050 34690
rect 10050 34638 10052 34690
rect 9996 34636 10052 34638
rect 10444 40348 10500 40404
rect 10556 40290 10612 40292
rect 10556 40238 10558 40290
rect 10558 40238 10610 40290
rect 10610 40238 10612 40290
rect 10556 40236 10612 40238
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 13468 41970 13524 41972
rect 13468 41918 13470 41970
rect 13470 41918 13522 41970
rect 13522 41918 13524 41970
rect 13468 41916 13524 41918
rect 16156 41916 16212 41972
rect 13244 41804 13300 41860
rect 14476 41858 14532 41860
rect 14476 41806 14478 41858
rect 14478 41806 14530 41858
rect 14530 41806 14532 41858
rect 14476 41804 14532 41806
rect 13356 40402 13412 40404
rect 13356 40350 13358 40402
rect 13358 40350 13410 40402
rect 13410 40350 13412 40402
rect 13356 40348 13412 40350
rect 17276 41970 17332 41972
rect 17276 41918 17278 41970
rect 17278 41918 17330 41970
rect 17330 41918 17332 41970
rect 17276 41916 17332 41918
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 16940 40402 16996 40404
rect 16940 40350 16942 40402
rect 16942 40350 16994 40402
rect 16994 40350 16996 40402
rect 16940 40348 16996 40350
rect 11116 38050 11172 38052
rect 11116 37998 11118 38050
rect 11118 37998 11170 38050
rect 11170 37998 11172 38050
rect 11116 37996 11172 37998
rect 14924 38556 14980 38612
rect 17612 40402 17668 40404
rect 17612 40350 17614 40402
rect 17614 40350 17666 40402
rect 17666 40350 17668 40402
rect 17612 40348 17668 40350
rect 20076 40348 20132 40404
rect 18956 40236 19012 40292
rect 24668 41804 24724 41860
rect 25900 41858 25956 41860
rect 25900 41806 25902 41858
rect 25902 41806 25954 41858
rect 25954 41806 25956 41858
rect 25900 41804 25956 41806
rect 20636 40460 20692 40516
rect 12908 37996 12964 38052
rect 14252 37996 14308 38052
rect 15820 37772 15876 37828
rect 10892 35868 10948 35924
rect 10332 34636 10388 34692
rect 8876 33964 8932 34020
rect 8540 33404 8596 33460
rect 9660 34018 9716 34020
rect 9660 33966 9662 34018
rect 9662 33966 9714 34018
rect 9714 33966 9716 34018
rect 9660 33964 9716 33966
rect 8540 31890 8596 31892
rect 8540 31838 8542 31890
rect 8542 31838 8594 31890
rect 8594 31838 8596 31890
rect 8540 31836 8596 31838
rect 9772 32620 9828 32676
rect 8988 31778 9044 31780
rect 8988 31726 8990 31778
rect 8990 31726 9042 31778
rect 9042 31726 9044 31778
rect 8988 31724 9044 31726
rect 9436 31554 9492 31556
rect 9436 31502 9438 31554
rect 9438 31502 9490 31554
rect 9490 31502 9492 31554
rect 9436 31500 9492 31502
rect 9212 30210 9268 30212
rect 9212 30158 9214 30210
rect 9214 30158 9266 30210
rect 9266 30158 9268 30210
rect 9212 30156 9268 30158
rect 11004 35026 11060 35028
rect 11004 34974 11006 35026
rect 11006 34974 11058 35026
rect 11058 34974 11060 35026
rect 11004 34972 11060 34974
rect 11116 34748 11172 34804
rect 10556 34188 10612 34244
rect 10220 33964 10276 34020
rect 10444 32172 10500 32228
rect 10220 30770 10276 30772
rect 10220 30718 10222 30770
rect 10222 30718 10274 30770
rect 10274 30718 10276 30770
rect 10220 30716 10276 30718
rect 10108 29484 10164 29540
rect 10668 31612 10724 31668
rect 10780 31724 10836 31780
rect 9436 29372 9492 29428
rect 10220 29426 10276 29428
rect 10220 29374 10222 29426
rect 10222 29374 10274 29426
rect 10274 29374 10276 29426
rect 10220 29372 10276 29374
rect 9772 28812 9828 28868
rect 9324 28754 9380 28756
rect 9324 28702 9326 28754
rect 9326 28702 9378 28754
rect 9378 28702 9380 28754
rect 9324 28700 9380 28702
rect 8764 28588 8820 28644
rect 10108 28642 10164 28644
rect 10108 28590 10110 28642
rect 10110 28590 10162 28642
rect 10162 28590 10164 28642
rect 10108 28588 10164 28590
rect 9996 27916 10052 27972
rect 8428 25788 8484 25844
rect 8764 25228 8820 25284
rect 8204 23378 8260 23380
rect 8204 23326 8206 23378
rect 8206 23326 8258 23378
rect 8258 23326 8260 23378
rect 8204 23324 8260 23326
rect 6188 22428 6244 22484
rect 6972 22988 7028 23044
rect 6300 22258 6356 22260
rect 6300 22206 6302 22258
rect 6302 22206 6354 22258
rect 6354 22206 6356 22258
rect 6300 22204 6356 22206
rect 5516 18508 5572 18564
rect 4956 18226 5012 18228
rect 4956 18174 4958 18226
rect 4958 18174 5010 18226
rect 5010 18174 5012 18226
rect 4956 18172 5012 18174
rect 5852 18284 5908 18340
rect 4844 15708 4900 15764
rect 4844 15372 4900 15428
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5740 17666 5796 17668
rect 5740 17614 5742 17666
rect 5742 17614 5794 17666
rect 5794 17614 5796 17666
rect 5740 17612 5796 17614
rect 5964 17724 6020 17780
rect 6524 18508 6580 18564
rect 6412 18172 6468 18228
rect 6860 19010 6916 19012
rect 6860 18958 6862 19010
rect 6862 18958 6914 19010
rect 6914 18958 6916 19010
rect 6860 18956 6916 18958
rect 7980 22988 8036 23044
rect 8428 22482 8484 22484
rect 8428 22430 8430 22482
rect 8430 22430 8482 22482
rect 8482 22430 8484 22482
rect 8428 22428 8484 22430
rect 7084 18844 7140 18900
rect 6636 18060 6692 18116
rect 6860 18450 6916 18452
rect 6860 18398 6862 18450
rect 6862 18398 6914 18450
rect 6914 18398 6916 18450
rect 6860 18396 6916 18398
rect 6748 18284 6804 18340
rect 7084 17724 7140 17780
rect 6748 17442 6804 17444
rect 6748 17390 6750 17442
rect 6750 17390 6802 17442
rect 6802 17390 6804 17442
rect 6748 17388 6804 17390
rect 7980 18226 8036 18228
rect 7980 18174 7982 18226
rect 7982 18174 8034 18226
rect 8034 18174 8036 18226
rect 7980 18172 8036 18174
rect 7756 18060 7812 18116
rect 7980 17724 8036 17780
rect 7420 17388 7476 17444
rect 7868 16098 7924 16100
rect 7868 16046 7870 16098
rect 7870 16046 7922 16098
rect 7922 16046 7924 16098
rect 7868 16044 7924 16046
rect 7756 15932 7812 15988
rect 7532 15874 7588 15876
rect 7532 15822 7534 15874
rect 7534 15822 7586 15874
rect 7586 15822 7588 15874
rect 7532 15820 7588 15822
rect 6860 15372 6916 15428
rect 7308 15314 7364 15316
rect 7308 15262 7310 15314
rect 7310 15262 7362 15314
rect 7362 15262 7364 15314
rect 7308 15260 7364 15262
rect 6860 14364 6916 14420
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2604 12290 2660 12292
rect 2604 12238 2606 12290
rect 2606 12238 2658 12290
rect 2658 12238 2660 12290
rect 2604 12236 2660 12238
rect 4732 12124 4788 12180
rect 6076 13020 6132 13076
rect 6300 12796 6356 12852
rect 6076 12178 6132 12180
rect 6076 12126 6078 12178
rect 6078 12126 6130 12178
rect 6130 12126 6132 12178
rect 6076 12124 6132 12126
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4508 9548 4564 9604
rect 3836 9042 3892 9044
rect 3836 8990 3838 9042
rect 3838 8990 3890 9042
rect 3890 8990 3892 9042
rect 3836 8988 3892 8990
rect 7756 14364 7812 14420
rect 7644 13020 7700 13076
rect 7756 12796 7812 12852
rect 7980 15260 8036 15316
rect 7644 12290 7700 12292
rect 7644 12238 7646 12290
rect 7646 12238 7698 12290
rect 7698 12238 7700 12290
rect 7644 12236 7700 12238
rect 6524 11116 6580 11172
rect 7196 11282 7252 11284
rect 7196 11230 7198 11282
rect 7198 11230 7250 11282
rect 7250 11230 7252 11282
rect 7196 11228 7252 11230
rect 7532 11170 7588 11172
rect 7532 11118 7534 11170
rect 7534 11118 7586 11170
rect 7586 11118 7588 11170
rect 7532 11116 7588 11118
rect 7644 10892 7700 10948
rect 7196 10610 7252 10612
rect 7196 10558 7198 10610
rect 7198 10558 7250 10610
rect 7250 10558 7252 10610
rect 7196 10556 7252 10558
rect 7868 12178 7924 12180
rect 7868 12126 7870 12178
rect 7870 12126 7922 12178
rect 7922 12126 7924 12178
rect 7868 12124 7924 12126
rect 7868 11116 7924 11172
rect 6748 9772 6804 9828
rect 6636 9602 6692 9604
rect 6636 9550 6638 9602
rect 6638 9550 6690 9602
rect 6690 9550 6692 9602
rect 6636 9548 6692 9550
rect 5180 8988 5236 9044
rect 7308 9826 7364 9828
rect 7308 9774 7310 9826
rect 7310 9774 7362 9826
rect 7362 9774 7364 9826
rect 7308 9772 7364 9774
rect 8204 16156 8260 16212
rect 8540 15986 8596 15988
rect 8540 15934 8542 15986
rect 8542 15934 8594 15986
rect 8594 15934 8596 15986
rect 8540 15932 8596 15934
rect 8652 15372 8708 15428
rect 9100 23938 9156 23940
rect 9100 23886 9102 23938
rect 9102 23886 9154 23938
rect 9154 23886 9156 23938
rect 9100 23884 9156 23886
rect 8876 23714 8932 23716
rect 8876 23662 8878 23714
rect 8878 23662 8930 23714
rect 8930 23662 8932 23714
rect 8876 23660 8932 23662
rect 9436 23996 9492 24052
rect 9212 23100 9268 23156
rect 9660 23660 9716 23716
rect 10780 28642 10836 28644
rect 10780 28590 10782 28642
rect 10782 28590 10834 28642
rect 10834 28590 10836 28642
rect 10780 28588 10836 28590
rect 9884 23100 9940 23156
rect 11676 34748 11732 34804
rect 11340 33964 11396 34020
rect 12012 34242 12068 34244
rect 12012 34190 12014 34242
rect 12014 34190 12066 34242
rect 12066 34190 12068 34242
rect 12012 34188 12068 34190
rect 12796 33964 12852 34020
rect 12124 33628 12180 33684
rect 12012 33516 12068 33572
rect 11900 32172 11956 32228
rect 11116 31724 11172 31780
rect 11452 31612 11508 31668
rect 11116 31388 11172 31444
rect 11116 30716 11172 30772
rect 12460 33628 12516 33684
rect 13804 33292 13860 33348
rect 12124 32786 12180 32788
rect 12124 32734 12126 32786
rect 12126 32734 12178 32786
rect 12178 32734 12180 32786
rect 12124 32732 12180 32734
rect 11228 30210 11284 30212
rect 11228 30158 11230 30210
rect 11230 30158 11282 30210
rect 11282 30158 11284 30210
rect 11228 30156 11284 30158
rect 11564 30098 11620 30100
rect 11564 30046 11566 30098
rect 11566 30046 11618 30098
rect 11618 30046 11620 30098
rect 11564 30044 11620 30046
rect 11676 29986 11732 29988
rect 11676 29934 11678 29986
rect 11678 29934 11730 29986
rect 11730 29934 11732 29986
rect 11676 29932 11732 29934
rect 11116 29372 11172 29428
rect 11676 29426 11732 29428
rect 11676 29374 11678 29426
rect 11678 29374 11730 29426
rect 11730 29374 11732 29426
rect 11676 29372 11732 29374
rect 11004 26514 11060 26516
rect 11004 26462 11006 26514
rect 11006 26462 11058 26514
rect 11058 26462 11060 26514
rect 11004 26460 11060 26462
rect 10892 23996 10948 24052
rect 10780 23938 10836 23940
rect 10780 23886 10782 23938
rect 10782 23886 10834 23938
rect 10834 23886 10836 23938
rect 10780 23884 10836 23886
rect 10220 22204 10276 22260
rect 9884 22092 9940 22148
rect 11228 25900 11284 25956
rect 11228 25228 11284 25284
rect 11228 23996 11284 24052
rect 11788 26514 11844 26516
rect 11788 26462 11790 26514
rect 11790 26462 11842 26514
rect 11842 26462 11844 26514
rect 11788 26460 11844 26462
rect 11452 25282 11508 25284
rect 11452 25230 11454 25282
rect 11454 25230 11506 25282
rect 11506 25230 11508 25282
rect 11452 25228 11508 25230
rect 11452 23772 11508 23828
rect 11228 23378 11284 23380
rect 11228 23326 11230 23378
rect 11230 23326 11282 23378
rect 11282 23326 11284 23378
rect 11228 23324 11284 23326
rect 11452 23378 11508 23380
rect 11452 23326 11454 23378
rect 11454 23326 11506 23378
rect 11506 23326 11508 23378
rect 11452 23324 11508 23326
rect 11228 23100 11284 23156
rect 9100 20748 9156 20804
rect 10668 20578 10724 20580
rect 10668 20526 10670 20578
rect 10670 20526 10722 20578
rect 10722 20526 10724 20578
rect 10668 20524 10724 20526
rect 11452 21532 11508 21588
rect 10892 20076 10948 20132
rect 9884 19852 9940 19908
rect 9548 18396 9604 18452
rect 9884 18450 9940 18452
rect 9884 18398 9886 18450
rect 9886 18398 9938 18450
rect 9938 18398 9940 18450
rect 9884 18396 9940 18398
rect 11228 18396 11284 18452
rect 12124 30098 12180 30100
rect 12124 30046 12126 30098
rect 12126 30046 12178 30098
rect 12178 30046 12180 30098
rect 12124 30044 12180 30046
rect 12124 28812 12180 28868
rect 12460 33180 12516 33236
rect 13020 33068 13076 33124
rect 13020 32786 13076 32788
rect 13020 32734 13022 32786
rect 13022 32734 13074 32786
rect 13074 32734 13076 32786
rect 13020 32732 13076 32734
rect 15148 36316 15204 36372
rect 15036 33234 15092 33236
rect 15036 33182 15038 33234
rect 15038 33182 15090 33234
rect 15090 33182 15092 33234
rect 15036 33180 15092 33182
rect 14700 33122 14756 33124
rect 14700 33070 14702 33122
rect 14702 33070 14754 33122
rect 14754 33070 14756 33122
rect 14700 33068 14756 33070
rect 13580 32172 13636 32228
rect 16604 38668 16660 38724
rect 18508 39506 18564 39508
rect 18508 39454 18510 39506
rect 18510 39454 18562 39506
rect 18562 39454 18564 39506
rect 18508 39452 18564 39454
rect 19068 39506 19124 39508
rect 19068 39454 19070 39506
rect 19070 39454 19122 39506
rect 19122 39454 19124 39506
rect 19068 39452 19124 39454
rect 19852 39506 19908 39508
rect 19852 39454 19854 39506
rect 19854 39454 19906 39506
rect 19906 39454 19908 39506
rect 19852 39452 19908 39454
rect 20188 39452 20244 39508
rect 18284 39394 18340 39396
rect 18284 39342 18286 39394
rect 18286 39342 18338 39394
rect 18338 39342 18340 39394
rect 18284 39340 18340 39342
rect 18844 39394 18900 39396
rect 18844 39342 18846 39394
rect 18846 39342 18898 39394
rect 18898 39342 18900 39394
rect 18844 39340 18900 39342
rect 20076 39394 20132 39396
rect 20076 39342 20078 39394
rect 20078 39342 20130 39394
rect 20130 39342 20132 39394
rect 20076 39340 20132 39342
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 17948 38668 18004 38724
rect 16380 37772 16436 37828
rect 20524 38946 20580 38948
rect 20524 38894 20526 38946
rect 20526 38894 20578 38946
rect 20578 38894 20580 38946
rect 20524 38892 20580 38894
rect 20188 38834 20244 38836
rect 20188 38782 20190 38834
rect 20190 38782 20242 38834
rect 20242 38782 20244 38834
rect 20188 38780 20244 38782
rect 20076 37938 20132 37940
rect 20076 37886 20078 37938
rect 20078 37886 20130 37938
rect 20130 37886 20132 37938
rect 20076 37884 20132 37886
rect 19180 37826 19236 37828
rect 19180 37774 19182 37826
rect 19182 37774 19234 37826
rect 19234 37774 19236 37826
rect 19180 37772 19236 37774
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 23660 40402 23716 40404
rect 23660 40350 23662 40402
rect 23662 40350 23714 40402
rect 23714 40350 23716 40402
rect 23660 40348 23716 40350
rect 23772 39452 23828 39508
rect 23548 38610 23604 38612
rect 23548 38558 23550 38610
rect 23550 38558 23602 38610
rect 23602 38558 23604 38610
rect 23548 38556 23604 38558
rect 20412 38274 20468 38276
rect 20412 38222 20414 38274
rect 20414 38222 20466 38274
rect 20466 38222 20468 38274
rect 20412 38220 20468 38222
rect 23772 38780 23828 38836
rect 20524 37938 20580 37940
rect 20524 37886 20526 37938
rect 20526 37886 20578 37938
rect 20578 37886 20580 37938
rect 20524 37884 20580 37886
rect 21420 37884 21476 37940
rect 19740 36482 19796 36484
rect 19740 36430 19742 36482
rect 19742 36430 19794 36482
rect 19794 36430 19796 36482
rect 19740 36428 19796 36430
rect 20188 36482 20244 36484
rect 20188 36430 20190 36482
rect 20190 36430 20242 36482
rect 20242 36430 20244 36482
rect 20188 36428 20244 36430
rect 18732 36316 18788 36372
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20524 36316 20580 36372
rect 20412 36258 20468 36260
rect 20412 36206 20414 36258
rect 20414 36206 20466 36258
rect 20466 36206 20468 36258
rect 20412 36204 20468 36206
rect 15820 34636 15876 34692
rect 20188 34914 20244 34916
rect 20188 34862 20190 34914
rect 20190 34862 20242 34914
rect 20242 34862 20244 34914
rect 20188 34860 20244 34862
rect 20412 35084 20468 35140
rect 16604 34636 16660 34692
rect 17164 34690 17220 34692
rect 17164 34638 17166 34690
rect 17166 34638 17218 34690
rect 17218 34638 17220 34690
rect 17164 34636 17220 34638
rect 18284 34636 18340 34692
rect 15484 33292 15540 33348
rect 15260 33122 15316 33124
rect 15260 33070 15262 33122
rect 15262 33070 15314 33122
rect 15314 33070 15316 33122
rect 15260 33068 15316 33070
rect 15036 32284 15092 32340
rect 14588 32060 14644 32116
rect 12572 31388 12628 31444
rect 15036 31164 15092 31220
rect 14588 30210 14644 30212
rect 14588 30158 14590 30210
rect 14590 30158 14642 30210
rect 14642 30158 14644 30210
rect 14588 30156 14644 30158
rect 14700 30044 14756 30100
rect 13468 28700 13524 28756
rect 12908 28028 12964 28084
rect 12908 26908 12964 26964
rect 13244 27746 13300 27748
rect 13244 27694 13246 27746
rect 13246 27694 13298 27746
rect 13298 27694 13300 27746
rect 13244 27692 13300 27694
rect 12348 26514 12404 26516
rect 12348 26462 12350 26514
rect 12350 26462 12402 26514
rect 12402 26462 12404 26514
rect 12348 26460 12404 26462
rect 12684 26236 12740 26292
rect 12012 25900 12068 25956
rect 13132 25900 13188 25956
rect 12012 23378 12068 23380
rect 12012 23326 12014 23378
rect 12014 23326 12066 23378
rect 12066 23326 12068 23378
rect 12012 23324 12068 23326
rect 12348 23378 12404 23380
rect 12348 23326 12350 23378
rect 12350 23326 12402 23378
rect 12402 23326 12404 23378
rect 12348 23324 12404 23326
rect 12684 23324 12740 23380
rect 11900 18450 11956 18452
rect 11900 18398 11902 18450
rect 11902 18398 11954 18450
rect 11954 18398 11956 18450
rect 11900 18396 11956 18398
rect 9100 16210 9156 16212
rect 9100 16158 9102 16210
rect 9102 16158 9154 16210
rect 9154 16158 9156 16210
rect 9100 16156 9156 16158
rect 9660 16044 9716 16100
rect 8876 15538 8932 15540
rect 8876 15486 8878 15538
rect 8878 15486 8930 15538
rect 8930 15486 8932 15538
rect 8876 15484 8932 15486
rect 11676 16882 11732 16884
rect 11676 16830 11678 16882
rect 11678 16830 11730 16882
rect 11730 16830 11732 16882
rect 11676 16828 11732 16830
rect 12348 18450 12404 18452
rect 12348 18398 12350 18450
rect 12350 18398 12402 18450
rect 12402 18398 12404 18450
rect 12348 18396 12404 18398
rect 13020 16098 13076 16100
rect 13020 16046 13022 16098
rect 13022 16046 13074 16098
rect 13074 16046 13076 16098
rect 13020 16044 13076 16046
rect 9884 15426 9940 15428
rect 9884 15374 9886 15426
rect 9886 15374 9938 15426
rect 9938 15374 9940 15426
rect 9884 15372 9940 15374
rect 9548 15314 9604 15316
rect 9548 15262 9550 15314
rect 9550 15262 9602 15314
rect 9602 15262 9604 15314
rect 9548 15260 9604 15262
rect 8764 15148 8820 15204
rect 9436 15148 9492 15204
rect 8764 12796 8820 12852
rect 8540 12738 8596 12740
rect 8540 12686 8542 12738
rect 8542 12686 8594 12738
rect 8594 12686 8596 12738
rect 8540 12684 8596 12686
rect 8428 12348 8484 12404
rect 8652 12178 8708 12180
rect 8652 12126 8654 12178
rect 8654 12126 8706 12178
rect 8706 12126 8708 12178
rect 8652 12124 8708 12126
rect 9100 12012 9156 12068
rect 8876 11452 8932 11508
rect 8316 11170 8372 11172
rect 8316 11118 8318 11170
rect 8318 11118 8370 11170
rect 8370 11118 8372 11170
rect 8316 11116 8372 11118
rect 8092 10892 8148 10948
rect 8876 11228 8932 11284
rect 10220 15260 10276 15316
rect 12460 15708 12516 15764
rect 12460 15260 12516 15316
rect 9660 14418 9716 14420
rect 9660 14366 9662 14418
rect 9662 14366 9714 14418
rect 9714 14366 9716 14418
rect 9660 14364 9716 14366
rect 9996 14252 10052 14308
rect 9660 12402 9716 12404
rect 9660 12350 9662 12402
rect 9662 12350 9714 12402
rect 9714 12350 9716 12402
rect 9660 12348 9716 12350
rect 9324 11506 9380 11508
rect 9324 11454 9326 11506
rect 9326 11454 9378 11506
rect 9378 11454 9380 11506
rect 9324 11452 9380 11454
rect 11564 12684 11620 12740
rect 12236 12290 12292 12292
rect 12236 12238 12238 12290
rect 12238 12238 12290 12290
rect 12290 12238 12292 12290
rect 12236 12236 12292 12238
rect 10220 11116 10276 11172
rect 11340 11340 11396 11396
rect 8092 10610 8148 10612
rect 8092 10558 8094 10610
rect 8094 10558 8146 10610
rect 8146 10558 8148 10610
rect 8092 10556 8148 10558
rect 11228 10610 11284 10612
rect 11228 10558 11230 10610
rect 11230 10558 11282 10610
rect 11282 10558 11284 10610
rect 11228 10556 11284 10558
rect 10780 9996 10836 10052
rect 7980 9772 8036 9828
rect 8092 9884 8148 9940
rect 11788 11228 11844 11284
rect 12236 11394 12292 11396
rect 12236 11342 12238 11394
rect 12238 11342 12290 11394
rect 12290 11342 12292 11394
rect 12236 11340 12292 11342
rect 11676 10556 11732 10612
rect 12348 11282 12404 11284
rect 12348 11230 12350 11282
rect 12350 11230 12402 11282
rect 12402 11230 12404 11282
rect 12348 11228 12404 11230
rect 12236 10556 12292 10612
rect 13692 27970 13748 27972
rect 13692 27918 13694 27970
rect 13694 27918 13746 27970
rect 13746 27918 13748 27970
rect 13692 27916 13748 27918
rect 14588 29538 14644 29540
rect 14588 29486 14590 29538
rect 14590 29486 14642 29538
rect 14642 29486 14644 29538
rect 14588 29484 14644 29486
rect 14364 28700 14420 28756
rect 14028 27692 14084 27748
rect 14924 28028 14980 28084
rect 14924 27858 14980 27860
rect 14924 27806 14926 27858
rect 14926 27806 14978 27858
rect 14978 27806 14980 27858
rect 14924 27804 14980 27806
rect 15484 32786 15540 32788
rect 15484 32734 15486 32786
rect 15486 32734 15538 32786
rect 15538 32734 15540 32786
rect 15484 32732 15540 32734
rect 15932 33964 15988 34020
rect 16380 34018 16436 34020
rect 16380 33966 16382 34018
rect 16382 33966 16434 34018
rect 16434 33966 16436 34018
rect 16380 33964 16436 33966
rect 15820 33292 15876 33348
rect 17276 33180 17332 33236
rect 17052 33122 17108 33124
rect 17052 33070 17054 33122
rect 17054 33070 17106 33122
rect 17106 33070 17108 33122
rect 17052 33068 17108 33070
rect 16380 32732 16436 32788
rect 15820 32674 15876 32676
rect 15820 32622 15822 32674
rect 15822 32622 15874 32674
rect 15874 32622 15876 32674
rect 15820 32620 15876 32622
rect 16044 32562 16100 32564
rect 16044 32510 16046 32562
rect 16046 32510 16098 32562
rect 16098 32510 16100 32562
rect 16044 32508 16100 32510
rect 16716 32620 16772 32676
rect 16268 32338 16324 32340
rect 16268 32286 16270 32338
rect 16270 32286 16322 32338
rect 16322 32286 16324 32338
rect 16268 32284 16324 32286
rect 15484 31724 15540 31780
rect 15820 30828 15876 30884
rect 16044 30210 16100 30212
rect 16044 30158 16046 30210
rect 16046 30158 16098 30210
rect 16098 30158 16100 30210
rect 16044 30156 16100 30158
rect 15596 30098 15652 30100
rect 15596 30046 15598 30098
rect 15598 30046 15650 30098
rect 15650 30046 15652 30098
rect 15596 30044 15652 30046
rect 15148 29484 15204 29540
rect 15260 27804 15316 27860
rect 16380 30882 16436 30884
rect 16380 30830 16382 30882
rect 16382 30830 16434 30882
rect 16434 30830 16436 30882
rect 16380 30828 16436 30830
rect 16268 29708 16324 29764
rect 16156 28700 16212 28756
rect 16492 29932 16548 29988
rect 15484 28642 15540 28644
rect 15484 28590 15486 28642
rect 15486 28590 15538 28642
rect 15538 28590 15540 28642
rect 15484 28588 15540 28590
rect 15372 27916 15428 27972
rect 14140 26850 14196 26852
rect 14140 26798 14142 26850
rect 14142 26798 14194 26850
rect 14194 26798 14196 26850
rect 14140 26796 14196 26798
rect 15372 26796 15428 26852
rect 13692 26684 13748 26740
rect 13580 24332 13636 24388
rect 15820 28530 15876 28532
rect 15820 28478 15822 28530
rect 15822 28478 15874 28530
rect 15874 28478 15876 28530
rect 15820 28476 15876 28478
rect 16156 27916 16212 27972
rect 15596 26572 15652 26628
rect 14252 24332 14308 24388
rect 13356 23324 13412 23380
rect 13244 15484 13300 15540
rect 15708 23884 15764 23940
rect 13692 22988 13748 23044
rect 13692 21868 13748 21924
rect 14588 21868 14644 21924
rect 13468 18396 13524 18452
rect 13132 15260 13188 15316
rect 12796 14252 12852 14308
rect 13468 13356 13524 13412
rect 12796 12290 12852 12292
rect 12796 12238 12798 12290
rect 12798 12238 12850 12290
rect 12850 12238 12852 12290
rect 12796 12236 12852 12238
rect 13468 12236 13524 12292
rect 13804 20524 13860 20580
rect 13692 20018 13748 20020
rect 13692 19966 13694 20018
rect 13694 19966 13746 20018
rect 13746 19966 13748 20018
rect 13692 19964 13748 19966
rect 13580 19852 13636 19908
rect 15820 27804 15876 27860
rect 15260 21586 15316 21588
rect 15260 21534 15262 21586
rect 15262 21534 15314 21586
rect 15314 21534 15316 21586
rect 15260 21532 15316 21534
rect 14700 21420 14756 21476
rect 15596 21474 15652 21476
rect 15596 21422 15598 21474
rect 15598 21422 15650 21474
rect 15650 21422 15652 21474
rect 15596 21420 15652 21422
rect 14476 20578 14532 20580
rect 14476 20526 14478 20578
rect 14478 20526 14530 20578
rect 14530 20526 14532 20578
rect 14476 20524 14532 20526
rect 13468 11228 13524 11284
rect 12684 10668 12740 10724
rect 11564 9996 11620 10052
rect 12124 9996 12180 10052
rect 12460 9996 12516 10052
rect 7084 9042 7140 9044
rect 7084 8990 7086 9042
rect 7086 8990 7138 9042
rect 7138 8990 7140 9042
rect 7084 8988 7140 8990
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 10892 8316 10948 8372
rect 11564 8370 11620 8372
rect 11564 8318 11566 8370
rect 11566 8318 11618 8370
rect 11618 8318 11620 8370
rect 11564 8316 11620 8318
rect 12908 9996 12964 10052
rect 12796 9548 12852 9604
rect 12572 8316 12628 8372
rect 12572 7980 12628 8036
rect 9996 6690 10052 6692
rect 9996 6638 9998 6690
rect 9998 6638 10050 6690
rect 10050 6638 10052 6690
rect 9996 6636 10052 6638
rect 12124 6636 12180 6692
rect 14140 18508 14196 18564
rect 14028 15426 14084 15428
rect 14028 15374 14030 15426
rect 14030 15374 14082 15426
rect 14082 15374 14084 15426
rect 14028 15372 14084 15374
rect 16044 27804 16100 27860
rect 16380 27804 16436 27860
rect 16268 26460 16324 26516
rect 17612 33068 17668 33124
rect 17836 32508 17892 32564
rect 16940 30940 16996 30996
rect 16716 29708 16772 29764
rect 16716 28812 16772 28868
rect 16828 26402 16884 26404
rect 16828 26350 16830 26402
rect 16830 26350 16882 26402
rect 16882 26350 16884 26402
rect 16828 26348 16884 26350
rect 16604 26290 16660 26292
rect 16604 26238 16606 26290
rect 16606 26238 16658 26290
rect 16658 26238 16660 26290
rect 16604 26236 16660 26238
rect 16044 23324 16100 23380
rect 16716 25340 16772 25396
rect 16268 24050 16324 24052
rect 16268 23998 16270 24050
rect 16270 23998 16322 24050
rect 16322 23998 16324 24050
rect 16268 23996 16324 23998
rect 16492 23884 16548 23940
rect 16044 20188 16100 20244
rect 14812 17388 14868 17444
rect 15708 17388 15764 17444
rect 15484 16828 15540 16884
rect 15932 16604 15988 16660
rect 14364 15820 14420 15876
rect 15260 14588 15316 14644
rect 16044 15820 16100 15876
rect 13804 14306 13860 14308
rect 13804 14254 13806 14306
rect 13806 14254 13858 14306
rect 13858 14254 13860 14306
rect 13804 14252 13860 14254
rect 13804 11900 13860 11956
rect 13692 11282 13748 11284
rect 13692 11230 13694 11282
rect 13694 11230 13746 11282
rect 13746 11230 13748 11282
rect 13692 11228 13748 11230
rect 14252 13356 14308 13412
rect 14812 12066 14868 12068
rect 14812 12014 14814 12066
rect 14814 12014 14866 12066
rect 14866 12014 14868 12066
rect 14812 12012 14868 12014
rect 15036 11954 15092 11956
rect 15036 11902 15038 11954
rect 15038 11902 15090 11954
rect 15090 11902 15092 11954
rect 15036 11900 15092 11902
rect 15260 11676 15316 11732
rect 15708 11340 15764 11396
rect 13804 10610 13860 10612
rect 13804 10558 13806 10610
rect 13806 10558 13858 10610
rect 13858 10558 13860 10610
rect 13804 10556 13860 10558
rect 16044 11676 16100 11732
rect 14028 10780 14084 10836
rect 15260 10610 15316 10612
rect 15260 10558 15262 10610
rect 15262 10558 15314 10610
rect 15314 10558 15316 10610
rect 15260 10556 15316 10558
rect 15932 10722 15988 10724
rect 15932 10670 15934 10722
rect 15934 10670 15986 10722
rect 15986 10670 15988 10722
rect 15932 10668 15988 10670
rect 14364 9996 14420 10052
rect 13692 9548 13748 9604
rect 15820 9996 15876 10052
rect 17948 30268 18004 30324
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 18508 33964 18564 34020
rect 18284 28700 18340 28756
rect 17836 27020 17892 27076
rect 17276 26572 17332 26628
rect 17388 26514 17444 26516
rect 17388 26462 17390 26514
rect 17390 26462 17442 26514
rect 17442 26462 17444 26514
rect 17388 26460 17444 26462
rect 17948 26402 18004 26404
rect 17948 26350 17950 26402
rect 17950 26350 18002 26402
rect 18002 26350 18004 26402
rect 17948 26348 18004 26350
rect 17276 25394 17332 25396
rect 17276 25342 17278 25394
rect 17278 25342 17330 25394
rect 17330 25342 17332 25394
rect 17276 25340 17332 25342
rect 18060 25340 18116 25396
rect 17276 23938 17332 23940
rect 17276 23886 17278 23938
rect 17278 23886 17330 23938
rect 17330 23886 17332 23938
rect 17276 23884 17332 23886
rect 16940 23436 16996 23492
rect 17388 23378 17444 23380
rect 17388 23326 17390 23378
rect 17390 23326 17442 23378
rect 17442 23326 17444 23378
rect 17388 23324 17444 23326
rect 17500 23266 17556 23268
rect 17500 23214 17502 23266
rect 17502 23214 17554 23266
rect 17554 23214 17556 23266
rect 17500 23212 17556 23214
rect 17724 23436 17780 23492
rect 17724 23154 17780 23156
rect 17724 23102 17726 23154
rect 17726 23102 17778 23154
rect 17778 23102 17780 23154
rect 17724 23100 17780 23102
rect 17500 21756 17556 21812
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20412 32844 20468 32900
rect 20300 32786 20356 32788
rect 20300 32734 20302 32786
rect 20302 32734 20354 32786
rect 20354 32734 20356 32786
rect 20300 32732 20356 32734
rect 19404 31612 19460 31668
rect 19068 31500 19124 31556
rect 18956 30604 19012 30660
rect 18508 27916 18564 27972
rect 18620 30268 18676 30324
rect 18844 30268 18900 30324
rect 19292 30994 19348 30996
rect 19292 30942 19294 30994
rect 19294 30942 19346 30994
rect 19346 30942 19348 30994
rect 19292 30940 19348 30942
rect 19516 32172 19572 32228
rect 19628 31836 19684 31892
rect 20076 31890 20132 31892
rect 20076 31838 20078 31890
rect 20078 31838 20130 31890
rect 20130 31838 20132 31890
rect 20076 31836 20132 31838
rect 21644 36482 21700 36484
rect 21644 36430 21646 36482
rect 21646 36430 21698 36482
rect 21698 36430 21700 36482
rect 21644 36428 21700 36430
rect 21868 36204 21924 36260
rect 25788 40348 25844 40404
rect 24220 40290 24276 40292
rect 24220 40238 24222 40290
rect 24222 40238 24274 40290
rect 24274 40238 24276 40290
rect 24220 40236 24276 40238
rect 24780 39058 24836 39060
rect 24780 39006 24782 39058
rect 24782 39006 24834 39058
rect 24834 39006 24836 39058
rect 24780 39004 24836 39006
rect 25676 40236 25732 40292
rect 24220 38220 24276 38276
rect 24556 38946 24612 38948
rect 24556 38894 24558 38946
rect 24558 38894 24610 38946
rect 24610 38894 24612 38946
rect 24556 38892 24612 38894
rect 25452 38220 25508 38276
rect 26460 39618 26516 39620
rect 26460 39566 26462 39618
rect 26462 39566 26514 39618
rect 26514 39566 26516 39618
rect 26460 39564 26516 39566
rect 26908 39618 26964 39620
rect 26908 39566 26910 39618
rect 26910 39566 26962 39618
rect 26962 39566 26964 39618
rect 26908 39564 26964 39566
rect 28476 40402 28532 40404
rect 28476 40350 28478 40402
rect 28478 40350 28530 40402
rect 28530 40350 28532 40402
rect 28476 40348 28532 40350
rect 31164 40402 31220 40404
rect 31164 40350 31166 40402
rect 31166 40350 31218 40402
rect 31218 40350 31220 40402
rect 31164 40348 31220 40350
rect 27804 39564 27860 39620
rect 29820 39618 29876 39620
rect 29820 39566 29822 39618
rect 29822 39566 29874 39618
rect 29874 39566 29876 39618
rect 29820 39564 29876 39566
rect 26460 39340 26516 39396
rect 27132 39340 27188 39396
rect 26124 38834 26180 38836
rect 26124 38782 26126 38834
rect 26126 38782 26178 38834
rect 26178 38782 26180 38834
rect 26124 38780 26180 38782
rect 23884 37436 23940 37492
rect 25228 37490 25284 37492
rect 25228 37438 25230 37490
rect 25230 37438 25282 37490
rect 25282 37438 25284 37490
rect 25228 37436 25284 37438
rect 23436 36428 23492 36484
rect 21868 35308 21924 35364
rect 22988 35308 23044 35364
rect 20636 34636 20692 34692
rect 20636 34130 20692 34132
rect 20636 34078 20638 34130
rect 20638 34078 20690 34130
rect 20690 34078 20692 34130
rect 20636 34076 20692 34078
rect 21084 33516 21140 33572
rect 21084 32732 21140 32788
rect 22764 34188 22820 34244
rect 22204 33516 22260 33572
rect 22204 32562 22260 32564
rect 22204 32510 22206 32562
rect 22206 32510 22258 32562
rect 22258 32510 22260 32562
rect 22204 32508 22260 32510
rect 22652 32450 22708 32452
rect 22652 32398 22654 32450
rect 22654 32398 22706 32450
rect 22706 32398 22708 32450
rect 22652 32396 22708 32398
rect 19852 31778 19908 31780
rect 19852 31726 19854 31778
rect 19854 31726 19906 31778
rect 19906 31726 19908 31778
rect 19852 31724 19908 31726
rect 20412 31666 20468 31668
rect 20412 31614 20414 31666
rect 20414 31614 20466 31666
rect 20466 31614 20468 31666
rect 20412 31612 20468 31614
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19628 31164 19684 31220
rect 19516 30268 19572 30324
rect 20636 30882 20692 30884
rect 20636 30830 20638 30882
rect 20638 30830 20690 30882
rect 20690 30830 20692 30882
rect 20636 30828 20692 30830
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20412 29260 20468 29316
rect 19404 28754 19460 28756
rect 19404 28702 19406 28754
rect 19406 28702 19458 28754
rect 19458 28702 19460 28754
rect 19404 28700 19460 28702
rect 19292 27916 19348 27972
rect 18732 26402 18788 26404
rect 18732 26350 18734 26402
rect 18734 26350 18786 26402
rect 18786 26350 18788 26402
rect 18732 26348 18788 26350
rect 18956 27746 19012 27748
rect 18956 27694 18958 27746
rect 18958 27694 19010 27746
rect 19010 27694 19012 27746
rect 18956 27692 19012 27694
rect 18956 26290 19012 26292
rect 18956 26238 18958 26290
rect 18958 26238 19010 26290
rect 19010 26238 19012 26290
rect 18956 26236 19012 26238
rect 21308 28476 21364 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20524 27746 20580 27748
rect 20524 27694 20526 27746
rect 20526 27694 20578 27746
rect 20578 27694 20580 27746
rect 20524 27692 20580 27694
rect 19740 27186 19796 27188
rect 19740 27134 19742 27186
rect 19742 27134 19794 27186
rect 19794 27134 19796 27186
rect 19740 27132 19796 27134
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19628 26402 19684 26404
rect 19628 26350 19630 26402
rect 19630 26350 19682 26402
rect 19682 26350 19684 26402
rect 19628 26348 19684 26350
rect 18396 24332 18452 24388
rect 18396 23436 18452 23492
rect 18396 23100 18452 23156
rect 19180 23772 19236 23828
rect 19180 23154 19236 23156
rect 19180 23102 19182 23154
rect 19182 23102 19234 23154
rect 19234 23102 19236 23154
rect 19180 23100 19236 23102
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 21756 27074 21812 27076
rect 21756 27022 21758 27074
rect 21758 27022 21810 27074
rect 21810 27022 21812 27074
rect 21756 27020 21812 27022
rect 22652 27020 22708 27076
rect 23324 34242 23380 34244
rect 23324 34190 23326 34242
rect 23326 34190 23378 34242
rect 23378 34190 23380 34242
rect 23324 34188 23380 34190
rect 24556 36988 24612 37044
rect 23660 36316 23716 36372
rect 25564 37042 25620 37044
rect 25564 36990 25566 37042
rect 25566 36990 25618 37042
rect 25618 36990 25620 37042
rect 25564 36988 25620 36990
rect 25788 36876 25844 36932
rect 24444 34914 24500 34916
rect 24444 34862 24446 34914
rect 24446 34862 24498 34914
rect 24498 34862 24500 34914
rect 24444 34860 24500 34862
rect 23548 34076 23604 34132
rect 24220 34690 24276 34692
rect 24220 34638 24222 34690
rect 24222 34638 24274 34690
rect 24274 34638 24276 34690
rect 24220 34636 24276 34638
rect 23884 34018 23940 34020
rect 23884 33966 23886 34018
rect 23886 33966 23938 34018
rect 23938 33966 23940 34018
rect 23884 33964 23940 33966
rect 23660 33906 23716 33908
rect 23660 33854 23662 33906
rect 23662 33854 23714 33906
rect 23714 33854 23716 33906
rect 23660 33852 23716 33854
rect 23100 32844 23156 32900
rect 22988 26796 23044 26852
rect 23772 26178 23828 26180
rect 23772 26126 23774 26178
rect 23774 26126 23826 26178
rect 23826 26126 23828 26178
rect 23772 26124 23828 26126
rect 23772 25788 23828 25844
rect 20412 23826 20468 23828
rect 20412 23774 20414 23826
rect 20414 23774 20466 23826
rect 20466 23774 20468 23826
rect 20412 23772 20468 23774
rect 21756 23772 21812 23828
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19740 23100 19796 23156
rect 23548 23826 23604 23828
rect 23548 23774 23550 23826
rect 23550 23774 23602 23826
rect 23602 23774 23604 23826
rect 23548 23772 23604 23774
rect 19852 22482 19908 22484
rect 19852 22430 19854 22482
rect 19854 22430 19906 22482
rect 19906 22430 19908 22482
rect 19852 22428 19908 22430
rect 21420 22482 21476 22484
rect 21420 22430 21422 22482
rect 21422 22430 21474 22482
rect 21474 22430 21476 22482
rect 21420 22428 21476 22430
rect 21980 22316 22036 22372
rect 18284 20636 18340 20692
rect 17612 20018 17668 20020
rect 17612 19966 17614 20018
rect 17614 19966 17666 20018
rect 17666 19966 17668 20018
rect 17612 19964 17668 19966
rect 18396 21756 18452 21812
rect 17948 17442 18004 17444
rect 17948 17390 17950 17442
rect 17950 17390 18002 17442
rect 18002 17390 18004 17442
rect 17948 17388 18004 17390
rect 18284 17164 18340 17220
rect 16604 16882 16660 16884
rect 16604 16830 16606 16882
rect 16606 16830 16658 16882
rect 16658 16830 16660 16882
rect 16604 16828 16660 16830
rect 17388 16658 17444 16660
rect 17388 16606 17390 16658
rect 17390 16606 17442 16658
rect 17442 16606 17444 16658
rect 17388 16604 17444 16606
rect 18844 20860 18900 20916
rect 19180 20690 19236 20692
rect 19180 20638 19182 20690
rect 19182 20638 19234 20690
rect 19234 20638 19236 20690
rect 19180 20636 19236 20638
rect 19180 20300 19236 20356
rect 18844 20130 18900 20132
rect 18844 20078 18846 20130
rect 18846 20078 18898 20130
rect 18898 20078 18900 20130
rect 18844 20076 18900 20078
rect 17948 16828 18004 16884
rect 18508 19964 18564 20020
rect 17836 16044 17892 16100
rect 16716 14588 16772 14644
rect 18620 17724 18676 17780
rect 19180 17778 19236 17780
rect 19180 17726 19182 17778
rect 19182 17726 19234 17778
rect 19234 17726 19236 17778
rect 19180 17724 19236 17726
rect 19404 20188 19460 20244
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19628 21532 19684 21588
rect 19628 20914 19684 20916
rect 19628 20862 19630 20914
rect 19630 20862 19682 20914
rect 19682 20862 19684 20914
rect 19628 20860 19684 20862
rect 19740 20524 19796 20580
rect 19852 20860 19908 20916
rect 19836 20410 19892 20412
rect 19628 20300 19684 20356
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19740 20188 19796 20244
rect 19628 19906 19684 19908
rect 19628 19854 19630 19906
rect 19630 19854 19682 19906
rect 19682 19854 19684 19906
rect 19628 19852 19684 19854
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 25228 34914 25284 34916
rect 25228 34862 25230 34914
rect 25230 34862 25282 34914
rect 25282 34862 25284 34914
rect 25228 34860 25284 34862
rect 27244 38834 27300 38836
rect 27244 38782 27246 38834
rect 27246 38782 27298 38834
rect 27298 38782 27300 38834
rect 27244 38780 27300 38782
rect 29708 38780 29764 38836
rect 26684 36876 26740 36932
rect 27132 36876 27188 36932
rect 30492 39506 30548 39508
rect 30492 39454 30494 39506
rect 30494 39454 30546 39506
rect 30546 39454 30548 39506
rect 30492 39452 30548 39454
rect 29820 38668 29876 38724
rect 30492 38668 30548 38724
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 33180 40402 33236 40404
rect 33180 40350 33182 40402
rect 33182 40350 33234 40402
rect 33234 40350 33236 40402
rect 33180 40348 33236 40350
rect 39900 41804 39956 41860
rect 36428 40402 36484 40404
rect 36428 40350 36430 40402
rect 36430 40350 36482 40402
rect 36482 40350 36484 40402
rect 36428 40348 36484 40350
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 38892 39394 38948 39396
rect 38892 39342 38894 39394
rect 38894 39342 38946 39394
rect 38946 39342 38948 39394
rect 38892 39340 38948 39342
rect 33852 39004 33908 39060
rect 38332 39058 38388 39060
rect 38332 39006 38334 39058
rect 38334 39006 38386 39058
rect 38386 39006 38388 39058
rect 38332 39004 38388 39006
rect 37324 38892 37380 38948
rect 31164 38668 31220 38724
rect 36764 38556 36820 38612
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34636 37884 34692 37940
rect 37212 37938 37268 37940
rect 37212 37886 37214 37938
rect 37214 37886 37266 37938
rect 37266 37886 37268 37938
rect 37212 37884 37268 37886
rect 37100 36988 37156 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 37100 36428 37156 36484
rect 26012 34636 26068 34692
rect 25340 34130 25396 34132
rect 25340 34078 25342 34130
rect 25342 34078 25394 34130
rect 25394 34078 25396 34130
rect 25340 34076 25396 34078
rect 25788 33964 25844 34020
rect 24892 33852 24948 33908
rect 25564 33906 25620 33908
rect 25564 33854 25566 33906
rect 25566 33854 25618 33906
rect 25618 33854 25620 33906
rect 25564 33852 25620 33854
rect 24892 32508 24948 32564
rect 25676 32450 25732 32452
rect 25676 32398 25678 32450
rect 25678 32398 25730 32450
rect 25730 32398 25732 32450
rect 25676 32396 25732 32398
rect 25788 31836 25844 31892
rect 25228 31778 25284 31780
rect 25228 31726 25230 31778
rect 25230 31726 25282 31778
rect 25282 31726 25284 31778
rect 25228 31724 25284 31726
rect 25564 31388 25620 31444
rect 36764 35698 36820 35700
rect 36764 35646 36766 35698
rect 36766 35646 36818 35698
rect 36818 35646 36820 35698
rect 36764 35644 36820 35646
rect 33404 35084 33460 35140
rect 31276 34802 31332 34804
rect 31276 34750 31278 34802
rect 31278 34750 31330 34802
rect 31330 34750 31332 34802
rect 31276 34748 31332 34750
rect 32060 34748 32116 34804
rect 30604 34636 30660 34692
rect 30828 34188 30884 34244
rect 26796 34076 26852 34132
rect 30156 34076 30212 34132
rect 29708 34018 29764 34020
rect 29708 33966 29710 34018
rect 29710 33966 29762 34018
rect 29762 33966 29764 34018
rect 29708 33964 29764 33966
rect 26348 31890 26404 31892
rect 26348 31838 26350 31890
rect 26350 31838 26402 31890
rect 26402 31838 26404 31890
rect 26348 31836 26404 31838
rect 26460 31724 26516 31780
rect 26124 31388 26180 31444
rect 26012 30994 26068 30996
rect 26012 30942 26014 30994
rect 26014 30942 26066 30994
rect 26066 30942 26068 30994
rect 26012 30940 26068 30942
rect 25564 30716 25620 30772
rect 25900 30098 25956 30100
rect 25900 30046 25902 30098
rect 25902 30046 25954 30098
rect 25954 30046 25956 30098
rect 25900 30044 25956 30046
rect 25788 29986 25844 29988
rect 25788 29934 25790 29986
rect 25790 29934 25842 29986
rect 25842 29934 25844 29986
rect 25788 29932 25844 29934
rect 29036 31106 29092 31108
rect 29036 31054 29038 31106
rect 29038 31054 29090 31106
rect 29090 31054 29092 31106
rect 29036 31052 29092 31054
rect 26908 30994 26964 30996
rect 26908 30942 26910 30994
rect 26910 30942 26962 30994
rect 26962 30942 26964 30994
rect 26908 30940 26964 30942
rect 26460 30716 26516 30772
rect 26684 30828 26740 30884
rect 26460 30492 26516 30548
rect 25564 29372 25620 29428
rect 24668 29314 24724 29316
rect 24668 29262 24670 29314
rect 24670 29262 24722 29314
rect 24722 29262 24724 29314
rect 24668 29260 24724 29262
rect 24220 21532 24276 21588
rect 23996 20242 24052 20244
rect 23996 20190 23998 20242
rect 23998 20190 24050 20242
rect 24050 20190 24052 20242
rect 23996 20188 24052 20190
rect 20636 19906 20692 19908
rect 20636 19854 20638 19906
rect 20638 19854 20690 19906
rect 20690 19854 20692 19906
rect 20636 19852 20692 19854
rect 20972 18396 21028 18452
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19292 17052 19348 17108
rect 19740 17052 19796 17108
rect 20636 17106 20692 17108
rect 20636 17054 20638 17106
rect 20638 17054 20690 17106
rect 20690 17054 20692 17106
rect 20636 17052 20692 17054
rect 20188 16828 20244 16884
rect 20972 16882 21028 16884
rect 20972 16830 20974 16882
rect 20974 16830 21026 16882
rect 21026 16830 21028 16882
rect 20972 16828 21028 16830
rect 21420 16716 21476 16772
rect 22988 20076 23044 20132
rect 23660 20130 23716 20132
rect 23660 20078 23662 20130
rect 23662 20078 23714 20130
rect 23714 20078 23716 20130
rect 23660 20076 23716 20078
rect 22988 18508 23044 18564
rect 22428 18450 22484 18452
rect 22428 18398 22430 18450
rect 22430 18398 22482 18450
rect 22482 18398 22484 18450
rect 22428 18396 22484 18398
rect 21644 16604 21700 16660
rect 19740 15820 19796 15876
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 22540 16604 22596 16660
rect 23660 17388 23716 17444
rect 24444 20748 24500 20804
rect 24556 20242 24612 20244
rect 24556 20190 24558 20242
rect 24558 20190 24610 20242
rect 24610 20190 24612 20242
rect 24556 20188 24612 20190
rect 23996 17554 24052 17556
rect 23996 17502 23998 17554
rect 23998 17502 24050 17554
rect 24050 17502 24052 17554
rect 23996 17500 24052 17502
rect 24556 17388 24612 17444
rect 24108 16940 24164 16996
rect 23772 16604 23828 16660
rect 20636 15148 20692 15204
rect 18508 14642 18564 14644
rect 18508 14590 18510 14642
rect 18510 14590 18562 14642
rect 18562 14590 18564 14642
rect 18508 14588 18564 14590
rect 19516 14588 19572 14644
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21756 15202 21812 15204
rect 21756 15150 21758 15202
rect 21758 15150 21810 15202
rect 21810 15150 21812 15202
rect 21756 15148 21812 15150
rect 22092 13580 22148 13636
rect 19852 13356 19908 13412
rect 20524 13356 20580 13412
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 17388 11394 17444 11396
rect 17388 11342 17390 11394
rect 17390 11342 17442 11394
rect 17442 11342 17444 11394
rect 17388 11340 17444 11342
rect 17612 11394 17668 11396
rect 17612 11342 17614 11394
rect 17614 11342 17666 11394
rect 17666 11342 17668 11394
rect 17612 11340 17668 11342
rect 16716 11282 16772 11284
rect 16716 11230 16718 11282
rect 16718 11230 16770 11282
rect 16770 11230 16772 11282
rect 16716 11228 16772 11230
rect 14588 9548 14644 9604
rect 17948 12012 18004 12068
rect 17836 11676 17892 11732
rect 17724 11228 17780 11284
rect 19852 12066 19908 12068
rect 19852 12014 19854 12066
rect 19854 12014 19906 12066
rect 19906 12014 19908 12066
rect 19852 12012 19908 12014
rect 18284 11676 18340 11732
rect 18060 11228 18116 11284
rect 18620 11282 18676 11284
rect 18620 11230 18622 11282
rect 18622 11230 18674 11282
rect 18674 11230 18676 11282
rect 18620 11228 18676 11230
rect 16604 10556 16660 10612
rect 17388 9660 17444 9716
rect 16492 9154 16548 9156
rect 16492 9102 16494 9154
rect 16494 9102 16546 9154
rect 16546 9102 16548 9154
rect 16492 9100 16548 9102
rect 18172 9714 18228 9716
rect 18172 9662 18174 9714
rect 18174 9662 18226 9714
rect 18226 9662 18228 9714
rect 18172 9660 18228 9662
rect 19068 9996 19124 10052
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 18844 9660 18900 9716
rect 17388 9100 17444 9156
rect 13580 8034 13636 8036
rect 13580 7982 13582 8034
rect 13582 7982 13634 8034
rect 13634 7982 13636 8034
rect 13580 7980 13636 7982
rect 13580 6690 13636 6692
rect 13580 6638 13582 6690
rect 13582 6638 13634 6690
rect 13634 6638 13636 6690
rect 13580 6636 13636 6638
rect 13692 6076 13748 6132
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19628 9212 19684 9268
rect 20524 9212 20580 9268
rect 21420 9266 21476 9268
rect 21420 9214 21422 9266
rect 21422 9214 21474 9266
rect 21474 9214 21476 9266
rect 21420 9212 21476 9214
rect 21868 9212 21924 9268
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 25228 27132 25284 27188
rect 25228 26796 25284 26852
rect 24892 26124 24948 26180
rect 24780 21532 24836 21588
rect 24780 20188 24836 20244
rect 25900 27020 25956 27076
rect 25564 26796 25620 26852
rect 25788 23212 25844 23268
rect 25676 22428 25732 22484
rect 25452 21586 25508 21588
rect 25452 21534 25454 21586
rect 25454 21534 25506 21586
rect 25506 21534 25508 21586
rect 25452 21532 25508 21534
rect 25452 20412 25508 20468
rect 25116 20188 25172 20244
rect 25676 17612 25732 17668
rect 25228 17554 25284 17556
rect 25228 17502 25230 17554
rect 25230 17502 25282 17554
rect 25282 17502 25284 17554
rect 25228 17500 25284 17502
rect 25676 16716 25732 16772
rect 25788 20412 25844 20468
rect 25228 15986 25284 15988
rect 25228 15934 25230 15986
rect 25230 15934 25282 15986
rect 25282 15934 25284 15986
rect 25228 15932 25284 15934
rect 25564 15820 25620 15876
rect 25340 15036 25396 15092
rect 22764 13634 22820 13636
rect 22764 13582 22766 13634
rect 22766 13582 22818 13634
rect 22818 13582 22820 13634
rect 22764 13580 22820 13582
rect 22876 13074 22932 13076
rect 22876 13022 22878 13074
rect 22878 13022 22930 13074
rect 22930 13022 22932 13074
rect 22876 13020 22932 13022
rect 23212 9884 23268 9940
rect 24332 13634 24388 13636
rect 24332 13582 24334 13634
rect 24334 13582 24386 13634
rect 24386 13582 24388 13634
rect 24332 13580 24388 13582
rect 24668 13522 24724 13524
rect 24668 13470 24670 13522
rect 24670 13470 24722 13522
rect 24722 13470 24724 13522
rect 24668 13468 24724 13470
rect 25452 13580 25508 13636
rect 24780 13020 24836 13076
rect 25340 13356 25396 13412
rect 30940 34130 30996 34132
rect 30940 34078 30942 34130
rect 30942 34078 30994 34130
rect 30994 34078 30996 34130
rect 30940 34076 30996 34078
rect 31388 34130 31444 34132
rect 31388 34078 31390 34130
rect 31390 34078 31442 34130
rect 31442 34078 31444 34130
rect 31388 34076 31444 34078
rect 31164 33964 31220 34020
rect 35980 35586 36036 35588
rect 35980 35534 35982 35586
rect 35982 35534 36034 35586
rect 36034 35534 36036 35586
rect 35980 35532 36036 35534
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 33852 34860 33908 34916
rect 35084 34860 35140 34916
rect 33852 34690 33908 34692
rect 33852 34638 33854 34690
rect 33854 34638 33906 34690
rect 33906 34638 33908 34690
rect 33852 34636 33908 34638
rect 34636 34636 34692 34692
rect 33404 34188 33460 34244
rect 31836 33964 31892 34020
rect 32284 34076 32340 34132
rect 30156 33068 30212 33124
rect 30380 31778 30436 31780
rect 30380 31726 30382 31778
rect 30382 31726 30434 31778
rect 30434 31726 30436 31778
rect 30380 31724 30436 31726
rect 32396 34018 32452 34020
rect 32396 33966 32398 34018
rect 32398 33966 32450 34018
rect 32450 33966 32452 34018
rect 32396 33964 32452 33966
rect 34524 33964 34580 34020
rect 33740 32786 33796 32788
rect 33740 32734 33742 32786
rect 33742 32734 33794 32786
rect 33794 32734 33796 32786
rect 33740 32732 33796 32734
rect 34188 32732 34244 32788
rect 29596 30716 29652 30772
rect 26796 30492 26852 30548
rect 27244 29932 27300 29988
rect 27356 30044 27412 30100
rect 30268 30940 30324 30996
rect 31388 31724 31444 31780
rect 30492 30828 30548 30884
rect 30604 30210 30660 30212
rect 30604 30158 30606 30210
rect 30606 30158 30658 30210
rect 30658 30158 30660 30210
rect 30604 30156 30660 30158
rect 29708 29932 29764 29988
rect 29820 29484 29876 29540
rect 27356 29036 27412 29092
rect 30380 29036 30436 29092
rect 30716 27298 30772 27300
rect 30716 27246 30718 27298
rect 30718 27246 30770 27298
rect 30770 27246 30772 27298
rect 30716 27244 30772 27246
rect 27020 26908 27076 26964
rect 30044 26962 30100 26964
rect 30044 26910 30046 26962
rect 30046 26910 30098 26962
rect 30098 26910 30100 26962
rect 30044 26908 30100 26910
rect 31276 30882 31332 30884
rect 31276 30830 31278 30882
rect 31278 30830 31330 30882
rect 31330 30830 31332 30882
rect 31276 30828 31332 30830
rect 31276 30210 31332 30212
rect 31276 30158 31278 30210
rect 31278 30158 31330 30210
rect 31330 30158 31332 30210
rect 31276 30156 31332 30158
rect 31052 29426 31108 29428
rect 31052 29374 31054 29426
rect 31054 29374 31106 29426
rect 31106 29374 31108 29426
rect 31052 29372 31108 29374
rect 30044 26348 30100 26404
rect 29820 26236 29876 26292
rect 29484 26124 29540 26180
rect 27692 24892 27748 24948
rect 29260 24946 29316 24948
rect 29260 24894 29262 24946
rect 29262 24894 29314 24946
rect 29314 24894 29316 24946
rect 29260 24892 29316 24894
rect 28700 24834 28756 24836
rect 28700 24782 28702 24834
rect 28702 24782 28754 24834
rect 28754 24782 28756 24834
rect 28700 24780 28756 24782
rect 28588 24722 28644 24724
rect 28588 24670 28590 24722
rect 28590 24670 28642 24722
rect 28642 24670 28644 24722
rect 28588 24668 28644 24670
rect 28252 23154 28308 23156
rect 28252 23102 28254 23154
rect 28254 23102 28306 23154
rect 28306 23102 28308 23154
rect 28252 23100 28308 23102
rect 26684 22482 26740 22484
rect 26684 22430 26686 22482
rect 26686 22430 26738 22482
rect 26738 22430 26740 22482
rect 26684 22428 26740 22430
rect 26124 21474 26180 21476
rect 26124 21422 26126 21474
rect 26126 21422 26178 21474
rect 26178 21422 26180 21474
rect 26124 21420 26180 21422
rect 27020 21420 27076 21476
rect 30268 26178 30324 26180
rect 30268 26126 30270 26178
rect 30270 26126 30322 26178
rect 30322 26126 30324 26178
rect 30268 26124 30324 26126
rect 29932 24834 29988 24836
rect 29932 24782 29934 24834
rect 29934 24782 29986 24834
rect 29986 24782 29988 24834
rect 29932 24780 29988 24782
rect 29596 24668 29652 24724
rect 31948 30156 32004 30212
rect 34076 31666 34132 31668
rect 34076 31614 34078 31666
rect 34078 31614 34130 31666
rect 34130 31614 34132 31666
rect 34076 31612 34132 31614
rect 32396 30156 32452 30212
rect 32060 30098 32116 30100
rect 32060 30046 32062 30098
rect 32062 30046 32114 30098
rect 32114 30046 32116 30098
rect 32060 30044 32116 30046
rect 33964 30716 34020 30772
rect 31276 29484 31332 29540
rect 31500 29426 31556 29428
rect 31500 29374 31502 29426
rect 31502 29374 31554 29426
rect 31554 29374 31556 29426
rect 31500 29372 31556 29374
rect 33628 29538 33684 29540
rect 33628 29486 33630 29538
rect 33630 29486 33682 29538
rect 33682 29486 33684 29538
rect 33628 29484 33684 29486
rect 33292 29426 33348 29428
rect 33292 29374 33294 29426
rect 33294 29374 33346 29426
rect 33346 29374 33348 29426
rect 33292 29372 33348 29374
rect 31836 27692 31892 27748
rect 31836 27244 31892 27300
rect 30716 26290 30772 26292
rect 30716 26238 30718 26290
rect 30718 26238 30770 26290
rect 30770 26238 30772 26290
rect 30716 26236 30772 26238
rect 31276 26290 31332 26292
rect 31276 26238 31278 26290
rect 31278 26238 31330 26290
rect 31330 26238 31332 26290
rect 31276 26236 31332 26238
rect 31612 26402 31668 26404
rect 31612 26350 31614 26402
rect 31614 26350 31666 26402
rect 31666 26350 31668 26402
rect 31612 26348 31668 26350
rect 31612 25228 31668 25284
rect 30380 23100 30436 23156
rect 34076 26908 34132 26964
rect 34860 31612 34916 31668
rect 34748 31218 34804 31220
rect 34748 31166 34750 31218
rect 34750 31166 34802 31218
rect 34802 31166 34804 31218
rect 34748 31164 34804 31166
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35756 32732 35812 32788
rect 36316 32732 36372 32788
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35532 31218 35588 31220
rect 35532 31166 35534 31218
rect 35534 31166 35586 31218
rect 35586 31166 35588 31218
rect 35532 31164 35588 31166
rect 34860 30994 34916 30996
rect 34860 30942 34862 30994
rect 34862 30942 34914 30994
rect 34914 30942 34916 30994
rect 34860 30940 34916 30942
rect 35084 30828 35140 30884
rect 35756 30994 35812 30996
rect 35756 30942 35758 30994
rect 35758 30942 35810 30994
rect 35810 30942 35812 30994
rect 35756 30940 35812 30942
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34860 27746 34916 27748
rect 34860 27694 34862 27746
rect 34862 27694 34914 27746
rect 34914 27694 34916 27746
rect 34860 27692 34916 27694
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34412 27020 34468 27076
rect 31948 26290 32004 26292
rect 31948 26238 31950 26290
rect 31950 26238 32002 26290
rect 32002 26238 32004 26290
rect 31948 26236 32004 26238
rect 32396 25900 32452 25956
rect 33852 24780 33908 24836
rect 31724 23324 31780 23380
rect 32396 23324 32452 23380
rect 28700 21474 28756 21476
rect 28700 21422 28702 21474
rect 28702 21422 28754 21474
rect 28754 21422 28756 21474
rect 28700 21420 28756 21422
rect 29596 21420 29652 21476
rect 31724 22876 31780 22932
rect 32284 22876 32340 22932
rect 26684 20802 26740 20804
rect 26684 20750 26686 20802
rect 26686 20750 26738 20802
rect 26738 20750 26740 20802
rect 26684 20748 26740 20750
rect 29820 20802 29876 20804
rect 29820 20750 29822 20802
rect 29822 20750 29874 20802
rect 29874 20750 29876 20802
rect 29820 20748 29876 20750
rect 33628 22370 33684 22372
rect 33628 22318 33630 22370
rect 33630 22318 33682 22370
rect 33682 22318 33684 22370
rect 33628 22316 33684 22318
rect 33180 21474 33236 21476
rect 33180 21422 33182 21474
rect 33182 21422 33234 21474
rect 33234 21422 33236 21474
rect 33180 21420 33236 21422
rect 31948 19068 32004 19124
rect 25900 17724 25956 17780
rect 26572 16828 26628 16884
rect 27804 17442 27860 17444
rect 27804 17390 27806 17442
rect 27806 17390 27858 17442
rect 27858 17390 27860 17442
rect 27804 17388 27860 17390
rect 27692 16994 27748 16996
rect 27692 16942 27694 16994
rect 27694 16942 27746 16994
rect 27746 16942 27748 16994
rect 27692 16940 27748 16942
rect 27356 16716 27412 16772
rect 26908 16098 26964 16100
rect 26908 16046 26910 16098
rect 26910 16046 26962 16098
rect 26962 16046 26964 16098
rect 26908 16044 26964 16046
rect 26796 15820 26852 15876
rect 26012 15036 26068 15092
rect 25564 13522 25620 13524
rect 25564 13470 25566 13522
rect 25566 13470 25618 13522
rect 25618 13470 25620 13522
rect 25564 13468 25620 13470
rect 26124 13356 26180 13412
rect 26236 12124 26292 12180
rect 26908 12124 26964 12180
rect 25340 11340 25396 11396
rect 25788 11228 25844 11284
rect 24108 9938 24164 9940
rect 24108 9886 24110 9938
rect 24110 9886 24162 9938
rect 24162 9886 24164 9938
rect 24108 9884 24164 9886
rect 22988 8652 23044 8708
rect 23436 9100 23492 9156
rect 26348 9324 26404 9380
rect 25340 9154 25396 9156
rect 25340 9102 25342 9154
rect 25342 9102 25394 9154
rect 25394 9102 25396 9154
rect 25340 9100 25396 9102
rect 24668 8988 24724 9044
rect 25676 9042 25732 9044
rect 25676 8990 25678 9042
rect 25678 8990 25730 9042
rect 25730 8990 25732 9042
rect 25676 8988 25732 8990
rect 23660 8652 23716 8708
rect 23212 8204 23268 8260
rect 26348 8428 26404 8484
rect 23548 8258 23604 8260
rect 23548 8206 23550 8258
rect 23550 8206 23602 8258
rect 23602 8206 23604 8258
rect 23548 8204 23604 8206
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 15372 6130 15428 6132
rect 15372 6078 15374 6130
rect 15374 6078 15426 6130
rect 15426 6078 15428 6130
rect 15372 6076 15428 6078
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 25788 6524 25844 6580
rect 24556 5964 24612 6020
rect 23324 5794 23380 5796
rect 23324 5742 23326 5794
rect 23326 5742 23378 5794
rect 23378 5742 23380 5794
rect 23324 5740 23380 5742
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 26236 6578 26292 6580
rect 26236 6526 26238 6578
rect 26238 6526 26290 6578
rect 26290 6526 26292 6578
rect 26236 6524 26292 6526
rect 25676 5740 25732 5796
rect 26796 6914 26852 6916
rect 26796 6862 26798 6914
rect 26798 6862 26850 6914
rect 26850 6862 26852 6914
rect 26796 6860 26852 6862
rect 27020 11228 27076 11284
rect 28588 17442 28644 17444
rect 28588 17390 28590 17442
rect 28590 17390 28642 17442
rect 28642 17390 28644 17442
rect 28588 17388 28644 17390
rect 28364 16716 28420 16772
rect 30044 18338 30100 18340
rect 30044 18286 30046 18338
rect 30046 18286 30098 18338
rect 30098 18286 30100 18338
rect 30044 18284 30100 18286
rect 31276 18284 31332 18340
rect 29484 17724 29540 17780
rect 28364 16044 28420 16100
rect 29148 16098 29204 16100
rect 29148 16046 29150 16098
rect 29150 16046 29202 16098
rect 29202 16046 29204 16098
rect 29148 16044 29204 16046
rect 29372 15874 29428 15876
rect 29372 15822 29374 15874
rect 29374 15822 29426 15874
rect 29426 15822 29428 15874
rect 29372 15820 29428 15822
rect 29260 15260 29316 15316
rect 30156 17388 30212 17444
rect 33852 17612 33908 17668
rect 31948 17052 32004 17108
rect 32060 16940 32116 16996
rect 30156 16828 30212 16884
rect 32508 16994 32564 16996
rect 32508 16942 32510 16994
rect 32510 16942 32562 16994
rect 32562 16942 32564 16994
rect 32508 16940 32564 16942
rect 33628 16940 33684 16996
rect 33292 16882 33348 16884
rect 33292 16830 33294 16882
rect 33294 16830 33346 16882
rect 33346 16830 33348 16882
rect 33292 16828 33348 16830
rect 29484 15484 29540 15540
rect 30604 15538 30660 15540
rect 30604 15486 30606 15538
rect 30606 15486 30658 15538
rect 30658 15486 30660 15538
rect 30604 15484 30660 15486
rect 30380 15314 30436 15316
rect 30380 15262 30382 15314
rect 30382 15262 30434 15314
rect 30434 15262 30436 15314
rect 30380 15260 30436 15262
rect 29820 15202 29876 15204
rect 29820 15150 29822 15202
rect 29822 15150 29874 15202
rect 29874 15150 29876 15202
rect 29820 15148 29876 15150
rect 29484 13356 29540 13412
rect 29708 12962 29764 12964
rect 29708 12910 29710 12962
rect 29710 12910 29762 12962
rect 29762 12910 29764 12962
rect 29708 12908 29764 12910
rect 30828 13468 30884 13524
rect 28140 12178 28196 12180
rect 28140 12126 28142 12178
rect 28142 12126 28194 12178
rect 28194 12126 28196 12178
rect 28140 12124 28196 12126
rect 29596 10668 29652 10724
rect 28924 10556 28980 10612
rect 27468 9772 27524 9828
rect 30380 12962 30436 12964
rect 30380 12910 30382 12962
rect 30382 12910 30434 12962
rect 30434 12910 30436 12962
rect 30380 12908 30436 12910
rect 32284 13468 32340 13524
rect 37548 38668 37604 38724
rect 37996 38610 38052 38612
rect 37996 38558 37998 38610
rect 37998 38558 38050 38610
rect 38050 38558 38052 38610
rect 37996 38556 38052 38558
rect 37772 37884 37828 37940
rect 37660 36482 37716 36484
rect 37660 36430 37662 36482
rect 37662 36430 37714 36482
rect 37714 36430 37716 36482
rect 37660 36428 37716 36430
rect 37996 36258 38052 36260
rect 37996 36206 37998 36258
rect 37998 36206 38050 36258
rect 38050 36206 38052 36258
rect 37996 36204 38052 36206
rect 37212 35586 37268 35588
rect 37212 35534 37214 35586
rect 37214 35534 37266 35586
rect 37266 35534 37268 35586
rect 37212 35532 37268 35534
rect 38108 35698 38164 35700
rect 38108 35646 38110 35698
rect 38110 35646 38162 35698
rect 38162 35646 38164 35698
rect 38108 35644 38164 35646
rect 37548 35532 37604 35588
rect 37100 34860 37156 34916
rect 37212 31948 37268 32004
rect 37212 31666 37268 31668
rect 37212 31614 37214 31666
rect 37214 31614 37266 31666
rect 37266 31614 37268 31666
rect 37212 31612 37268 31614
rect 36988 30210 37044 30212
rect 36988 30158 36990 30210
rect 36990 30158 37042 30210
rect 37042 30158 37044 30210
rect 36988 30156 37044 30158
rect 37100 30098 37156 30100
rect 37100 30046 37102 30098
rect 37102 30046 37154 30098
rect 37154 30046 37156 30098
rect 37100 30044 37156 30046
rect 37100 28588 37156 28644
rect 38780 38722 38836 38724
rect 38780 38670 38782 38722
rect 38782 38670 38834 38722
rect 38834 38670 38836 38722
rect 38780 38668 38836 38670
rect 39900 38946 39956 38948
rect 39900 38894 39902 38946
rect 39902 38894 39954 38946
rect 39954 38894 39956 38946
rect 39900 38892 39956 38894
rect 39228 37884 39284 37940
rect 40124 38834 40180 38836
rect 40124 38782 40126 38834
rect 40126 38782 40178 38834
rect 40178 38782 40180 38834
rect 40124 38780 40180 38782
rect 41132 41858 41188 41860
rect 41132 41806 41134 41858
rect 41134 41806 41186 41858
rect 41186 41806 41188 41858
rect 41132 41804 41188 41806
rect 41580 40236 41636 40292
rect 40460 39340 40516 39396
rect 40908 39004 40964 39060
rect 38780 35644 38836 35700
rect 39340 36988 39396 37044
rect 38220 34636 38276 34692
rect 37884 30044 37940 30100
rect 38108 31836 38164 31892
rect 37548 28700 37604 28756
rect 37772 28642 37828 28644
rect 37772 28590 37774 28642
rect 37774 28590 37826 28642
rect 37826 28590 37828 28642
rect 37772 28588 37828 28590
rect 40348 37938 40404 37940
rect 40348 37886 40350 37938
rect 40350 37886 40402 37938
rect 40402 37886 40404 37938
rect 40348 37884 40404 37886
rect 40236 36988 40292 37044
rect 40012 36204 40068 36260
rect 39452 35698 39508 35700
rect 39452 35646 39454 35698
rect 39454 35646 39506 35698
rect 39506 35646 39508 35698
rect 39452 35644 39508 35646
rect 39788 35532 39844 35588
rect 40236 35586 40292 35588
rect 40236 35534 40238 35586
rect 40238 35534 40290 35586
rect 40290 35534 40292 35586
rect 40236 35532 40292 35534
rect 40348 35084 40404 35140
rect 40796 36258 40852 36260
rect 40796 36206 40798 36258
rect 40798 36206 40850 36258
rect 40850 36206 40852 36258
rect 40796 36204 40852 36206
rect 40684 36092 40740 36148
rect 41356 39058 41412 39060
rect 41356 39006 41358 39058
rect 41358 39006 41410 39058
rect 41410 39006 41412 39058
rect 41356 39004 41412 39006
rect 41692 39058 41748 39060
rect 41692 39006 41694 39058
rect 41694 39006 41746 39058
rect 41746 39006 41748 39058
rect 41692 39004 41748 39006
rect 41580 38892 41636 38948
rect 41132 37938 41188 37940
rect 41132 37886 41134 37938
rect 41134 37886 41186 37938
rect 41186 37886 41188 37938
rect 41132 37884 41188 37886
rect 43932 40290 43988 40292
rect 43932 40238 43934 40290
rect 43934 40238 43986 40290
rect 43986 40238 43988 40290
rect 43932 40236 43988 40238
rect 42028 39340 42084 39396
rect 42140 38834 42196 38836
rect 42140 38782 42142 38834
rect 42142 38782 42194 38834
rect 42194 38782 42196 38834
rect 42140 38780 42196 38782
rect 41132 36204 41188 36260
rect 43820 36204 43876 36260
rect 41020 36092 41076 36148
rect 40348 34690 40404 34692
rect 40348 34638 40350 34690
rect 40350 34638 40402 34690
rect 40402 34638 40404 34690
rect 40348 34636 40404 34638
rect 40012 33346 40068 33348
rect 40012 33294 40014 33346
rect 40014 33294 40066 33346
rect 40066 33294 40068 33346
rect 40012 33292 40068 33294
rect 39340 31612 39396 31668
rect 39564 31836 39620 31892
rect 40460 33404 40516 33460
rect 40908 35698 40964 35700
rect 40908 35646 40910 35698
rect 40910 35646 40962 35698
rect 40962 35646 40964 35698
rect 40908 35644 40964 35646
rect 40348 31836 40404 31892
rect 40908 33346 40964 33348
rect 40908 33294 40910 33346
rect 40910 33294 40962 33346
rect 40962 33294 40964 33346
rect 40908 33292 40964 33294
rect 40572 31612 40628 31668
rect 38556 29372 38612 29428
rect 36092 28364 36148 28420
rect 35756 27692 35812 27748
rect 35756 27074 35812 27076
rect 35756 27022 35758 27074
rect 35758 27022 35810 27074
rect 35810 27022 35812 27074
rect 35756 27020 35812 27022
rect 37996 28418 38052 28420
rect 37996 28366 37998 28418
rect 37998 28366 38050 28418
rect 38050 28366 38052 28418
rect 37996 28364 38052 28366
rect 35644 26514 35700 26516
rect 35644 26462 35646 26514
rect 35646 26462 35698 26514
rect 35698 26462 35700 26514
rect 35644 26460 35700 26462
rect 34860 25900 34916 25956
rect 34300 21756 34356 21812
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35532 24892 35588 24948
rect 35644 25228 35700 25284
rect 37436 27020 37492 27076
rect 36428 26460 36484 26516
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 36092 23660 36148 23716
rect 35308 23266 35364 23268
rect 35308 23214 35310 23266
rect 35310 23214 35362 23266
rect 35362 23214 35364 23266
rect 35308 23212 35364 23214
rect 35644 23154 35700 23156
rect 35644 23102 35646 23154
rect 35646 23102 35698 23154
rect 35698 23102 35700 23154
rect 35644 23100 35700 23102
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35420 22540 35476 22596
rect 35308 21810 35364 21812
rect 35308 21758 35310 21810
rect 35310 21758 35362 21810
rect 35362 21758 35364 21810
rect 35308 21756 35364 21758
rect 36204 23436 36260 23492
rect 36092 22540 36148 22596
rect 37884 25618 37940 25620
rect 37884 25566 37886 25618
rect 37886 25566 37938 25618
rect 37938 25566 37940 25618
rect 37884 25564 37940 25566
rect 38668 27746 38724 27748
rect 38668 27694 38670 27746
rect 38670 27694 38722 27746
rect 38722 27694 38724 27746
rect 38668 27692 38724 27694
rect 38220 25564 38276 25620
rect 38668 25564 38724 25620
rect 36540 24946 36596 24948
rect 36540 24894 36542 24946
rect 36542 24894 36594 24946
rect 36594 24894 36596 24946
rect 36540 24892 36596 24894
rect 39788 29484 39844 29540
rect 39004 28700 39060 28756
rect 39340 27692 39396 27748
rect 39228 24668 39284 24724
rect 36540 23660 36596 23716
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35644 19010 35700 19012
rect 35644 18958 35646 19010
rect 35646 18958 35698 19010
rect 35698 18958 35700 19010
rect 35644 18956 35700 18958
rect 35756 18508 35812 18564
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35308 17666 35364 17668
rect 35308 17614 35310 17666
rect 35310 17614 35362 17666
rect 35362 17614 35364 17666
rect 35308 17612 35364 17614
rect 36092 19010 36148 19012
rect 36092 18958 36094 19010
rect 36094 18958 36146 19010
rect 36146 18958 36148 19010
rect 36092 18956 36148 18958
rect 36428 18396 36484 18452
rect 36428 17778 36484 17780
rect 36428 17726 36430 17778
rect 36430 17726 36482 17778
rect 36482 17726 36484 17778
rect 36428 17724 36484 17726
rect 35868 17612 35924 17668
rect 30268 12850 30324 12852
rect 30268 12798 30270 12850
rect 30270 12798 30322 12850
rect 30322 12798 30324 12850
rect 30268 12796 30324 12798
rect 30604 12348 30660 12404
rect 32956 12908 33012 12964
rect 31948 12796 32004 12852
rect 31388 12178 31444 12180
rect 31388 12126 31390 12178
rect 31390 12126 31442 12178
rect 31442 12126 31444 12178
rect 31388 12124 31444 12126
rect 30492 11282 30548 11284
rect 30492 11230 30494 11282
rect 30494 11230 30546 11282
rect 30546 11230 30548 11282
rect 30492 11228 30548 11230
rect 30380 10722 30436 10724
rect 30380 10670 30382 10722
rect 30382 10670 30434 10722
rect 30434 10670 30436 10722
rect 30380 10668 30436 10670
rect 32844 12850 32900 12852
rect 32844 12798 32846 12850
rect 32846 12798 32898 12850
rect 32898 12798 32900 12850
rect 32844 12796 32900 12798
rect 32060 12348 32116 12404
rect 32060 11228 32116 11284
rect 32396 12012 32452 12068
rect 31948 10668 32004 10724
rect 30044 10610 30100 10612
rect 30044 10558 30046 10610
rect 30046 10558 30098 10610
rect 30098 10558 30100 10610
rect 30044 10556 30100 10558
rect 29372 9826 29428 9828
rect 29372 9774 29374 9826
rect 29374 9774 29426 9826
rect 29426 9774 29428 9826
rect 29372 9772 29428 9774
rect 27580 9154 27636 9156
rect 27580 9102 27582 9154
rect 27582 9102 27634 9154
rect 27634 9102 27636 9154
rect 27580 9100 27636 9102
rect 28364 9154 28420 9156
rect 28364 9102 28366 9154
rect 28366 9102 28418 9154
rect 28418 9102 28420 9154
rect 28364 9100 28420 9102
rect 27132 8652 27188 8708
rect 27580 8652 27636 8708
rect 28252 8316 28308 8372
rect 27804 8258 27860 8260
rect 27804 8206 27806 8258
rect 27806 8206 27858 8258
rect 27858 8206 27860 8258
rect 27804 8204 27860 8206
rect 26572 6300 26628 6356
rect 26460 6018 26516 6020
rect 26460 5966 26462 6018
rect 26462 5966 26514 6018
rect 26514 5966 26516 6018
rect 26460 5964 26516 5966
rect 26908 6300 26964 6356
rect 26908 5628 26964 5684
rect 27132 6578 27188 6580
rect 27132 6526 27134 6578
rect 27134 6526 27186 6578
rect 27186 6526 27188 6578
rect 27132 6524 27188 6526
rect 28476 8204 28532 8260
rect 28700 8988 28756 9044
rect 29484 8370 29540 8372
rect 29484 8318 29486 8370
rect 29486 8318 29538 8370
rect 29538 8318 29540 8370
rect 29484 8316 29540 8318
rect 29932 8316 29988 8372
rect 31612 8370 31668 8372
rect 31612 8318 31614 8370
rect 31614 8318 31666 8370
rect 31666 8318 31668 8370
rect 31612 8316 31668 8318
rect 32508 11394 32564 11396
rect 32508 11342 32510 11394
rect 32510 11342 32562 11394
rect 32562 11342 32564 11394
rect 32508 11340 32564 11342
rect 33068 12738 33124 12740
rect 33068 12686 33070 12738
rect 33070 12686 33122 12738
rect 33122 12686 33124 12738
rect 33068 12684 33124 12686
rect 33068 12348 33124 12404
rect 33964 12962 34020 12964
rect 33964 12910 33966 12962
rect 33966 12910 34018 12962
rect 34018 12910 34020 12962
rect 33964 12908 34020 12910
rect 33740 12348 33796 12404
rect 33516 11394 33572 11396
rect 33516 11342 33518 11394
rect 33518 11342 33570 11394
rect 33570 11342 33572 11394
rect 33516 11340 33572 11342
rect 34748 11340 34804 11396
rect 35980 17554 36036 17556
rect 35980 17502 35982 17554
rect 35982 17502 36034 17554
rect 36034 17502 36036 17554
rect 35980 17500 36036 17502
rect 37212 23100 37268 23156
rect 36540 17500 36596 17556
rect 36764 22316 36820 22372
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 37100 22370 37156 22372
rect 37100 22318 37102 22370
rect 37102 22318 37154 22370
rect 37154 22318 37156 22370
rect 37100 22316 37156 22318
rect 39004 22876 39060 22932
rect 41692 35586 41748 35588
rect 41692 35534 41694 35586
rect 41694 35534 41746 35586
rect 41746 35534 41748 35586
rect 41692 35532 41748 35534
rect 43820 33458 43876 33460
rect 43820 33406 43822 33458
rect 43822 33406 43874 33458
rect 43874 33406 43876 33458
rect 43820 33404 43876 33406
rect 41020 32844 41076 32900
rect 41692 32786 41748 32788
rect 41692 32734 41694 32786
rect 41694 32734 41746 32786
rect 41746 32734 41748 32786
rect 41692 32732 41748 32734
rect 41580 31666 41636 31668
rect 41580 31614 41582 31666
rect 41582 31614 41634 31666
rect 41634 31614 41636 31666
rect 41580 31612 41636 31614
rect 41692 29708 41748 29764
rect 42476 29708 42532 29764
rect 40348 29426 40404 29428
rect 40348 29374 40350 29426
rect 40350 29374 40402 29426
rect 40402 29374 40404 29426
rect 40348 29372 40404 29374
rect 41468 28700 41524 28756
rect 42588 29260 42644 29316
rect 40572 28476 40628 28532
rect 40236 25618 40292 25620
rect 40236 25566 40238 25618
rect 40238 25566 40290 25618
rect 40290 25566 40292 25618
rect 40236 25564 40292 25566
rect 39788 24892 39844 24948
rect 41132 25564 41188 25620
rect 40012 24834 40068 24836
rect 40012 24782 40014 24834
rect 40014 24782 40066 24834
rect 40066 24782 40068 24834
rect 40012 24780 40068 24782
rect 39900 24108 39956 24164
rect 39676 23154 39732 23156
rect 39676 23102 39678 23154
rect 39678 23102 39730 23154
rect 39730 23102 39732 23154
rect 39676 23100 39732 23102
rect 39116 20412 39172 20468
rect 39564 20076 39620 20132
rect 38892 19122 38948 19124
rect 38892 19070 38894 19122
rect 38894 19070 38946 19122
rect 38946 19070 38948 19122
rect 38892 19068 38948 19070
rect 40684 25452 40740 25508
rect 42364 28530 42420 28532
rect 42364 28478 42366 28530
rect 42366 28478 42418 28530
rect 42418 28478 42420 28530
rect 42364 28476 42420 28478
rect 43820 29314 43876 29316
rect 43820 29262 43822 29314
rect 43822 29262 43874 29314
rect 43874 29262 43876 29314
rect 43820 29260 43876 29262
rect 44044 25618 44100 25620
rect 44044 25566 44046 25618
rect 44046 25566 44098 25618
rect 44098 25566 44100 25618
rect 44044 25564 44100 25566
rect 42364 24780 42420 24836
rect 41804 24668 41860 24724
rect 42028 24108 42084 24164
rect 40572 20076 40628 20132
rect 39900 19068 39956 19124
rect 41692 19964 41748 20020
rect 37324 17612 37380 17668
rect 36988 17554 37044 17556
rect 36988 17502 36990 17554
rect 36990 17502 37042 17554
rect 37042 17502 37044 17554
rect 36988 17500 37044 17502
rect 41804 19852 41860 19908
rect 42364 19852 42420 19908
rect 41692 19180 41748 19236
rect 41132 19068 41188 19124
rect 41020 18562 41076 18564
rect 41020 18510 41022 18562
rect 41022 18510 41074 18562
rect 41074 18510 41076 18562
rect 41020 18508 41076 18510
rect 44044 19906 44100 19908
rect 44044 19854 44046 19906
rect 44046 19854 44098 19906
rect 44098 19854 44100 19906
rect 44044 19852 44100 19854
rect 42476 19234 42532 19236
rect 42476 19182 42478 19234
rect 42478 19182 42530 19234
rect 42530 19182 42532 19234
rect 42476 19180 42532 19182
rect 41580 18396 41636 18452
rect 43372 18396 43428 18452
rect 36764 16994 36820 16996
rect 36764 16942 36766 16994
rect 36766 16942 36818 16994
rect 36818 16942 36820 16994
rect 36764 16940 36820 16942
rect 37212 17442 37268 17444
rect 37212 17390 37214 17442
rect 37214 17390 37266 17442
rect 37266 17390 37268 17442
rect 37212 17388 37268 17390
rect 37100 15820 37156 15876
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 40460 17442 40516 17444
rect 40460 17390 40462 17442
rect 40462 17390 40514 17442
rect 40514 17390 40516 17442
rect 40460 17388 40516 17390
rect 40124 15874 40180 15876
rect 40124 15822 40126 15874
rect 40126 15822 40178 15874
rect 40178 15822 40180 15874
rect 40124 15820 40180 15822
rect 40460 15820 40516 15876
rect 36428 14306 36484 14308
rect 36428 14254 36430 14306
rect 36430 14254 36482 14306
rect 36482 14254 36484 14306
rect 36428 14252 36484 14254
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 33068 11282 33124 11284
rect 33068 11230 33070 11282
rect 33070 11230 33122 11282
rect 33122 11230 33124 11282
rect 33068 11228 33124 11230
rect 35196 12684 35252 12740
rect 35868 12012 35924 12068
rect 37324 14252 37380 14308
rect 36428 12066 36484 12068
rect 36428 12014 36430 12066
rect 36430 12014 36482 12066
rect 36482 12014 36484 12066
rect 36428 12012 36484 12014
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34972 8428 35028 8484
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 27804 6860 27860 6916
rect 27804 6578 27860 6580
rect 27804 6526 27806 6578
rect 27806 6526 27858 6578
rect 27858 6526 27860 6578
rect 27804 6524 27860 6526
rect 27020 4508 27076 4564
rect 27804 5682 27860 5684
rect 27804 5630 27806 5682
rect 27806 5630 27858 5682
rect 27858 5630 27860 5682
rect 27804 5628 27860 5630
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 30268 4562 30324 4564
rect 30268 4510 30270 4562
rect 30270 4510 30322 4562
rect 30322 4510 30324 4562
rect 30268 4508 30324 4510
rect 27468 4172 27524 4228
rect 29820 4226 29876 4228
rect 29820 4174 29822 4226
rect 29822 4174 29874 4226
rect 29874 4174 29876 4226
rect 29820 4172 29876 4174
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
<< metal3 >>
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 12674 41916 12684 41972
rect 12740 41916 13468 41972
rect 13524 41916 13534 41972
rect 16146 41916 16156 41972
rect 16212 41916 17276 41972
rect 17332 41916 17342 41972
rect 13234 41804 13244 41860
rect 13300 41804 14476 41860
rect 14532 41804 14542 41860
rect 24658 41804 24668 41860
rect 24724 41804 25900 41860
rect 25956 41804 25966 41860
rect 39890 41804 39900 41860
rect 39956 41804 41132 41860
rect 41188 41804 41198 41860
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 5618 40460 5628 40516
rect 5684 40460 8764 40516
rect 8820 40460 20636 40516
rect 20692 40460 20702 40516
rect 4946 40348 4956 40404
rect 5012 40348 5740 40404
rect 5796 40348 8316 40404
rect 8372 40348 9772 40404
rect 9828 40348 10444 40404
rect 10500 40348 10510 40404
rect 13346 40348 13356 40404
rect 13412 40348 16940 40404
rect 16996 40348 17612 40404
rect 17668 40348 17678 40404
rect 20066 40348 20076 40404
rect 20132 40348 23660 40404
rect 23716 40348 23726 40404
rect 25778 40348 25788 40404
rect 25844 40348 28476 40404
rect 28532 40348 28542 40404
rect 31154 40348 31164 40404
rect 31220 40348 33180 40404
rect 33236 40348 36428 40404
rect 36484 40348 36494 40404
rect 10546 40236 10556 40292
rect 10612 40236 18956 40292
rect 19012 40236 19022 40292
rect 24210 40236 24220 40292
rect 24276 40236 25676 40292
rect 25732 40236 25742 40292
rect 41570 40236 41580 40292
rect 41636 40236 43932 40292
rect 43988 40236 43998 40292
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 4722 39676 4732 39732
rect 4788 39676 6972 39732
rect 7028 39676 7038 39732
rect 7746 39676 7756 39732
rect 7812 39676 8764 39732
rect 8820 39676 8830 39732
rect 26450 39564 26460 39620
rect 26516 39564 26908 39620
rect 26964 39564 27804 39620
rect 27860 39564 29820 39620
rect 29876 39564 29886 39620
rect 18498 39452 18508 39508
rect 18564 39452 19068 39508
rect 19124 39452 19852 39508
rect 19908 39452 20188 39508
rect 20244 39452 20254 39508
rect 23762 39452 23772 39508
rect 23828 39452 30492 39508
rect 30548 39452 30558 39508
rect 18274 39340 18284 39396
rect 18340 39340 18844 39396
rect 18900 39340 20076 39396
rect 20132 39340 26460 39396
rect 26516 39340 27132 39396
rect 27188 39340 27198 39396
rect 38882 39340 38892 39396
rect 38948 39340 40460 39396
rect 40516 39340 42028 39396
rect 42084 39340 42094 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 24770 39004 24780 39060
rect 24836 39004 33852 39060
rect 33908 39004 33918 39060
rect 38322 39004 38332 39060
rect 38388 39004 40908 39060
rect 40964 39004 41356 39060
rect 41412 39004 41692 39060
rect 41748 39004 41758 39060
rect 20514 38892 20524 38948
rect 20580 38892 24556 38948
rect 24612 38892 24622 38948
rect 37314 38892 37324 38948
rect 37380 38892 39900 38948
rect 39956 38892 41580 38948
rect 41636 38892 41646 38948
rect 20132 38724 20188 38836
rect 20244 38780 20254 38836
rect 23762 38780 23772 38836
rect 23828 38780 26124 38836
rect 26180 38780 27244 38836
rect 27300 38780 29708 38836
rect 29764 38780 29774 38836
rect 40114 38780 40124 38836
rect 40180 38780 42140 38836
rect 42196 38780 42206 38836
rect 16594 38668 16604 38724
rect 16660 38668 17948 38724
rect 18004 38668 20188 38724
rect 29810 38668 29820 38724
rect 29876 38668 30492 38724
rect 30548 38668 31164 38724
rect 31220 38668 31230 38724
rect 37538 38668 37548 38724
rect 37604 38668 38780 38724
rect 38836 38668 38846 38724
rect 14914 38556 14924 38612
rect 14980 38556 23548 38612
rect 23604 38556 23614 38612
rect 36754 38556 36764 38612
rect 36820 38556 37996 38612
rect 38052 38556 38062 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 20402 38220 20412 38276
rect 20468 38220 24220 38276
rect 24276 38220 25452 38276
rect 25508 38220 25518 38276
rect 1810 38108 1820 38164
rect 1876 38108 2268 38164
rect 2324 38108 5740 38164
rect 5796 38108 5806 38164
rect 11106 37996 11116 38052
rect 11172 37996 12908 38052
rect 12964 37996 14252 38052
rect 14308 37996 14318 38052
rect 2930 37884 2940 37940
rect 2996 37884 5068 37940
rect 5124 37884 5134 37940
rect 20066 37884 20076 37940
rect 20132 37884 20524 37940
rect 20580 37884 21420 37940
rect 21476 37884 21486 37940
rect 34626 37884 34636 37940
rect 34692 37884 37212 37940
rect 37268 37884 37772 37940
rect 37828 37884 37838 37940
rect 39218 37884 39228 37940
rect 39284 37884 40348 37940
rect 40404 37884 41132 37940
rect 41188 37884 41198 37940
rect 15810 37772 15820 37828
rect 15876 37772 16380 37828
rect 16436 37772 19180 37828
rect 19236 37772 19246 37828
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 2594 37436 2604 37492
rect 2660 37436 4620 37492
rect 4676 37436 4686 37492
rect 23874 37436 23884 37492
rect 23940 37436 25228 37492
rect 25284 37436 25294 37492
rect 4386 37212 4396 37268
rect 4452 37212 5628 37268
rect 5684 37212 5694 37268
rect 24546 36988 24556 37044
rect 24612 36988 25564 37044
rect 25620 36988 25630 37044
rect 37090 36988 37100 37044
rect 37156 36988 39340 37044
rect 39396 36988 40236 37044
rect 40292 36988 40302 37044
rect 25778 36876 25788 36932
rect 25844 36876 26684 36932
rect 26740 36876 27132 36932
rect 27188 36876 27198 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 4834 36652 4844 36708
rect 4900 36652 7420 36708
rect 7476 36652 7486 36708
rect 7746 36652 7756 36708
rect 7812 36652 9548 36708
rect 9604 36652 9614 36708
rect 6178 36428 6188 36484
rect 6244 36428 19740 36484
rect 19796 36428 20188 36484
rect 20244 36428 20254 36484
rect 21634 36428 21644 36484
rect 21700 36428 23436 36484
rect 23492 36428 23502 36484
rect 37090 36428 37100 36484
rect 37156 36428 37660 36484
rect 37716 36428 37726 36484
rect 6962 36316 6972 36372
rect 7028 36316 7980 36372
rect 8036 36316 15148 36372
rect 15204 36316 15214 36372
rect 18722 36316 18732 36372
rect 18788 36316 20524 36372
rect 20580 36316 23660 36372
rect 23716 36316 23726 36372
rect 20402 36204 20412 36260
rect 20468 36204 21868 36260
rect 21924 36204 21934 36260
rect 37986 36204 37996 36260
rect 38052 36204 40012 36260
rect 40068 36204 40078 36260
rect 40786 36204 40796 36260
rect 40852 36204 41132 36260
rect 41188 36204 43820 36260
rect 43876 36204 43886 36260
rect 40674 36092 40684 36148
rect 40740 36092 41020 36148
rect 41076 36092 41086 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 9874 35868 9884 35924
rect 9940 35868 10892 35924
rect 10948 35868 10958 35924
rect 36754 35644 36764 35700
rect 36820 35644 38108 35700
rect 38164 35644 38780 35700
rect 38836 35644 39452 35700
rect 39508 35644 40908 35700
rect 40964 35644 40974 35700
rect 8418 35532 8428 35588
rect 8484 35532 9660 35588
rect 9716 35532 9726 35588
rect 35970 35532 35980 35588
rect 36036 35532 37212 35588
rect 37268 35532 37278 35588
rect 37538 35532 37548 35588
rect 37604 35532 39788 35588
rect 39844 35532 39854 35588
rect 40226 35532 40236 35588
rect 40292 35532 41692 35588
rect 41748 35532 41758 35588
rect 5282 35420 5292 35476
rect 5348 35420 6972 35476
rect 7028 35420 7038 35476
rect 5170 35308 5180 35364
rect 5236 35308 8540 35364
rect 8596 35308 8606 35364
rect 21858 35308 21868 35364
rect 21924 35308 22988 35364
rect 23044 35308 23054 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 8866 35084 8876 35140
rect 8932 35084 20412 35140
rect 20468 35084 20478 35140
rect 33394 35084 33404 35140
rect 33460 35084 40348 35140
rect 40404 35084 40414 35140
rect 9314 34972 9324 35028
rect 9380 34972 11004 35028
rect 11060 34972 11070 35028
rect 7746 34860 7756 34916
rect 7812 34860 9772 34916
rect 9828 34860 9838 34916
rect 20178 34860 20188 34916
rect 20244 34860 24444 34916
rect 24500 34860 25228 34916
rect 25284 34860 25294 34916
rect 33842 34860 33852 34916
rect 33908 34860 35084 34916
rect 35140 34860 37100 34916
rect 37156 34860 37166 34916
rect 10098 34748 10108 34804
rect 10164 34748 11116 34804
rect 11172 34748 11676 34804
rect 11732 34748 11742 34804
rect 31266 34748 31276 34804
rect 31332 34748 32060 34804
rect 32116 34748 32126 34804
rect 9986 34636 9996 34692
rect 10052 34636 10332 34692
rect 10388 34636 10398 34692
rect 15810 34636 15820 34692
rect 15876 34636 16604 34692
rect 16660 34636 17164 34692
rect 17220 34636 18284 34692
rect 18340 34636 18350 34692
rect 18508 34636 20636 34692
rect 20692 34636 20702 34692
rect 24210 34636 24220 34692
rect 24276 34636 26012 34692
rect 26068 34636 26078 34692
rect 30594 34636 30604 34692
rect 30660 34636 33852 34692
rect 33908 34636 34636 34692
rect 34692 34636 34702 34692
rect 38210 34636 38220 34692
rect 38276 34636 40348 34692
rect 40404 34636 40414 34692
rect 18508 34580 18564 34636
rect 8754 34524 8764 34580
rect 8820 34524 9548 34580
rect 9604 34524 18564 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 7634 34300 7644 34356
rect 7700 34300 8540 34356
rect 8596 34300 8606 34356
rect 10546 34188 10556 34244
rect 10612 34188 12012 34244
rect 12068 34188 12078 34244
rect 22754 34188 22764 34244
rect 22820 34188 23324 34244
rect 23380 34188 25396 34244
rect 30818 34188 30828 34244
rect 30884 34188 33404 34244
rect 33460 34188 33470 34244
rect 25340 34132 25396 34188
rect 20626 34076 20636 34132
rect 20692 34076 23548 34132
rect 23604 34076 23614 34132
rect 25330 34076 25340 34132
rect 25396 34076 26796 34132
rect 26852 34076 26862 34132
rect 30146 34076 30156 34132
rect 30212 34076 30940 34132
rect 30996 34076 31006 34132
rect 31378 34076 31388 34132
rect 31444 34076 32284 34132
rect 32340 34076 32350 34132
rect 8866 33964 8876 34020
rect 8932 33964 9660 34020
rect 9716 33964 10220 34020
rect 10276 33964 10286 34020
rect 11330 33964 11340 34020
rect 11396 33964 12796 34020
rect 12852 33964 15932 34020
rect 15988 33964 16380 34020
rect 16436 33964 18508 34020
rect 18564 33964 18574 34020
rect 23874 33964 23884 34020
rect 23940 33964 25788 34020
rect 25844 33964 25854 34020
rect 29698 33964 29708 34020
rect 29764 33964 31164 34020
rect 31220 33964 31230 34020
rect 31826 33964 31836 34020
rect 31892 33964 32396 34020
rect 32452 33964 34524 34020
rect 34580 33964 34590 34020
rect 2930 33852 2940 33908
rect 2996 33852 6972 33908
rect 7028 33852 7038 33908
rect 23650 33852 23660 33908
rect 23716 33852 24892 33908
rect 24948 33852 25564 33908
rect 25620 33852 25630 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 12114 33628 12124 33684
rect 12180 33628 12460 33684
rect 12516 33628 12526 33684
rect 5730 33516 5740 33572
rect 5796 33516 12012 33572
rect 12068 33516 12078 33572
rect 21074 33516 21084 33572
rect 21140 33516 22204 33572
rect 22260 33516 22270 33572
rect 8372 33404 8540 33460
rect 8596 33404 20188 33460
rect 8372 33348 8428 33404
rect 20132 33348 20188 33404
rect 31892 33348 31948 33964
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 40450 33404 40460 33460
rect 40516 33404 43820 33460
rect 43876 33404 43886 33460
rect 7298 33292 7308 33348
rect 7364 33292 8204 33348
rect 8260 33292 8428 33348
rect 13794 33292 13804 33348
rect 13860 33292 15484 33348
rect 15540 33292 15820 33348
rect 15876 33292 15886 33348
rect 20132 33292 31948 33348
rect 40002 33292 40012 33348
rect 40068 33292 40908 33348
rect 40964 33292 40974 33348
rect 12450 33180 12460 33236
rect 12516 33180 15036 33236
rect 15092 33180 17276 33236
rect 17332 33180 17342 33236
rect 6626 33068 6636 33124
rect 6692 33068 7756 33124
rect 7812 33068 7822 33124
rect 13010 33068 13020 33124
rect 13076 33068 14700 33124
rect 14756 33068 15260 33124
rect 15316 33068 17052 33124
rect 17108 33068 17612 33124
rect 17668 33068 30156 33124
rect 30212 33068 30222 33124
rect 5058 32956 5068 33012
rect 5124 32956 5134 33012
rect 5068 32676 5124 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 20402 32844 20412 32900
rect 20468 32844 23100 32900
rect 23156 32844 23166 32900
rect 41010 32844 41020 32900
rect 41076 32844 41086 32900
rect 41020 32788 41076 32844
rect 12114 32732 12124 32788
rect 12180 32732 13020 32788
rect 13076 32732 13086 32788
rect 15474 32732 15484 32788
rect 15540 32732 16380 32788
rect 16436 32732 16446 32788
rect 20290 32732 20300 32788
rect 20356 32732 21084 32788
rect 21140 32732 21150 32788
rect 33730 32732 33740 32788
rect 33796 32732 34188 32788
rect 34244 32732 35756 32788
rect 35812 32732 35822 32788
rect 36306 32732 36316 32788
rect 36372 32732 41692 32788
rect 41748 32732 41758 32788
rect 5068 32620 7756 32676
rect 7812 32620 9772 32676
rect 9828 32620 9838 32676
rect 15810 32620 15820 32676
rect 15876 32620 16716 32676
rect 16772 32620 16782 32676
rect 16034 32508 16044 32564
rect 16100 32508 17836 32564
rect 17892 32508 17902 32564
rect 22194 32508 22204 32564
rect 22260 32508 24892 32564
rect 24948 32508 24958 32564
rect 3042 32396 3052 32452
rect 3108 32396 6972 32452
rect 7028 32396 7038 32452
rect 22642 32396 22652 32452
rect 22708 32396 25676 32452
rect 25732 32396 25742 32452
rect 15026 32284 15036 32340
rect 15092 32284 16268 32340
rect 16324 32284 16334 32340
rect 10434 32172 10444 32228
rect 10500 32172 11900 32228
rect 11956 32172 13580 32228
rect 13636 32172 19516 32228
rect 19572 32172 19582 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 6738 32060 6748 32116
rect 6804 32060 14588 32116
rect 14644 32060 14654 32116
rect 37202 31948 37212 32004
rect 37268 31948 37278 32004
rect 37212 31892 37268 31948
rect 6178 31836 6188 31892
rect 6244 31836 6860 31892
rect 6916 31836 8540 31892
rect 8596 31836 8606 31892
rect 19618 31836 19628 31892
rect 19684 31836 20076 31892
rect 20132 31836 20142 31892
rect 25778 31836 25788 31892
rect 25844 31836 26348 31892
rect 26404 31836 26414 31892
rect 37212 31836 38108 31892
rect 38164 31836 39564 31892
rect 39620 31836 40348 31892
rect 40404 31836 40414 31892
rect 8082 31724 8092 31780
rect 8148 31724 8988 31780
rect 9044 31724 9054 31780
rect 10770 31724 10780 31780
rect 10836 31724 11116 31780
rect 11172 31724 11182 31780
rect 15474 31724 15484 31780
rect 15540 31724 19852 31780
rect 19908 31724 19918 31780
rect 25218 31724 25228 31780
rect 25284 31724 26460 31780
rect 26516 31724 26526 31780
rect 30370 31724 30380 31780
rect 30436 31724 31388 31780
rect 31444 31724 31454 31780
rect 10658 31612 10668 31668
rect 10724 31612 11452 31668
rect 11508 31612 11518 31668
rect 19394 31612 19404 31668
rect 19460 31612 20412 31668
rect 20468 31612 20478 31668
rect 34066 31612 34076 31668
rect 34132 31612 34860 31668
rect 34916 31612 34926 31668
rect 37202 31612 37212 31668
rect 37268 31612 39340 31668
rect 39396 31612 39406 31668
rect 40562 31612 40572 31668
rect 40628 31612 41580 31668
rect 41636 31612 41646 31668
rect 9426 31500 9436 31556
rect 9492 31500 19068 31556
rect 19124 31500 19134 31556
rect 11106 31388 11116 31444
rect 11172 31388 12572 31444
rect 12628 31388 12638 31444
rect 25554 31388 25564 31444
rect 25620 31388 26124 31444
rect 26180 31388 26190 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 15026 31164 15036 31220
rect 15092 31164 19628 31220
rect 19684 31164 19694 31220
rect 34738 31164 34748 31220
rect 34804 31164 35532 31220
rect 35588 31164 35598 31220
rect 26572 31052 29036 31108
rect 29092 31052 29102 31108
rect 26572 30996 26628 31052
rect 16930 30940 16940 30996
rect 16996 30940 19292 30996
rect 19348 30940 19358 30996
rect 26002 30940 26012 30996
rect 26068 30940 26628 30996
rect 26898 30940 26908 30996
rect 26964 30940 30268 30996
rect 30324 30940 30334 30996
rect 34850 30940 34860 30996
rect 34916 30940 35756 30996
rect 35812 30940 35822 30996
rect 15810 30828 15820 30884
rect 15876 30828 16380 30884
rect 16436 30828 20636 30884
rect 20692 30828 26684 30884
rect 26740 30828 30492 30884
rect 30548 30828 30558 30884
rect 31266 30828 31276 30884
rect 31332 30828 35084 30884
rect 35140 30828 35150 30884
rect 30492 30772 30548 30828
rect 10210 30716 10220 30772
rect 10276 30716 11116 30772
rect 11172 30716 11182 30772
rect 25554 30716 25564 30772
rect 25620 30716 26460 30772
rect 26516 30716 26526 30772
rect 29586 30716 29596 30772
rect 29652 30716 29662 30772
rect 30492 30716 33964 30772
rect 34020 30716 34030 30772
rect 29596 30660 29652 30716
rect 6850 30604 6860 30660
rect 6916 30604 7420 30660
rect 7476 30604 7486 30660
rect 18946 30604 18956 30660
rect 19012 30604 29652 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 26450 30492 26460 30548
rect 26516 30492 26796 30548
rect 26852 30492 26862 30548
rect 17938 30268 17948 30324
rect 18004 30268 18620 30324
rect 18676 30268 18686 30324
rect 18834 30268 18844 30324
rect 18900 30268 19516 30324
rect 19572 30268 19582 30324
rect 6626 30156 6636 30212
rect 6692 30156 9212 30212
rect 9268 30156 9278 30212
rect 11218 30156 11228 30212
rect 11284 30156 11294 30212
rect 14578 30156 14588 30212
rect 14644 30156 16044 30212
rect 16100 30156 16110 30212
rect 30594 30156 30604 30212
rect 30660 30156 30670 30212
rect 31266 30156 31276 30212
rect 31332 30156 31948 30212
rect 32004 30156 32014 30212
rect 32386 30156 32396 30212
rect 32452 30156 36988 30212
rect 37044 30156 37054 30212
rect 11228 30100 11284 30156
rect 30604 30100 30660 30156
rect 7074 30044 7084 30100
rect 7140 30044 11284 30100
rect 11554 30044 11564 30100
rect 11620 30044 12124 30100
rect 12180 30044 12190 30100
rect 14690 30044 14700 30100
rect 14756 30044 15596 30100
rect 15652 30044 15662 30100
rect 25890 30044 25900 30100
rect 25956 30044 27356 30100
rect 27412 30044 27422 30100
rect 30604 30044 32060 30100
rect 32116 30044 37100 30100
rect 37156 30044 37884 30100
rect 37940 30044 37950 30100
rect 11666 29932 11676 29988
rect 11732 29932 16492 29988
rect 16548 29932 16558 29988
rect 25778 29932 25788 29988
rect 25844 29932 27244 29988
rect 27300 29932 29708 29988
rect 29764 29932 29774 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 16258 29708 16268 29764
rect 16324 29708 16716 29764
rect 16772 29708 16782 29764
rect 41682 29708 41692 29764
rect 41748 29708 42476 29764
rect 42532 29708 42542 29764
rect 10098 29484 10108 29540
rect 10164 29484 11172 29540
rect 14578 29484 14588 29540
rect 14644 29484 15148 29540
rect 15204 29484 15214 29540
rect 29810 29484 29820 29540
rect 29876 29484 31276 29540
rect 31332 29484 31342 29540
rect 33618 29484 33628 29540
rect 33684 29484 39788 29540
rect 39844 29484 39854 29540
rect 11116 29428 11172 29484
rect 4722 29372 4732 29428
rect 4788 29372 5964 29428
rect 6020 29372 6636 29428
rect 6692 29372 6702 29428
rect 9426 29372 9436 29428
rect 9492 29372 10220 29428
rect 10276 29372 10286 29428
rect 11106 29372 11116 29428
rect 11172 29372 11676 29428
rect 11732 29372 25564 29428
rect 25620 29372 31052 29428
rect 31108 29372 31500 29428
rect 31556 29372 33292 29428
rect 33348 29372 33358 29428
rect 38546 29372 38556 29428
rect 38612 29372 40348 29428
rect 40404 29372 40414 29428
rect 6402 29260 6412 29316
rect 6468 29260 7420 29316
rect 7476 29260 7486 29316
rect 20402 29260 20412 29316
rect 20468 29260 24668 29316
rect 24724 29260 24734 29316
rect 42578 29260 42588 29316
rect 42644 29260 43820 29316
rect 43876 29260 43886 29316
rect 27346 29036 27356 29092
rect 27412 29036 30380 29092
rect 30436 29036 30446 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 6738 28812 6748 28868
rect 6804 28812 7756 28868
rect 7812 28812 9772 28868
rect 9828 28812 9838 28868
rect 12114 28812 12124 28868
rect 12180 28812 16716 28868
rect 16772 28812 16782 28868
rect 9314 28700 9324 28756
rect 9380 28700 13468 28756
rect 13524 28700 13534 28756
rect 14354 28700 14364 28756
rect 14420 28700 16156 28756
rect 16212 28700 16222 28756
rect 18274 28700 18284 28756
rect 18340 28700 19404 28756
rect 19460 28700 19470 28756
rect 37538 28700 37548 28756
rect 37604 28700 39004 28756
rect 39060 28700 41468 28756
rect 41524 28700 41534 28756
rect 8754 28588 8764 28644
rect 8820 28588 10108 28644
rect 10164 28588 10174 28644
rect 10770 28588 10780 28644
rect 10836 28588 15484 28644
rect 15540 28588 15550 28644
rect 37090 28588 37100 28644
rect 37156 28588 37772 28644
rect 37828 28588 37838 28644
rect 15810 28476 15820 28532
rect 15876 28476 21308 28532
rect 21364 28476 21374 28532
rect 40562 28476 40572 28532
rect 40628 28476 42364 28532
rect 42420 28476 42430 28532
rect 36082 28364 36092 28420
rect 36148 28364 37996 28420
rect 38052 28364 38062 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 12898 28028 12908 28084
rect 12964 28028 14924 28084
rect 14980 28028 14990 28084
rect 9986 27916 9996 27972
rect 10052 27916 13692 27972
rect 13748 27916 13758 27972
rect 15362 27916 15372 27972
rect 15428 27916 16156 27972
rect 16212 27916 16222 27972
rect 18498 27916 18508 27972
rect 18564 27916 19292 27972
rect 19348 27916 19358 27972
rect 14914 27804 14924 27860
rect 14980 27804 15260 27860
rect 15316 27804 15820 27860
rect 15876 27804 15886 27860
rect 16034 27804 16044 27860
rect 16100 27804 16380 27860
rect 16436 27804 16446 27860
rect 13234 27692 13244 27748
rect 13300 27692 14028 27748
rect 14084 27692 14094 27748
rect 18946 27692 18956 27748
rect 19012 27692 20524 27748
rect 20580 27692 20590 27748
rect 31826 27692 31836 27748
rect 31892 27692 34860 27748
rect 34916 27692 35756 27748
rect 35812 27692 35822 27748
rect 38658 27692 38668 27748
rect 38724 27692 39340 27748
rect 39396 27692 39406 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 30706 27244 30716 27300
rect 30772 27244 31836 27300
rect 31892 27244 31902 27300
rect 19730 27132 19740 27188
rect 19796 27132 25228 27188
rect 25284 27132 25294 27188
rect 17826 27020 17836 27076
rect 17892 27020 21756 27076
rect 21812 27020 22652 27076
rect 22708 27020 22718 27076
rect 25890 27020 25900 27076
rect 25956 27020 34412 27076
rect 34468 27020 34478 27076
rect 35746 27020 35756 27076
rect 35812 27020 37436 27076
rect 37492 27020 37502 27076
rect 2594 26908 2604 26964
rect 2660 26908 3724 26964
rect 3780 26908 3790 26964
rect 12898 26908 12908 26964
rect 12964 26908 13748 26964
rect 27010 26908 27020 26964
rect 27076 26908 30044 26964
rect 30100 26908 34076 26964
rect 34132 26908 34142 26964
rect 13692 26740 13748 26908
rect 14130 26796 14140 26852
rect 14196 26796 15372 26852
rect 15428 26796 15438 26852
rect 22978 26796 22988 26852
rect 23044 26796 25228 26852
rect 25284 26796 25564 26852
rect 25620 26796 25630 26852
rect 13682 26684 13692 26740
rect 13748 26684 13758 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 15586 26572 15596 26628
rect 15652 26572 17276 26628
rect 17332 26572 17342 26628
rect 10994 26460 11004 26516
rect 11060 26460 11788 26516
rect 11844 26460 12348 26516
rect 12404 26460 12414 26516
rect 16258 26460 16268 26516
rect 16324 26460 17388 26516
rect 17444 26460 17454 26516
rect 35634 26460 35644 26516
rect 35700 26460 36428 26516
rect 36484 26460 36494 26516
rect 16818 26348 16828 26404
rect 16884 26348 17948 26404
rect 18004 26348 18732 26404
rect 18788 26348 19628 26404
rect 19684 26348 30044 26404
rect 30100 26348 31612 26404
rect 31668 26348 31678 26404
rect 6738 26236 6748 26292
rect 6804 26236 7084 26292
rect 7140 26236 12684 26292
rect 12740 26236 16604 26292
rect 16660 26236 18956 26292
rect 19012 26236 19022 26292
rect 29810 26236 29820 26292
rect 29876 26236 30716 26292
rect 30772 26236 30782 26292
rect 31266 26236 31276 26292
rect 31332 26236 31948 26292
rect 32004 26236 32014 26292
rect 2594 26124 2604 26180
rect 2660 26124 4060 26180
rect 4116 26124 4126 26180
rect 4722 26124 4732 26180
rect 4788 26124 5964 26180
rect 6020 26124 6030 26180
rect 6626 26124 6636 26180
rect 6692 26124 7308 26180
rect 7364 26124 7374 26180
rect 23762 26124 23772 26180
rect 23828 26124 24892 26180
rect 24948 26124 24958 26180
rect 29474 26124 29484 26180
rect 29540 26124 30268 26180
rect 30324 26124 30334 26180
rect 11218 25900 11228 25956
rect 11284 25900 12012 25956
rect 12068 25900 13132 25956
rect 13188 25900 32396 25956
rect 32452 25900 34860 25956
rect 34916 25900 34926 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 8418 25788 8428 25844
rect 8484 25788 23772 25844
rect 23828 25788 23838 25844
rect 4386 25564 4396 25620
rect 4452 25564 5852 25620
rect 5908 25564 5918 25620
rect 37874 25564 37884 25620
rect 37940 25564 37950 25620
rect 38210 25564 38220 25620
rect 38276 25564 38668 25620
rect 38724 25564 40236 25620
rect 40292 25564 41132 25620
rect 41188 25564 41198 25620
rect 43652 25564 44044 25620
rect 44100 25564 44110 25620
rect 37884 25508 37940 25564
rect 43652 25508 43708 25564
rect 37884 25452 40684 25508
rect 40740 25452 43708 25508
rect 6514 25340 6524 25396
rect 6580 25340 6748 25396
rect 6804 25340 6814 25396
rect 16706 25340 16716 25396
rect 16772 25340 17276 25396
rect 17332 25340 18060 25396
rect 18116 25340 18126 25396
rect 7298 25228 7308 25284
rect 7364 25228 7756 25284
rect 7812 25228 8764 25284
rect 8820 25228 8830 25284
rect 11218 25228 11228 25284
rect 11284 25228 11452 25284
rect 11508 25228 11518 25284
rect 31602 25228 31612 25284
rect 31668 25228 35644 25284
rect 35700 25228 35710 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 27682 24892 27692 24948
rect 27748 24892 29260 24948
rect 29316 24892 29326 24948
rect 35522 24892 35532 24948
rect 35588 24892 36540 24948
rect 36596 24892 39788 24948
rect 39844 24892 39854 24948
rect 28690 24780 28700 24836
rect 28756 24780 29932 24836
rect 29988 24780 33852 24836
rect 33908 24780 33918 24836
rect 40002 24780 40012 24836
rect 40068 24780 42364 24836
rect 42420 24780 42430 24836
rect 5394 24668 5404 24724
rect 5460 24668 6076 24724
rect 6132 24668 6142 24724
rect 28578 24668 28588 24724
rect 28644 24668 29596 24724
rect 29652 24668 29662 24724
rect 39218 24668 39228 24724
rect 39284 24668 41804 24724
rect 41860 24668 41870 24724
rect 4050 24556 4060 24612
rect 4116 24556 6300 24612
rect 6356 24556 6366 24612
rect 13570 24332 13580 24388
rect 13636 24332 14252 24388
rect 14308 24332 18396 24388
rect 18452 24332 18462 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 39890 24108 39900 24164
rect 39956 24108 42028 24164
rect 42084 24108 42094 24164
rect 9426 23996 9436 24052
rect 9492 23996 10892 24052
rect 10948 23996 11228 24052
rect 11284 23996 16268 24052
rect 16324 23996 16334 24052
rect 9090 23884 9100 23940
rect 9156 23884 10780 23940
rect 10836 23884 11508 23940
rect 15698 23884 15708 23940
rect 15764 23884 16492 23940
rect 16548 23884 17276 23940
rect 17332 23884 17342 23940
rect 11452 23828 11508 23884
rect 11442 23772 11452 23828
rect 11508 23772 11518 23828
rect 19170 23772 19180 23828
rect 19236 23772 20412 23828
rect 20468 23772 20478 23828
rect 21746 23772 21756 23828
rect 21812 23772 23548 23828
rect 23604 23772 23614 23828
rect 6178 23660 6188 23716
rect 6244 23660 8876 23716
rect 8932 23660 9660 23716
rect 9716 23660 9726 23716
rect 36082 23660 36092 23716
rect 36148 23660 36540 23716
rect 36596 23660 36606 23716
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 16930 23436 16940 23492
rect 16996 23436 17724 23492
rect 17780 23436 18396 23492
rect 18452 23436 18462 23492
rect 36194 23436 36204 23492
rect 36260 23436 38668 23492
rect 6066 23324 6076 23380
rect 6132 23324 8204 23380
rect 8260 23324 11228 23380
rect 11284 23324 11294 23380
rect 11442 23324 11452 23380
rect 11508 23324 12012 23380
rect 12068 23324 12078 23380
rect 12338 23324 12348 23380
rect 12404 23324 12684 23380
rect 12740 23324 13356 23380
rect 13412 23324 13422 23380
rect 16034 23324 16044 23380
rect 16100 23324 17388 23380
rect 17444 23324 17454 23380
rect 31714 23324 31724 23380
rect 31780 23324 32396 23380
rect 32452 23324 32462 23380
rect 12348 23156 12404 23324
rect 17490 23212 17500 23268
rect 17556 23212 19236 23268
rect 25778 23212 25788 23268
rect 25844 23212 35308 23268
rect 35364 23212 35374 23268
rect 19180 23156 19236 23212
rect 38612 23156 38668 23436
rect 9202 23100 9212 23156
rect 9268 23100 9884 23156
rect 9940 23100 9950 23156
rect 11218 23100 11228 23156
rect 11284 23100 12404 23156
rect 17714 23100 17724 23156
rect 17780 23100 18396 23156
rect 18452 23100 18462 23156
rect 19170 23100 19180 23156
rect 19236 23100 19740 23156
rect 19796 23100 19806 23156
rect 28242 23100 28252 23156
rect 28308 23100 30380 23156
rect 30436 23100 30446 23156
rect 35634 23100 35644 23156
rect 35700 23100 37212 23156
rect 37268 23100 37278 23156
rect 38612 23100 39676 23156
rect 39732 23100 39742 23156
rect 6962 22988 6972 23044
rect 7028 22988 7980 23044
rect 8036 22988 13692 23044
rect 13748 22988 13758 23044
rect 31714 22876 31724 22932
rect 31780 22876 32284 22932
rect 32340 22876 39004 22932
rect 39060 22876 39070 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 35410 22540 35420 22596
rect 35476 22540 36092 22596
rect 36148 22540 36158 22596
rect 4162 22428 4172 22484
rect 4228 22428 5740 22484
rect 5796 22428 5806 22484
rect 6178 22428 6188 22484
rect 6244 22428 8428 22484
rect 8484 22428 8494 22484
rect 19842 22428 19852 22484
rect 19908 22428 21420 22484
rect 21476 22428 21486 22484
rect 25666 22428 25676 22484
rect 25732 22428 26684 22484
rect 26740 22428 26750 22484
rect 1698 22316 1708 22372
rect 1764 22316 21980 22372
rect 22036 22316 22046 22372
rect 33618 22316 33628 22372
rect 33684 22316 36764 22372
rect 36820 22316 37100 22372
rect 37156 22316 37166 22372
rect 6290 22204 6300 22260
rect 6356 22204 10220 22260
rect 10276 22204 10286 22260
rect 2594 22092 2604 22148
rect 2660 22092 4060 22148
rect 4116 22092 4126 22148
rect 4834 22092 4844 22148
rect 4900 22092 5852 22148
rect 5908 22092 9884 22148
rect 9940 22092 9950 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 13682 21868 13692 21924
rect 13748 21868 14588 21924
rect 14644 21868 14654 21924
rect 17490 21756 17500 21812
rect 17556 21756 18396 21812
rect 18452 21756 18462 21812
rect 34290 21756 34300 21812
rect 34356 21756 35308 21812
rect 35364 21756 35374 21812
rect 11442 21532 11452 21588
rect 11508 21532 15260 21588
rect 15316 21532 19628 21588
rect 19684 21532 19694 21588
rect 24210 21532 24220 21588
rect 24276 21532 24780 21588
rect 24836 21532 25452 21588
rect 25508 21532 28756 21588
rect 28700 21476 28756 21532
rect 14690 21420 14700 21476
rect 14756 21420 15596 21476
rect 15652 21420 15662 21476
rect 26114 21420 26124 21476
rect 26180 21420 27020 21476
rect 27076 21420 27086 21476
rect 28690 21420 28700 21476
rect 28756 21420 29596 21476
rect 29652 21420 33180 21476
rect 33236 21420 33246 21476
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 18834 20860 18844 20916
rect 18900 20860 19628 20916
rect 19684 20860 19852 20916
rect 19908 20860 19918 20916
rect 9090 20748 9100 20804
rect 9156 20748 24444 20804
rect 24500 20748 26684 20804
rect 26740 20748 29820 20804
rect 29876 20748 29886 20804
rect 18274 20636 18284 20692
rect 18340 20636 19180 20692
rect 19236 20636 19246 20692
rect 3826 20524 3836 20580
rect 3892 20524 10668 20580
rect 10724 20524 13804 20580
rect 13860 20524 14476 20580
rect 14532 20524 14542 20580
rect 19618 20524 19628 20580
rect 19684 20524 19740 20580
rect 19796 20524 19806 20580
rect 25442 20412 25452 20468
rect 25508 20412 25788 20468
rect 25844 20412 39116 20468
rect 39172 20412 39182 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 19170 20300 19180 20356
rect 19236 20300 19628 20356
rect 19684 20300 19694 20356
rect 3332 20188 5348 20244
rect 16034 20188 16044 20244
rect 16100 20188 19404 20244
rect 19460 20188 19470 20244
rect 19618 20188 19628 20244
rect 19684 20188 19740 20244
rect 19796 20188 19806 20244
rect 23986 20188 23996 20244
rect 24052 20188 24556 20244
rect 24612 20188 24780 20244
rect 24836 20188 25116 20244
rect 25172 20188 25182 20244
rect 3332 20020 3388 20188
rect 1922 19964 1932 20020
rect 1988 19964 3388 20020
rect 5292 19908 5348 20188
rect 10882 20076 10892 20132
rect 10948 20076 18844 20132
rect 18900 20076 18910 20132
rect 22978 20076 22988 20132
rect 23044 20076 23660 20132
rect 23716 20076 23726 20132
rect 39554 20076 39564 20132
rect 39620 20076 40572 20132
rect 40628 20076 41748 20132
rect 41692 20020 41748 20076
rect 13682 19964 13692 20020
rect 13748 19964 17612 20020
rect 17668 19964 18508 20020
rect 18564 19964 18574 20020
rect 41682 19964 41692 20020
rect 41748 19964 41758 20020
rect 5282 19852 5292 19908
rect 5348 19852 9884 19908
rect 9940 19852 13580 19908
rect 13636 19852 13646 19908
rect 19618 19852 19628 19908
rect 19684 19852 20636 19908
rect 20692 19852 20702 19908
rect 41794 19852 41804 19908
rect 41860 19852 42364 19908
rect 42420 19852 44044 19908
rect 44100 19852 44110 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41682 19180 41692 19236
rect 41748 19180 42476 19236
rect 42532 19180 42542 19236
rect 31938 19068 31948 19124
rect 32004 19068 38892 19124
rect 38948 19068 38958 19124
rect 39890 19068 39900 19124
rect 39956 19068 41132 19124
rect 41188 19068 41198 19124
rect 6850 18956 6860 19012
rect 6916 18956 6926 19012
rect 35634 18956 35644 19012
rect 35700 18956 36092 19012
rect 36148 18956 36158 19012
rect 6860 18900 6916 18956
rect 6860 18844 7084 18900
rect 7140 18844 7150 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 5506 18508 5516 18564
rect 5572 18508 6524 18564
rect 6580 18508 7140 18564
rect 14130 18508 14140 18564
rect 14196 18508 22988 18564
rect 23044 18508 23054 18564
rect 35746 18508 35756 18564
rect 35812 18508 41020 18564
rect 41076 18508 41086 18564
rect 7084 18452 7140 18508
rect 4946 18396 4956 18452
rect 5012 18396 6860 18452
rect 6916 18396 6926 18452
rect 7084 18396 9548 18452
rect 9604 18396 9614 18452
rect 9874 18396 9884 18452
rect 9940 18396 11228 18452
rect 11284 18396 11294 18452
rect 11890 18396 11900 18452
rect 11956 18396 12348 18452
rect 12404 18396 13468 18452
rect 13524 18396 13534 18452
rect 20962 18396 20972 18452
rect 21028 18396 22428 18452
rect 22484 18396 22494 18452
rect 36418 18396 36428 18452
rect 36484 18396 41580 18452
rect 41636 18396 43372 18452
rect 43428 18396 43438 18452
rect 5842 18284 5852 18340
rect 5908 18284 6748 18340
rect 6804 18284 6814 18340
rect 30034 18284 30044 18340
rect 30100 18284 31276 18340
rect 31332 18284 31342 18340
rect 2594 18172 2604 18228
rect 2660 18172 4956 18228
rect 5012 18172 5022 18228
rect 6402 18172 6412 18228
rect 6468 18172 7980 18228
rect 8036 18172 8046 18228
rect 6626 18060 6636 18116
rect 6692 18060 7756 18116
rect 7812 18060 7822 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 5954 17724 5964 17780
rect 6020 17724 7084 17780
rect 7140 17724 7980 17780
rect 8036 17724 8046 17780
rect 18610 17724 18620 17780
rect 18676 17724 19180 17780
rect 19236 17724 25900 17780
rect 25956 17724 29484 17780
rect 29540 17724 29550 17780
rect 35308 17724 36428 17780
rect 36484 17724 36494 17780
rect 35308 17668 35364 17724
rect 4722 17612 4732 17668
rect 4788 17612 5740 17668
rect 5796 17612 5806 17668
rect 25666 17612 25676 17668
rect 25732 17612 28644 17668
rect 33842 17612 33852 17668
rect 33908 17612 35308 17668
rect 35364 17612 35374 17668
rect 35858 17612 35868 17668
rect 35924 17612 37324 17668
rect 37380 17612 37390 17668
rect 23986 17500 23996 17556
rect 24052 17500 25228 17556
rect 25284 17500 25294 17556
rect 28588 17444 28644 17612
rect 35970 17500 35980 17556
rect 36036 17500 36540 17556
rect 36596 17500 36988 17556
rect 37044 17500 37054 17556
rect 6738 17388 6748 17444
rect 6804 17388 7420 17444
rect 7476 17388 7486 17444
rect 14802 17388 14812 17444
rect 14868 17388 15708 17444
rect 15764 17388 17948 17444
rect 18004 17388 18014 17444
rect 23650 17388 23660 17444
rect 23716 17388 24556 17444
rect 24612 17388 27804 17444
rect 27860 17388 27870 17444
rect 28578 17388 28588 17444
rect 28644 17388 30156 17444
rect 30212 17388 30222 17444
rect 37202 17388 37212 17444
rect 37268 17388 40460 17444
rect 40516 17388 40526 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 17948 17164 18284 17220
rect 18340 17164 18350 17220
rect 17948 16884 18004 17164
rect 19282 17052 19292 17108
rect 19348 17052 19740 17108
rect 19796 17052 20636 17108
rect 20692 17052 20702 17108
rect 29932 17052 31948 17108
rect 32004 17052 32014 17108
rect 24098 16940 24108 16996
rect 24164 16940 27692 16996
rect 27748 16940 27758 16996
rect 29932 16884 29988 17052
rect 32050 16940 32060 16996
rect 32116 16940 32508 16996
rect 32564 16940 33628 16996
rect 33684 16940 36764 16996
rect 36820 16940 36830 16996
rect 11666 16828 11676 16884
rect 11732 16828 15484 16884
rect 15540 16828 16604 16884
rect 16660 16828 16670 16884
rect 17938 16828 17948 16884
rect 18004 16828 18014 16884
rect 20178 16828 20188 16884
rect 20244 16828 20972 16884
rect 21028 16828 26572 16884
rect 26628 16828 29988 16884
rect 30146 16828 30156 16884
rect 30212 16828 33292 16884
rect 33348 16828 33358 16884
rect 16604 16772 16660 16828
rect 16604 16716 21420 16772
rect 21476 16716 25676 16772
rect 25732 16716 25742 16772
rect 27346 16716 27356 16772
rect 27412 16716 28364 16772
rect 28420 16716 28430 16772
rect 15922 16604 15932 16660
rect 15988 16604 17388 16660
rect 17444 16604 17454 16660
rect 21634 16604 21644 16660
rect 21700 16604 22540 16660
rect 22596 16604 23772 16660
rect 23828 16604 23838 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 8194 16156 8204 16212
rect 8260 16156 9100 16212
rect 9156 16156 9166 16212
rect 7858 16044 7868 16100
rect 7924 16044 9660 16100
rect 9716 16044 9726 16100
rect 13010 16044 13020 16100
rect 13076 16044 17836 16100
rect 17892 16044 17902 16100
rect 26852 15988 26908 16100
rect 26964 16044 26974 16100
rect 28354 16044 28364 16100
rect 28420 16044 29148 16100
rect 29204 16044 29214 16100
rect 7746 15932 7756 15988
rect 7812 15932 8540 15988
rect 8596 15932 8606 15988
rect 25218 15932 25228 15988
rect 25284 15932 26908 15988
rect 2706 15820 2716 15876
rect 2772 15820 7532 15876
rect 7588 15820 7598 15876
rect 14354 15820 14364 15876
rect 14420 15820 16044 15876
rect 16100 15820 19740 15876
rect 19796 15820 19806 15876
rect 25554 15820 25564 15876
rect 25620 15820 26796 15876
rect 26852 15820 29372 15876
rect 29428 15820 29438 15876
rect 37090 15820 37100 15876
rect 37156 15820 40124 15876
rect 40180 15820 40460 15876
rect 40516 15820 40526 15876
rect 4834 15708 4844 15764
rect 4900 15708 12460 15764
rect 12516 15708 12526 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 8866 15484 8876 15540
rect 8932 15484 13244 15540
rect 13300 15484 13310 15540
rect 29474 15484 29484 15540
rect 29540 15484 30604 15540
rect 30660 15484 30670 15540
rect 4834 15372 4844 15428
rect 4900 15372 6860 15428
rect 6916 15372 8652 15428
rect 8708 15372 9884 15428
rect 9940 15372 9950 15428
rect 14018 15372 14028 15428
rect 14084 15372 14094 15428
rect 7298 15260 7308 15316
rect 7364 15260 7980 15316
rect 8036 15260 8046 15316
rect 9538 15260 9548 15316
rect 9604 15260 10220 15316
rect 10276 15260 10286 15316
rect 12450 15260 12460 15316
rect 12516 15260 13132 15316
rect 13188 15260 13198 15316
rect 14028 15204 14084 15372
rect 29250 15260 29260 15316
rect 29316 15260 30380 15316
rect 30436 15260 30446 15316
rect 29820 15204 29876 15260
rect 8754 15148 8764 15204
rect 8820 15148 9436 15204
rect 9492 15148 14084 15204
rect 20626 15148 20636 15204
rect 20692 15148 21756 15204
rect 21812 15148 21822 15204
rect 29810 15148 29820 15204
rect 29876 15148 29886 15204
rect 25330 15036 25340 15092
rect 25396 15036 26012 15092
rect 26068 15036 26078 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 15250 14588 15260 14644
rect 15316 14588 16716 14644
rect 16772 14588 18508 14644
rect 18564 14588 19516 14644
rect 19572 14588 19582 14644
rect 6850 14364 6860 14420
rect 6916 14364 7756 14420
rect 7812 14364 9660 14420
rect 9716 14364 9726 14420
rect 9986 14252 9996 14308
rect 10052 14252 12796 14308
rect 12852 14252 13804 14308
rect 13860 14252 13870 14308
rect 36418 14252 36428 14308
rect 36484 14252 37324 14308
rect 37380 14252 37390 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 22082 13580 22092 13636
rect 22148 13580 22764 13636
rect 22820 13580 24332 13636
rect 24388 13580 25452 13636
rect 25508 13580 25518 13636
rect 24658 13468 24668 13524
rect 24724 13468 25564 13524
rect 25620 13468 25630 13524
rect 30818 13468 30828 13524
rect 30884 13468 32284 13524
rect 32340 13468 32350 13524
rect 13458 13356 13468 13412
rect 13524 13356 14252 13412
rect 14308 13356 14318 13412
rect 19842 13356 19852 13412
rect 19908 13356 20524 13412
rect 20580 13356 20590 13412
rect 25330 13356 25340 13412
rect 25396 13356 26124 13412
rect 26180 13356 29484 13412
rect 29540 13356 29550 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 6066 13020 6076 13076
rect 6132 13020 7644 13076
rect 7700 13020 7710 13076
rect 22866 13020 22876 13076
rect 22932 13020 24780 13076
rect 24836 13020 24846 13076
rect 29698 12908 29708 12964
rect 29764 12908 30380 12964
rect 30436 12908 30446 12964
rect 32946 12908 32956 12964
rect 33012 12908 33964 12964
rect 34020 12908 34030 12964
rect 6290 12796 6300 12852
rect 6356 12796 7756 12852
rect 7812 12796 8764 12852
rect 8820 12796 8830 12852
rect 30258 12796 30268 12852
rect 30324 12796 31948 12852
rect 32004 12796 32844 12852
rect 32900 12796 32910 12852
rect 8530 12684 8540 12740
rect 8596 12684 11564 12740
rect 11620 12684 11630 12740
rect 33058 12684 33068 12740
rect 33124 12684 35196 12740
rect 35252 12684 35262 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 8418 12348 8428 12404
rect 8484 12348 9660 12404
rect 9716 12348 9726 12404
rect 30594 12348 30604 12404
rect 30660 12348 32060 12404
rect 32116 12348 33068 12404
rect 33124 12348 33740 12404
rect 33796 12348 33806 12404
rect 2594 12236 2604 12292
rect 2660 12236 7644 12292
rect 7700 12236 7710 12292
rect 12226 12236 12236 12292
rect 12292 12236 12796 12292
rect 12852 12236 13468 12292
rect 13524 12236 13534 12292
rect 4722 12124 4732 12180
rect 4788 12124 6076 12180
rect 6132 12124 6142 12180
rect 7858 12124 7868 12180
rect 7924 12124 8652 12180
rect 8708 12124 8718 12180
rect 26226 12124 26236 12180
rect 26292 12124 26908 12180
rect 26964 12124 28140 12180
rect 28196 12124 31388 12180
rect 31444 12124 31454 12180
rect 9090 12012 9100 12068
rect 9156 12012 14812 12068
rect 14868 12012 14878 12068
rect 17938 12012 17948 12068
rect 18004 12012 19852 12068
rect 19908 12012 19918 12068
rect 32386 12012 32396 12068
rect 32452 12012 35868 12068
rect 35924 12012 36428 12068
rect 36484 12012 36494 12068
rect 13794 11900 13804 11956
rect 13860 11900 15036 11956
rect 15092 11900 15102 11956
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 15250 11676 15260 11732
rect 15316 11676 16044 11732
rect 16100 11676 17836 11732
rect 17892 11676 18284 11732
rect 18340 11676 18350 11732
rect 8866 11452 8876 11508
rect 8932 11452 9324 11508
rect 9380 11452 9390 11508
rect 11330 11340 11340 11396
rect 11396 11340 12236 11396
rect 12292 11340 12302 11396
rect 15698 11340 15708 11396
rect 15764 11340 17388 11396
rect 17444 11340 17454 11396
rect 17602 11340 17612 11396
rect 17668 11340 25340 11396
rect 25396 11340 25406 11396
rect 32498 11340 32508 11396
rect 32564 11340 33516 11396
rect 33572 11340 34748 11396
rect 34804 11340 34814 11396
rect 7186 11228 7196 11284
rect 7252 11228 8876 11284
rect 8932 11228 8942 11284
rect 11778 11228 11788 11284
rect 11844 11228 12348 11284
rect 12404 11228 13468 11284
rect 13524 11228 13692 11284
rect 13748 11228 13758 11284
rect 16706 11228 16716 11284
rect 16772 11228 17724 11284
rect 17780 11228 17790 11284
rect 18050 11228 18060 11284
rect 18116 11228 18620 11284
rect 18676 11228 18686 11284
rect 25778 11228 25788 11284
rect 25844 11228 27020 11284
rect 27076 11228 27086 11284
rect 30482 11228 30492 11284
rect 30548 11228 32060 11284
rect 32116 11228 33068 11284
rect 33124 11228 33134 11284
rect 6514 11116 6524 11172
rect 6580 11116 7532 11172
rect 7588 11116 7598 11172
rect 7858 11116 7868 11172
rect 7924 11116 8316 11172
rect 8372 11116 10220 11172
rect 10276 11116 10286 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 7634 10892 7644 10948
rect 7700 10892 8092 10948
rect 8148 10892 8158 10948
rect 14018 10780 14028 10836
rect 14084 10780 14094 10836
rect 14028 10724 14084 10780
rect 12674 10668 12684 10724
rect 12740 10668 15932 10724
rect 15988 10668 15998 10724
rect 29586 10668 29596 10724
rect 29652 10668 30380 10724
rect 30436 10668 31948 10724
rect 32004 10668 32014 10724
rect 7186 10556 7196 10612
rect 7252 10556 8092 10612
rect 8148 10556 8158 10612
rect 11218 10556 11228 10612
rect 11284 10556 11676 10612
rect 11732 10556 11742 10612
rect 12226 10556 12236 10612
rect 12292 10556 13804 10612
rect 13860 10556 13870 10612
rect 15250 10556 15260 10612
rect 15316 10556 16604 10612
rect 16660 10556 16670 10612
rect 28914 10556 28924 10612
rect 28980 10556 30044 10612
rect 30100 10556 30110 10612
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 10770 9996 10780 10052
rect 10836 9996 11564 10052
rect 11620 9996 12124 10052
rect 12180 9996 12190 10052
rect 12450 9996 12460 10052
rect 12516 9996 12908 10052
rect 12964 9996 14364 10052
rect 14420 9996 14430 10052
rect 15810 9996 15820 10052
rect 15876 9996 19068 10052
rect 19124 9996 19134 10052
rect 8082 9884 8092 9940
rect 8148 9884 23212 9940
rect 23268 9884 24108 9940
rect 24164 9884 24174 9940
rect 6738 9772 6748 9828
rect 6804 9772 7308 9828
rect 7364 9772 7980 9828
rect 8036 9772 8046 9828
rect 27458 9772 27468 9828
rect 27524 9772 29372 9828
rect 29428 9772 29438 9828
rect 17378 9660 17388 9716
rect 17444 9660 18172 9716
rect 18228 9660 18844 9716
rect 18900 9660 18910 9716
rect 4498 9548 4508 9604
rect 4564 9548 6636 9604
rect 6692 9548 6702 9604
rect 12786 9548 12796 9604
rect 12852 9548 13692 9604
rect 13748 9548 14588 9604
rect 14644 9548 14654 9604
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 20300 9324 26348 9380
rect 26404 9324 26414 9380
rect 20300 9268 20356 9324
rect 19618 9212 19628 9268
rect 19684 9212 20356 9268
rect 20514 9212 20524 9268
rect 20580 9212 21420 9268
rect 21476 9212 21868 9268
rect 21924 9212 21934 9268
rect 16482 9100 16492 9156
rect 16548 9100 17388 9156
rect 17444 9100 17454 9156
rect 23426 9100 23436 9156
rect 23492 9100 25340 9156
rect 25396 9100 27580 9156
rect 27636 9100 28364 9156
rect 28420 9100 28430 9156
rect 3826 8988 3836 9044
rect 3892 8988 5180 9044
rect 5236 8988 7084 9044
rect 7140 8988 7150 9044
rect 24658 8988 24668 9044
rect 24724 8988 25676 9044
rect 25732 8988 28700 9044
rect 28756 8988 28766 9044
rect 22978 8652 22988 8708
rect 23044 8652 23660 8708
rect 23716 8652 27132 8708
rect 27188 8652 27580 8708
rect 27636 8652 27646 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 26338 8428 26348 8484
rect 26404 8428 34972 8484
rect 35028 8428 35038 8484
rect 10882 8316 10892 8372
rect 10948 8316 11564 8372
rect 11620 8316 12572 8372
rect 12628 8316 12638 8372
rect 28242 8316 28252 8372
rect 28308 8316 29484 8372
rect 29540 8316 29550 8372
rect 29922 8316 29932 8372
rect 29988 8316 31612 8372
rect 31668 8316 31678 8372
rect 23202 8204 23212 8260
rect 23268 8204 23548 8260
rect 23604 8204 23614 8260
rect 27794 8204 27804 8260
rect 27860 8204 28476 8260
rect 28532 8204 28542 8260
rect 12562 7980 12572 8036
rect 12628 7980 13580 8036
rect 13636 7980 13646 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 26786 6860 26796 6916
rect 26852 6860 27804 6916
rect 27860 6860 27870 6916
rect 9986 6636 9996 6692
rect 10052 6636 12124 6692
rect 12180 6636 13580 6692
rect 13636 6636 13646 6692
rect 25778 6524 25788 6580
rect 25844 6524 26236 6580
rect 26292 6524 27132 6580
rect 27188 6524 27804 6580
rect 27860 6524 27870 6580
rect 26562 6300 26572 6356
rect 26628 6300 26908 6356
rect 26964 6300 26974 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 13682 6076 13692 6132
rect 13748 6076 15372 6132
rect 15428 6076 15438 6132
rect 24546 5964 24556 6020
rect 24612 5964 26460 6020
rect 26516 5964 26526 6020
rect 23314 5740 23324 5796
rect 23380 5740 25676 5796
rect 25732 5740 25742 5796
rect 26898 5628 26908 5684
rect 26964 5628 27804 5684
rect 27860 5628 27870 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 27010 4508 27020 4564
rect 27076 4508 30268 4564
rect 30324 4508 30334 4564
rect 27458 4172 27468 4228
rect 27524 4172 29820 4228
rect 29876 4172 29886 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19628 20524 19684 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 19628 20188 19684 20244
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 42396
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 19808 42364 20128 42396
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19628 20580 19684 20590
rect 19628 20244 19684 20524
rect 19628 20178 19684 20188
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 41580 35488 42396
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _330_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31696 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _331_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32144 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _332_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32256 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _333_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29680 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _334_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31584 0 -1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _335_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27216 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _336_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26208 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _337_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14112 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _338_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _339_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _340_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _341_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8400 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _342_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _343_
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _344_
timestamp 1698431365
transform -1 0 30016 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _345_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25760 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _346_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20160 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _347_
timestamp 1698431365
transform 1 0 14336 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _348_
timestamp 1698431365
transform 1 0 5040 0 -1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _349_
timestamp 1698431365
transform 1 0 6496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _350_
timestamp 1698431365
transform 1 0 9184 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _351_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10640 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _352_
timestamp 1698431365
transform 1 0 13664 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _353_
timestamp 1698431365
transform -1 0 15680 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _354_
timestamp 1698431365
transform -1 0 14560 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _355_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15120 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _356_
timestamp 1698431365
transform 1 0 9632 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _357_
timestamp 1698431365
transform -1 0 22512 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _358_
timestamp 1698431365
transform -1 0 16016 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _359_
timestamp 1698431365
transform -1 0 16912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _360_
timestamp 1698431365
transform -1 0 17808 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _361_
timestamp 1698431365
transform 1 0 14448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _362_
timestamp 1698431365
transform 1 0 15456 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _363_
timestamp 1698431365
transform -1 0 16464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _364_
timestamp 1698431365
transform -1 0 17696 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _365_
timestamp 1698431365
transform -1 0 16464 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _366_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _367_
timestamp 1698431365
transform 1 0 6832 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _368_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _369_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11760 0 1 29792
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _370_
timestamp 1698431365
transform 1 0 14896 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _371_
timestamp 1698431365
transform 1 0 19264 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _372_
timestamp 1698431365
transform -1 0 31920 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _373_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31136 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _374_
timestamp 1698431365
transform -1 0 26096 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _375_
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _376_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25648 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _377_
timestamp 1698431365
transform -1 0 22848 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _378_
timestamp 1698431365
transform 1 0 8624 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _379_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _380_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _381_
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _382_
timestamp 1698431365
transform -1 0 20272 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _383_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22064 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _384_
timestamp 1698431365
transform -1 0 26768 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _385_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26096 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _386_
timestamp 1698431365
transform 1 0 25536 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _387_
timestamp 1698431365
transform -1 0 26768 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _388_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _389_
timestamp 1698431365
transform -1 0 26992 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _390_
timestamp 1698431365
transform 1 0 19936 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _391_
timestamp 1698431365
transform -1 0 20832 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _392_
timestamp 1698431365
transform 1 0 22960 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _393_
timestamp 1698431365
transform -1 0 22064 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _394_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _395_
timestamp 1698431365
transform -1 0 20496 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _396_
timestamp 1698431365
transform 1 0 18704 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _397_
timestamp 1698431365
transform -1 0 24752 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _398_
timestamp 1698431365
transform -1 0 21392 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _399_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25984 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _400_
timestamp 1698431365
transform -1 0 24864 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _401_
timestamp 1698431365
transform -1 0 20720 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _402_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24192 0 1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _403_
timestamp 1698431365
transform -1 0 25984 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _404_
timestamp 1698431365
transform -1 0 24528 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _405_
timestamp 1698431365
transform 1 0 26992 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _406_
timestamp 1698431365
transform 1 0 25424 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _407_
timestamp 1698431365
transform 1 0 23296 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _408_
timestamp 1698431365
transform 1 0 20048 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _409_
timestamp 1698431365
transform 1 0 24304 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _410_
timestamp 1698431365
transform -1 0 24304 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _411_
timestamp 1698431365
transform -1 0 15120 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _412_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _413_
timestamp 1698431365
transform -1 0 24192 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _414_
timestamp 1698431365
transform 1 0 22064 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _415_
timestamp 1698431365
transform -1 0 22288 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _416_
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _417_
timestamp 1698431365
transform -1 0 26656 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _418_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _419_
timestamp 1698431365
transform -1 0 25984 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _420_
timestamp 1698431365
transform 1 0 26992 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _421_
timestamp 1698431365
transform 1 0 25424 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _422_
timestamp 1698431365
transform 1 0 34608 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _423_
timestamp 1698431365
transform 1 0 27328 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _424_
timestamp 1698431365
transform 1 0 26096 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _425_
timestamp 1698431365
transform 1 0 27664 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _426_
timestamp 1698431365
transform -1 0 26656 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _427_
timestamp 1698431365
transform -1 0 26208 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _428_
timestamp 1698431365
transform -1 0 27328 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _429_
timestamp 1698431365
transform -1 0 28112 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _430_
timestamp 1698431365
transform -1 0 22848 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _431_
timestamp 1698431365
transform -1 0 23520 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _432_
timestamp 1698431365
transform -1 0 22960 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _433_
timestamp 1698431365
transform -1 0 25872 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _434_
timestamp 1698431365
transform 1 0 23072 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _435_
timestamp 1698431365
transform -1 0 23856 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _436_
timestamp 1698431365
transform 1 0 22848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _437_
timestamp 1698431365
transform 1 0 28000 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _438_
timestamp 1698431365
transform 1 0 29904 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _439_
timestamp 1698431365
transform 1 0 27104 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _440_
timestamp 1698431365
transform 1 0 29232 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _441_
timestamp 1698431365
transform -1 0 34272 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _442_
timestamp 1698431365
transform 1 0 32704 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _443_
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _444_
timestamp 1698431365
transform 1 0 30128 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _445_
timestamp 1698431365
transform -1 0 30912 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _446_
timestamp 1698431365
transform -1 0 30128 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _447_
timestamp 1698431365
transform -1 0 30016 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _448_
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _449_
timestamp 1698431365
transform 1 0 30016 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _450_
timestamp 1698431365
transform -1 0 30352 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _451_
timestamp 1698431365
transform -1 0 29008 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _452_
timestamp 1698431365
transform -1 0 24304 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _453_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _454_
timestamp 1698431365
transform 1 0 31248 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _455_
timestamp 1698431365
transform 1 0 31920 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _456_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _457_
timestamp 1698431365
transform 1 0 35616 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _458_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27216 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _459_
timestamp 1698431365
transform -1 0 32704 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _460_
timestamp 1698431365
transform 1 0 39088 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _461_
timestamp 1698431365
transform -1 0 38304 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _462_
timestamp 1698431365
transform -1 0 39536 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _463_
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _464_
timestamp 1698431365
transform 1 0 33936 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _465_
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _466_
timestamp 1698431365
transform 1 0 35168 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _467_
timestamp 1698431365
transform -1 0 35392 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _468_
timestamp 1698431365
transform 1 0 38864 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _469_
timestamp 1698431365
transform -1 0 37408 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _470_
timestamp 1698431365
transform -1 0 36176 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _471_
timestamp 1698431365
transform 1 0 36960 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _472_
timestamp 1698431365
transform -1 0 37408 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _473_
timestamp 1698431365
transform 1 0 36960 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _474_
timestamp 1698431365
transform 1 0 35840 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _475_
timestamp 1698431365
transform 1 0 39872 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _476_
timestamp 1698431365
transform 1 0 40880 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _477_
timestamp 1698431365
transform 1 0 39648 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _478_
timestamp 1698431365
transform -1 0 42336 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _479_
timestamp 1698431365
transform 1 0 40880 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _480_
timestamp 1698431365
transform 1 0 40096 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _481_
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _482_
timestamp 1698431365
transform 1 0 37520 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _483_
timestamp 1698431365
transform 1 0 40544 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _484_
timestamp 1698431365
transform -1 0 40544 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _485_
timestamp 1698431365
transform -1 0 40880 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _486_
timestamp 1698431365
transform 1 0 36960 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _487_
timestamp 1698431365
transform 1 0 37744 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _488_
timestamp 1698431365
transform 1 0 41440 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _489_
timestamp 1698431365
transform 1 0 40208 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _490_
timestamp 1698431365
transform 1 0 41104 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _491_
timestamp 1698431365
transform 1 0 39536 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _492_
timestamp 1698431365
transform -1 0 42112 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _493_
timestamp 1698431365
transform 1 0 39088 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _494_
timestamp 1698431365
transform 1 0 42224 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _495_
timestamp 1698431365
transform -1 0 42224 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _496_
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _497_
timestamp 1698431365
transform -1 0 42672 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _498_
timestamp 1698431365
transform 1 0 39312 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _499_
timestamp 1698431365
transform -1 0 42112 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _500_
timestamp 1698431365
transform 1 0 31808 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _501_
timestamp 1698431365
transform -1 0 36960 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _502_
timestamp 1698431365
transform -1 0 35504 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _503_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36176 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _504_
timestamp 1698431365
transform -1 0 35056 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _505_
timestamp 1698431365
transform 1 0 40208 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _506_
timestamp 1698431365
transform -1 0 41888 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _507_
timestamp 1698431365
transform -1 0 41664 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _508_
timestamp 1698431365
transform 1 0 35168 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _509_
timestamp 1698431365
transform -1 0 36400 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _510_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _511_
timestamp 1698431365
transform 1 0 37296 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _512_
timestamp 1698431365
transform -1 0 38304 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _513_
timestamp 1698431365
transform -1 0 36848 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _514_
timestamp 1698431365
transform -1 0 36624 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _515_
timestamp 1698431365
transform -1 0 35616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _516_
timestamp 1698431365
transform -1 0 42560 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _517_
timestamp 1698431365
transform 1 0 40432 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _518_
timestamp 1698431365
transform 1 0 41440 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _519_
timestamp 1698431365
transform 1 0 31136 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _520_
timestamp 1698431365
transform 1 0 35728 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _521_
timestamp 1698431365
transform 1 0 38976 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _522_
timestamp 1698431365
transform 1 0 39200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _523_
timestamp 1698431365
transform -1 0 18144 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _524_
timestamp 1698431365
transform -1 0 18928 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _525_
timestamp 1698431365
transform -1 0 15456 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _526_
timestamp 1698431365
transform -1 0 14000 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _527_
timestamp 1698431365
transform 1 0 14336 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _528_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _529_
timestamp 1698431365
transform 1 0 9968 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _530_
timestamp 1698431365
transform 1 0 10976 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _531_
timestamp 1698431365
transform 1 0 12544 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _532_
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _533_
timestamp 1698431365
transform 1 0 17808 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _534_
timestamp 1698431365
transform -1 0 17696 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _535_
timestamp 1698431365
transform 1 0 18704 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _536_
timestamp 1698431365
transform -1 0 12096 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _537_
timestamp 1698431365
transform 1 0 10976 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _538_
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _539_
timestamp 1698431365
transform 1 0 19040 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _540_
timestamp 1698431365
transform 1 0 20496 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _541_
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _542_
timestamp 1698431365
transform 1 0 18144 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _543_
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _544_
timestamp 1698431365
transform 1 0 19152 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _545_
timestamp 1698431365
transform 1 0 21280 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _546_
timestamp 1698431365
transform -1 0 14336 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _547_
timestamp 1698431365
transform -1 0 18144 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _548_
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _549_
timestamp 1698431365
transform -1 0 16128 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _550_
timestamp 1698431365
transform -1 0 14896 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _551_
timestamp 1698431365
transform -1 0 12544 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _552_
timestamp 1698431365
transform 1 0 7728 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _553_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17472 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _554_
timestamp 1698431365
transform 1 0 10304 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _555_
timestamp 1698431365
transform 1 0 10864 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _556_
timestamp 1698431365
transform -1 0 11088 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _557_
timestamp 1698431365
transform -1 0 10080 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _558_
timestamp 1698431365
transform -1 0 9184 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _559_
timestamp 1698431365
transform -1 0 8512 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _560_
timestamp 1698431365
transform -1 0 6832 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _561_
timestamp 1698431365
transform -1 0 4256 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _562_
timestamp 1698431365
transform -1 0 9520 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _563_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _564_
timestamp 1698431365
transform -1 0 6496 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _565_
timestamp 1698431365
transform -1 0 4368 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _566_
timestamp 1698431365
transform -1 0 13888 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _567_
timestamp 1698431365
transform 1 0 5376 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _568_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11648 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _569_
timestamp 1698431365
transform 1 0 5152 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _570_
timestamp 1698431365
transform -1 0 6496 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _571_
timestamp 1698431365
transform -1 0 4592 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _572_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _573_
timestamp 1698431365
transform -1 0 6608 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _574_
timestamp 1698431365
transform 1 0 6272 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _575_
timestamp 1698431365
transform -1 0 7392 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _576_
timestamp 1698431365
transform 1 0 5488 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _577_
timestamp 1698431365
transform -1 0 5488 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _578_
timestamp 1698431365
transform -1 0 8848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _579_
timestamp 1698431365
transform -1 0 10976 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _580_
timestamp 1698431365
transform 1 0 6832 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _581_
timestamp 1698431365
transform 1 0 7392 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _582_
timestamp 1698431365
transform -1 0 8288 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _583_
timestamp 1698431365
transform 1 0 9520 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _584_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _585_
timestamp 1698431365
transform -1 0 24976 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _586_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7280 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _587_
timestamp 1698431365
transform -1 0 7616 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _588_
timestamp 1698431365
transform 1 0 6496 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _589_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20384 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _590_
timestamp 1698431365
transform -1 0 20272 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _591_
timestamp 1698431365
transform -1 0 14560 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _592_
timestamp 1698431365
transform 1 0 7056 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _593_
timestamp 1698431365
transform 1 0 7056 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _594_
timestamp 1698431365
transform -1 0 6944 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _595_
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _596_
timestamp 1698431365
transform -1 0 8960 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _597_
timestamp 1698431365
transform 1 0 7952 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _598_
timestamp 1698431365
transform -1 0 9072 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _599_
timestamp 1698431365
transform 1 0 7392 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _600_
timestamp 1698431365
transform 1 0 7616 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _601_
timestamp 1698431365
transform -1 0 14000 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _602_
timestamp 1698431365
transform 1 0 11536 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _603_
timestamp 1698431365
transform 1 0 10080 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _604_
timestamp 1698431365
transform -1 0 11984 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _605_
timestamp 1698431365
transform -1 0 11312 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _606_
timestamp 1698431365
transform -1 0 14784 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _607_
timestamp 1698431365
transform 1 0 12096 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _608_
timestamp 1698431365
transform 1 0 12320 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _609_
timestamp 1698431365
transform 1 0 12096 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _610_
timestamp 1698431365
transform 1 0 12208 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _611_
timestamp 1698431365
transform -1 0 15456 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _612_
timestamp 1698431365
transform 1 0 15792 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _613_
timestamp 1698431365
transform 1 0 13552 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _614_
timestamp 1698431365
transform 1 0 14672 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _615_
timestamp 1698431365
transform 1 0 16576 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _616_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17024 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _617_
timestamp 1698431365
transform 1 0 18256 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _618_
timestamp 1698431365
transform -1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _619_
timestamp 1698431365
transform 1 0 15568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _620_
timestamp 1698431365
transform -1 0 19600 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _621_
timestamp 1698431365
transform 1 0 18032 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _622_
timestamp 1698431365
transform -1 0 13104 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _623_
timestamp 1698431365
transform -1 0 11424 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _624_
timestamp 1698431365
transform -1 0 10304 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _625_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _626_
timestamp 1698431365
transform -1 0 4928 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _627_
timestamp 1698431365
transform -1 0 9072 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _628_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _629_
timestamp 1698431365
transform -1 0 5376 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _630_
timestamp 1698431365
transform 1 0 12208 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _631_
timestamp 1698431365
transform -1 0 19376 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _632_
timestamp 1698431365
transform 1 0 12544 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _633_
timestamp 1698431365
transform 1 0 11536 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _634_
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _635_
timestamp 1698431365
transform -1 0 25760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _636_
timestamp 1698431365
transform 1 0 18704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _637_
timestamp 1698431365
transform 1 0 16240 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _638_
timestamp 1698431365
transform 1 0 14896 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _639_
timestamp 1698431365
transform 1 0 15232 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _640_
timestamp 1698431365
transform 1 0 11424 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _641_
timestamp 1698431365
transform -1 0 12544 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _642_
timestamp 1698431365
transform 1 0 11648 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _643_
timestamp 1698431365
transform 1 0 6384 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _644_
timestamp 1698431365
transform -1 0 7952 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _645_
timestamp 1698431365
transform 1 0 10640 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _646_
timestamp 1698431365
transform -1 0 10640 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _647_
timestamp 1698431365
transform 1 0 10640 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _648_
timestamp 1698431365
transform 1 0 6720 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _649_
timestamp 1698431365
transform 1 0 6496 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _650_
timestamp 1698431365
transform -1 0 32032 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _651_
timestamp 1698431365
transform -1 0 30688 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _652_
timestamp 1698431365
transform 1 0 30016 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _653_
timestamp 1698431365
transform 1 0 29568 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _654_
timestamp 1698431365
transform 1 0 28448 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _655_
timestamp 1698431365
transform 1 0 29008 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _656_
timestamp 1698431365
transform -1 0 28784 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _657_
timestamp 1698431365
transform -1 0 27552 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _658_
timestamp 1698431365
transform 1 0 30576 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _659_
timestamp 1698431365
transform 1 0 31584 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _660_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13104 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _661_
timestamp 1698431365
transform 1 0 9632 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _662_
timestamp 1698431365
transform -1 0 26656 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _663_
timestamp 1698431365
transform 1 0 27552 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _664_
timestamp 1698431365
transform 1 0 29568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _665_
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _666_
timestamp 1698431365
transform 1 0 17472 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _667_
timestamp 1698431365
transform 1 0 19712 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _668_
timestamp 1698431365
transform -1 0 25984 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _669_
timestamp 1698431365
transform 1 0 26768 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _670_
timestamp 1698431365
transform 1 0 21504 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _671_
timestamp 1698431365
transform 1 0 21616 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _672_
timestamp 1698431365
transform -1 0 32592 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _673_
timestamp 1698431365
transform -1 0 36176 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _674_
timestamp 1698431365
transform 1 0 27888 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _675_
timestamp 1698431365
transform -1 0 32256 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _676_
timestamp 1698431365
transform 1 0 24304 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _677_
timestamp 1698431365
transform -1 0 30688 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _678_
timestamp 1698431365
transform 1 0 15680 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _679_
timestamp 1698431365
transform 1 0 4704 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _680_
timestamp 1698431365
transform -1 0 37968 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _681_
timestamp 1698431365
transform 1 0 34832 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _682_
timestamp 1698431365
transform -1 0 36960 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _683_
timestamp 1698431365
transform 1 0 40880 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _684_
timestamp 1698431365
transform -1 0 42336 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _685_
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _686_
timestamp 1698431365
transform -1 0 37744 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _687_
timestamp 1698431365
transform 1 0 40768 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _688_
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _689_
timestamp 1698431365
transform 1 0 40992 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _690_
timestamp 1698431365
transform 1 0 33376 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _691_
timestamp 1698431365
transform 1 0 40320 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _692_
timestamp 1698431365
transform 1 0 37184 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _693_
timestamp 1698431365
transform 1 0 33376 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _694_
timestamp 1698431365
transform 1 0 40992 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _695_
timestamp 1698431365
transform 1 0 38752 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _696_
timestamp 1698431365
transform 1 0 15008 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _697_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23408 0 -1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _698_
timestamp 1698431365
transform -1 0 24528 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _699_
timestamp 1698431365
transform 1 0 13440 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _700_
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _701_
timestamp 1698431365
transform 1 0 1680 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _702_
timestamp 1698431365
transform 1 0 1680 0 -1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _703_
timestamp 1698431365
transform 1 0 1680 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _704_
timestamp 1698431365
transform 1 0 1680 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _705_
timestamp 1698431365
transform 1 0 1792 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _706_
timestamp 1698431365
transform 1 0 3584 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _707_
timestamp 1698431365
transform 1 0 1680 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _708_
timestamp 1698431365
transform 1 0 9744 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _709_
timestamp 1698431365
transform 1 0 11872 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _710_
timestamp 1698431365
transform -1 0 20832 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _711_
timestamp 1698431365
transform -1 0 20496 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _712_
timestamp 1698431365
transform 1 0 1680 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _713_
timestamp 1698431365
transform 1 0 2016 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _714_
timestamp 1698431365
transform 1 0 19600 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _715_
timestamp 1698431365
transform -1 0 16912 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _716_
timestamp 1698431365
transform 1 0 10752 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _717_
timestamp 1698431365
transform 1 0 2016 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _718_
timestamp 1698431365
transform -1 0 10864 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _719_
timestamp 1698431365
transform 1 0 2128 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _720_
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _721_
timestamp 1698431365
transform 1 0 26768 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _722_
timestamp 1698431365
transform 1 0 25200 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _723_
timestamp 1698431365
transform 1 0 30352 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__A3 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__A4
timestamp 1698431365
transform 1 0 15456 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__B
timestamp 1698431365
transform 1 0 20384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__A1
timestamp 1698431365
transform -1 0 15344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__A2
timestamp 1698431365
transform -1 0 13328 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__I
timestamp 1698431365
transform 1 0 17136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__I
timestamp 1698431365
transform 1 0 14224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__A1
timestamp 1698431365
transform 1 0 14560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__B2
timestamp 1698431365
transform -1 0 15456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__I
timestamp 1698431365
transform 1 0 6608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__B1
timestamp 1698431365
transform -1 0 12208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__379__I
timestamp 1698431365
transform -1 0 19936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__I
timestamp 1698431365
transform 1 0 19712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__A1
timestamp 1698431365
transform 1 0 26544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__B
timestamp 1698431365
transform -1 0 24192 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A1
timestamp 1698431365
transform -1 0 25536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__I
timestamp 1698431365
transform -1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__I
timestamp 1698431365
transform 1 0 22960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__I
timestamp 1698431365
transform -1 0 23856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__I
timestamp 1698431365
transform 1 0 25760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__I
timestamp 1698431365
transform 1 0 34384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__A1
timestamp 1698431365
transform 1 0 25872 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__A1
timestamp 1698431365
transform -1 0 23072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__B
timestamp 1698431365
transform 1 0 24080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__B
timestamp 1698431365
transform 1 0 32480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__B
timestamp 1698431365
transform -1 0 30016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__I
timestamp 1698431365
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__I
timestamp 1698431365
transform 1 0 31024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__I
timestamp 1698431365
transform -1 0 32032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__I
timestamp 1698431365
transform 1 0 38864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__I
timestamp 1698431365
transform 1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__I
timestamp 1698431365
transform 1 0 33712 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__I
timestamp 1698431365
transform -1 0 33152 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__I
timestamp 1698431365
transform 1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A1
timestamp 1698431365
transform -1 0 34832 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__I
timestamp 1698431365
transform -1 0 35840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__493__I
timestamp 1698431365
transform 1 0 38864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__I
timestamp 1698431365
transform 1 0 39088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__A1
timestamp 1698431365
transform -1 0 34944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__C
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__A1
timestamp 1698431365
transform 1 0 35616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__C
timestamp 1698431365
transform 1 0 37184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__C
timestamp 1698431365
transform 1 0 35280 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__A2
timestamp 1698431365
transform -1 0 35728 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__A2
timestamp 1698431365
transform 1 0 38752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__526__A1
timestamp 1698431365
transform 1 0 14224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__I
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A2
timestamp 1698431365
transform -1 0 9968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__A2
timestamp 1698431365
transform 1 0 12320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__C
timestamp 1698431365
transform 1 0 19152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__I
timestamp 1698431365
transform 1 0 19600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__A1
timestamp 1698431365
transform 1 0 12320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__B2
timestamp 1698431365
transform -1 0 19040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__I
timestamp 1698431365
transform 1 0 14560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__553__A3
timestamp 1698431365
transform 1 0 17696 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__566__I
timestamp 1698431365
transform 1 0 14784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__571__A1
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__576__B
timestamp 1698431365
transform 1 0 6832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__I
timestamp 1698431365
transform 1 0 24080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__586__C
timestamp 1698431365
transform 1 0 9072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__A1
timestamp 1698431365
transform -1 0 20720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__A2
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__592__B2
timestamp 1698431365
transform -1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__593__B
timestamp 1698431365
transform 1 0 7952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__598__B2
timestamp 1698431365
transform 1 0 9296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__C
timestamp 1698431365
transform 1 0 9632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__B
timestamp 1698431365
transform -1 0 12880 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__605__A1
timestamp 1698431365
transform 1 0 11536 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__610__A1
timestamp 1698431365
transform 1 0 13552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__620__A1
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__A1
timestamp 1698431365
transform 1 0 11648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__624__A1
timestamp 1698431365
transform -1 0 10752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__625__S
timestamp 1698431365
transform 1 0 6944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__626__A1
timestamp 1698431365
transform 1 0 5600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__A2
timestamp 1698431365
transform 1 0 9632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__A2
timestamp 1698431365
transform 1 0 10976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__B2
timestamp 1698431365
transform 1 0 6944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__C
timestamp 1698431365
transform -1 0 9968 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__A1
timestamp 1698431365
transform 1 0 19600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__A2
timestamp 1698431365
transform 1 0 17024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__635__I
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__636__B
timestamp 1698431365
transform -1 0 19824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__637__A1
timestamp 1698431365
transform 1 0 17920 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__638__A2
timestamp 1698431365
transform 1 0 14672 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__639__B
timestamp 1698431365
transform 1 0 16352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__640__A1
timestamp 1698431365
transform 1 0 13104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__641__A2
timestamp 1698431365
transform -1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__642__B
timestamp 1698431365
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__643__A1
timestamp 1698431365
transform -1 0 7392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__644__C
timestamp 1698431365
transform 1 0 8176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__645__A1
timestamp 1698431365
transform 1 0 11424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__A2
timestamp 1698431365
transform 1 0 10640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__B
timestamp 1698431365
transform 1 0 12432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__648__A1
timestamp 1698431365
transform 1 0 7728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__649__C
timestamp 1698431365
transform 1 0 8512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__650__A2
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__651__A1
timestamp 1698431365
transform 1 0 29792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__652__A2
timestamp 1698431365
transform 1 0 31248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__654__A1
timestamp 1698431365
transform 1 0 29904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__A1
timestamp 1698431365
transform 1 0 26656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__658__A1
timestamp 1698431365
transform 1 0 29680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__658__B1
timestamp 1698431365
transform 1 0 30128 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__659__A1
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__660__CLK
timestamp 1698431365
transform 1 0 16352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__661__CLK
timestamp 1698431365
transform 1 0 12880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__662__CLK
timestamp 1698431365
transform 1 0 26880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__663__CLK
timestamp 1698431365
transform -1 0 31248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__664__CLK
timestamp 1698431365
transform 1 0 33040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__665__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__666__CLK
timestamp 1698431365
transform -1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__667__CLK
timestamp 1698431365
transform 1 0 19488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__668__CLK
timestamp 1698431365
transform 1 0 26208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__669__CLK
timestamp 1698431365
transform 1 0 30240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__670__CLK
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__671__CLK
timestamp 1698431365
transform 1 0 21392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__672__CLK
timestamp 1698431365
transform -1 0 33040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__CLK
timestamp 1698431365
transform 1 0 31360 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__676__CLK
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__677__CLK
timestamp 1698431365
transform 1 0 30912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__CLK
timestamp 1698431365
transform 1 0 19152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__679__CLK
timestamp 1698431365
transform -1 0 8400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__679__D
timestamp 1698431365
transform -1 0 8848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__680__CLK
timestamp 1698431365
transform 1 0 38192 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__CLK
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__CLK
timestamp 1698431365
transform 1 0 38080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__683__CLK
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__684__CLK
timestamp 1698431365
transform 1 0 38864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__685__CLK
timestamp 1698431365
transform 1 0 39424 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__CLK
timestamp 1698431365
transform 1 0 38752 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__687__CLK
timestamp 1698431365
transform 1 0 39984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__688__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__690__CLK
timestamp 1698431365
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__691__CLK
timestamp 1698431365
transform 1 0 40096 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__692__CLK
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__693__CLK
timestamp 1698431365
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__694__CLK
timestamp 1698431365
transform 1 0 40208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__695__CLK
timestamp 1698431365
transform -1 0 38752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__696__CLK
timestamp 1698431365
transform 1 0 18480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__697__CLK
timestamp 1698431365
transform 1 0 23632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__CLK
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__699__CLK
timestamp 1698431365
transform -1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__700__CLK
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__702__CLK
timestamp 1698431365
transform -1 0 5600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__703__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__704__CLK
timestamp 1698431365
transform 1 0 4928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__705__CLK
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__706__CLK
timestamp 1698431365
transform 1 0 7056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__CLK
timestamp 1698431365
transform 1 0 13552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__CLK
timestamp 1698431365
transform 1 0 15344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__CLK
timestamp 1698431365
transform 1 0 20720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__CLK
timestamp 1698431365
transform 1 0 5712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__CLK
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__714__CLK
timestamp 1698431365
transform 1 0 19376 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__715__CLK
timestamp 1698431365
transform 1 0 17136 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__CLK
timestamp 1698431365
transform 1 0 14224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__717__CLK
timestamp 1698431365
transform 1 0 5712 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__718__CLK
timestamp 1698431365
transform 1 0 11088 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__719__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__720__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__721__CLK
timestamp 1698431365
transform 1 0 30016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__722__CLK
timestamp 1698431365
transform 1 0 28672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__723__CLK
timestamp 1698431365
transform 1 0 33824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 22064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 21392 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 16352 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 20608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 33376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 30576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 33600 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22064 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1698431365
transform 1 0 10752 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1698431365
transform 1 0 15344 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1698431365
transform -1 0 16128 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 14000 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1698431365
transform 1 0 30576 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_376 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_174
timestamp 1698431365
transform 1 0 20832 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_182
timestamp 1698431365
transform 1 0 21728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_186 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22176 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_193 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22960 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_224 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_226
timestamp 1698431365
transform 1 0 26656 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_256
timestamp 1698431365
transform 1 0 30016 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_260
timestamp 1698431365
transform 1 0 30464 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_179
timestamp 1698431365
transform 1 0 21392 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_209
timestamp 1698431365
transform 1 0 24752 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_383
timestamp 1698431365
transform 1 0 44240 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_88
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_92
timestamp 1698431365
transform 1 0 11648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_123
timestamp 1698431365
transform 1 0 15120 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_127
timestamp 1698431365
transform 1 0 15568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_135
timestamp 1698431365
transform 1 0 16464 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_174
timestamp 1698431365
transform 1 0 20832 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_198
timestamp 1698431365
transform 1 0 23520 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_216
timestamp 1698431365
transform 1 0 25536 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_226
timestamp 1698431365
transform 1 0 26656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_228
timestamp 1698431365
transform 1 0 26880 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_241
timestamp 1698431365
transform 1 0 28336 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_273
timestamp 1698431365
transform 1 0 31920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_277
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_73
timestamp 1698431365
transform 1 0 9520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_111
timestamp 1698431365
transform 1 0 13776 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_209
timestamp 1698431365
transform 1 0 24752 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_217
timestamp 1698431365
transform 1 0 25648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_237
timestamp 1698431365
transform 1 0 27888 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_383
timestamp 1698431365
transform 1 0 44240 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_171
timestamp 1698431365
transform 1 0 20496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_175
timestamp 1698431365
transform 1 0 20944 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_191
timestamp 1698431365
transform 1 0 22736 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_194
timestamp 1698431365
transform 1 0 23072 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_218
timestamp 1698431365
transform 1 0 25760 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_256
timestamp 1698431365
transform 1 0 30016 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_272
timestamp 1698431365
transform 1 0 31808 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_77
timestamp 1698431365
transform 1 0 9968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_81
timestamp 1698431365
transform 1 0 10416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_89
timestamp 1698431365
transform 1 0 11312 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_93
timestamp 1698431365
transform 1 0 11760 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_111
timestamp 1698431365
transform 1 0 13776 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_143
timestamp 1698431365
transform 1 0 17360 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_147
timestamp 1698431365
transform 1 0 17808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_155
timestamp 1698431365
transform 1 0 18704 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_185
timestamp 1698431365
transform 1 0 22064 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_200
timestamp 1698431365
transform 1 0 23744 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_232
timestamp 1698431365
transform 1 0 27328 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_239
timestamp 1698431365
transform 1 0 28112 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_249
timestamp 1698431365
transform 1 0 29232 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_279
timestamp 1698431365
transform 1 0 32592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_283
timestamp 1698431365
transform 1 0 33040 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_18
timestamp 1698431365
transform 1 0 3360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_49
timestamp 1698431365
transform 1 0 6832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_53
timestamp 1698431365
transform 1 0 7280 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_104
timestamp 1698431365
transform 1 0 12992 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_112
timestamp 1698431365
transform 1 0 13888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_120
timestamp 1698431365
transform 1 0 14784 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_128
timestamp 1698431365
transform 1 0 15680 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_132
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_174
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_178
timestamp 1698431365
transform 1 0 21280 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_219
timestamp 1698431365
transform 1 0 25872 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_227
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_229
timestamp 1698431365
transform 1 0 26992 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_248
timestamp 1698431365
transform 1 0 29120 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_41
timestamp 1698431365
transform 1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_43
timestamp 1698431365
transform 1 0 6160 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_56
timestamp 1698431365
transform 1 0 7616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_58
timestamp 1698431365
transform 1 0 7840 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_61
timestamp 1698431365
transform 1 0 8176 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_93
timestamp 1698431365
transform 1 0 11760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_95
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_113
timestamp 1698431365
transform 1 0 14000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_163
timestamp 1698431365
transform 1 0 19600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_167
timestamp 1698431365
transform 1 0 20048 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_201
timestamp 1698431365
transform 1 0 23856 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_205
timestamp 1698431365
transform 1 0 24304 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_237
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_257
timestamp 1698431365
transform 1 0 30128 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_289
timestamp 1698431365
transform 1 0 33712 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_305
timestamp 1698431365
transform 1 0 35504 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_383
timestamp 1698431365
transform 1 0 44240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_50
timestamp 1698431365
transform 1 0 6944 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_76
timestamp 1698431365
transform 1 0 9856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_95
timestamp 1698431365
transform 1 0 11984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_97
timestamp 1698431365
transform 1 0 12208 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_106
timestamp 1698431365
transform 1 0 13216 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_126
timestamp 1698431365
transform 1 0 15456 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_135
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_244
timestamp 1698431365
transform 1 0 28672 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_252
timestamp 1698431365
transform 1 0 29568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_254
timestamp 1698431365
transform 1 0 29792 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_261
timestamp 1698431365
transform 1 0 30576 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_73
timestamp 1698431365
transform 1 0 9520 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_89
timestamp 1698431365
transform 1 0 11312 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_93
timestamp 1698431365
transform 1 0 11760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_95
timestamp 1698431365
transform 1 0 11984 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_114
timestamp 1698431365
transform 1 0 14112 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_130
timestamp 1698431365
transform 1 0 15904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_134
timestamp 1698431365
transform 1 0 16352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_158
timestamp 1698431365
transform 1 0 19040 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_253
timestamp 1698431365
transform 1 0 29680 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_264
timestamp 1698431365
transform 1 0 30912 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_272
timestamp 1698431365
transform 1 0 31808 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_276
timestamp 1698431365
transform 1 0 32256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_288
timestamp 1698431365
transform 1 0 33600 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_304
timestamp 1698431365
transform 1 0 35392 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_312
timestamp 1698431365
transform 1 0 36288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_383
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_32
timestamp 1698431365
transform 1 0 4928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_36
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_46
timestamp 1698431365
transform 1 0 6496 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_76
timestamp 1698431365
transform 1 0 9856 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_84
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_88
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_90
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_99
timestamp 1698431365
transform 1 0 12432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_103
timestamp 1698431365
transform 1 0 12880 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_134
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_174
timestamp 1698431365
transform 1 0 20832 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_236
timestamp 1698431365
transform 1 0 27776 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_266
timestamp 1698431365
transform 1 0 31136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_270
timestamp 1698431365
transform 1 0 31584 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_311
timestamp 1698431365
transform 1 0 36176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_315
timestamp 1698431365
transform 1 0 36624 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_347
timestamp 1698431365
transform 1 0 40208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_53
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_55
timestamp 1698431365
transform 1 0 7504 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_66
timestamp 1698431365
transform 1 0 8736 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_98
timestamp 1698431365
transform 1 0 12320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_189
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_220
timestamp 1698431365
transform 1 0 25984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_224
timestamp 1698431365
transform 1 0 26432 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_240
timestamp 1698431365
transform 1 0 28224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_265
timestamp 1698431365
transform 1 0 31024 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_273
timestamp 1698431365
transform 1 0 31920 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_277
timestamp 1698431365
transform 1 0 32368 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_279
timestamp 1698431365
transform 1 0 32592 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_294
timestamp 1698431365
transform 1 0 34272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_296
timestamp 1698431365
transform 1 0 34496 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_305
timestamp 1698431365
transform 1 0 35504 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_313
timestamp 1698431365
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_383
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_34
timestamp 1698431365
transform 1 0 5152 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_50
timestamp 1698431365
transform 1 0 6944 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_54
timestamp 1698431365
transform 1 0 7392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_62
timestamp 1698431365
transform 1 0 8288 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_158
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_193
timestamp 1698431365
transform 1 0 22960 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_201
timestamp 1698431365
transform 1 0 23856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_203
timestamp 1698431365
transform 1 0 24080 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_226
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_258
timestamp 1698431365
transform 1 0 30240 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_294
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_297
timestamp 1698431365
transform 1 0 34608 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_329
timestamp 1698431365
transform 1 0 38192 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_345
timestamp 1698431365
transform 1 0 39984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_30
timestamp 1698431365
transform 1 0 4704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_32
timestamp 1698431365
transform 1 0 4928 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_69
timestamp 1698431365
transform 1 0 9072 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_79
timestamp 1698431365
transform 1 0 10192 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_95
timestamp 1698431365
transform 1 0 11984 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_113
timestamp 1698431365
transform 1 0 14000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_117
timestamp 1698431365
transform 1 0 14448 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_121
timestamp 1698431365
transform 1 0 14896 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_151
timestamp 1698431365
transform 1 0 18256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_155
timestamp 1698431365
transform 1 0 18704 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_209
timestamp 1698431365
transform 1 0 24752 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_217
timestamp 1698431365
transform 1 0 25648 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_220
timestamp 1698431365
transform 1 0 25984 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_236
timestamp 1698431365
transform 1 0 27776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_251
timestamp 1698431365
transform 1 0 29456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_253
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_256
timestamp 1698431365
transform 1 0 30016 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_288
timestamp 1698431365
transform 1 0 33600 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_304
timestamp 1698431365
transform 1 0 35392 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_319
timestamp 1698431365
transform 1 0 37072 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_349
timestamp 1698431365
transform 1 0 40432 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_383
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_96
timestamp 1698431365
transform 1 0 12096 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_118
timestamp 1698431365
transform 1 0 14560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_122
timestamp 1698431365
transform 1 0 15008 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_174
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_178
timestamp 1698431365
transform 1 0 21280 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_180
timestamp 1698431365
transform 1 0 21504 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_187
timestamp 1698431365
transform 1 0 22288 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_203
timestamp 1698431365
transform 1 0 24080 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698431365
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_244
timestamp 1698431365
transform 1 0 28672 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_264
timestamp 1698431365
transform 1 0 30912 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_286
timestamp 1698431365
transform 1 0 33376 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_318
timestamp 1698431365
transform 1 0 36960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_320
timestamp 1698431365
transform 1 0 37184 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_325
timestamp 1698431365
transform 1 0 37744 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_341
timestamp 1698431365
transform 1 0 39536 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_67
timestamp 1698431365
transform 1 0 8848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_71
timestamp 1698431365
transform 1 0 9296 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_79
timestamp 1698431365
transform 1 0 10192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_86
timestamp 1698431365
transform 1 0 10976 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_94
timestamp 1698431365
transform 1 0 11872 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_123
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_181
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_197
timestamp 1698431365
transform 1 0 23408 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_205
timestamp 1698431365
transform 1 0 24304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_207
timestamp 1698431365
transform 1 0 24528 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_231
timestamp 1698431365
transform 1 0 27216 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_239
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_284
timestamp 1698431365
transform 1 0 33152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_321
timestamp 1698431365
transform 1 0 37296 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_337
timestamp 1698431365
transform 1 0 39088 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_345
timestamp 1698431365
transform 1 0 39984 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_377
timestamp 1698431365
transform 1 0 43568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_383
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_18
timestamp 1698431365
transform 1 0 3360 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_26
timestamp 1698431365
transform 1 0 4256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_30
timestamp 1698431365
transform 1 0 4704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_34
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_134
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_151
timestamp 1698431365
transform 1 0 18256 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_159
timestamp 1698431365
transform 1 0 19152 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_169
timestamp 1698431365
transform 1 0 20272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_173
timestamp 1698431365
transform 1 0 20720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_177
timestamp 1698431365
transform 1 0 21168 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_191
timestamp 1698431365
transform 1 0 22736 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_195
timestamp 1698431365
transform 1 0 23184 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_203
timestamp 1698431365
transform 1 0 24080 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698431365
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_228
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_232
timestamp 1698431365
transform 1 0 27328 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_332
timestamp 1698431365
transform 1 0 38528 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_43
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_54
timestamp 1698431365
transform 1 0 7392 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_86
timestamp 1698431365
transform 1 0 10976 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_102
timestamp 1698431365
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_139
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_157
timestamp 1698431365
transform 1 0 18928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_161
timestamp 1698431365
transform 1 0 19376 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_169
timestamp 1698431365
transform 1 0 20272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_193
timestamp 1698431365
transform 1 0 22960 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_197
timestamp 1698431365
transform 1 0 23408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_234
timestamp 1698431365
transform 1 0 27552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_238
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_327
timestamp 1698431365
transform 1 0 37968 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_343
timestamp 1698431365
transform 1 0 39760 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_360
timestamp 1698431365
transform 1 0 41664 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_376
timestamp 1698431365
transform 1 0 43456 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_26
timestamp 1698431365
transform 1 0 4256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_30
timestamp 1698431365
transform 1 0 4704 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_62
timestamp 1698431365
transform 1 0 8288 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_78
timestamp 1698431365
transform 1 0 10080 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_86
timestamp 1698431365
transform 1 0 10976 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_96
timestamp 1698431365
transform 1 0 12096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_100
timestamp 1698431365
transform 1 0 12544 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_122
timestamp 1698431365
transform 1 0 15008 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_158
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_197
timestamp 1698431365
transform 1 0 23408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_201
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_244
timestamp 1698431365
transform 1 0 28672 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_252
timestamp 1698431365
transform 1 0 29568 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_259
timestamp 1698431365
transform 1 0 30352 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_275
timestamp 1698431365
transform 1 0 32144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_318
timestamp 1698431365
transform 1 0 36960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_322
timestamp 1698431365
transform 1 0 37408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_338
timestamp 1698431365
transform 1 0 39200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_362
timestamp 1698431365
transform 1 0 41888 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_378
timestamp 1698431365
transform 1 0 43680 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_382
timestamp 1698431365
transform 1 0 44128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_47
timestamp 1698431365
transform 1 0 6608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_51
timestamp 1698431365
transform 1 0 7056 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_83
timestamp 1698431365
transform 1 0 10640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_85
timestamp 1698431365
transform 1 0 10864 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_92
timestamp 1698431365
transform 1 0 11648 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_100
timestamp 1698431365
transform 1 0 12544 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_109
timestamp 1698431365
transform 1 0 13552 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_116
timestamp 1698431365
transform 1 0 14336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_120
timestamp 1698431365
transform 1 0 14784 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_152
timestamp 1698431365
transform 1 0 18368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_158
timestamp 1698431365
transform 1 0 19040 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_279
timestamp 1698431365
transform 1 0 32592 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_295
timestamp 1698431365
transform 1 0 34384 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_303
timestamp 1698431365
transform 1 0 35280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_305
timestamp 1698431365
transform 1 0 35504 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698431365
transform 1 0 36400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_333
timestamp 1698431365
transform 1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_343
timestamp 1698431365
transform 1 0 39760 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_351
timestamp 1698431365
transform 1 0 40656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_355
timestamp 1698431365
transform 1 0 41104 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_369
timestamp 1698431365
transform 1 0 42672 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_377
timestamp 1698431365
transform 1 0 43568 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_381
timestamp 1698431365
transform 1 0 44016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_105
timestamp 1698431365
transform 1 0 13104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_107
timestamp 1698431365
transform 1 0 13328 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698431365
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_167
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_177
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_193
timestamp 1698431365
transform 1 0 22960 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_197
timestamp 1698431365
transform 1 0 23408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_204
timestamp 1698431365
transform 1 0 24192 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_330
timestamp 1698431365
transform 1 0 38304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_334
timestamp 1698431365
transform 1 0 38752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_336
timestamp 1698431365
transform 1 0 38976 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_345
timestamp 1698431365
transform 1 0 39984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_383
timestamp 1698431365
transform 1 0 44240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_69
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_77
timestamp 1698431365
transform 1 0 9968 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_87
timestamp 1698431365
transform 1 0 11088 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_103
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_111
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_121
timestamp 1698431365
transform 1 0 14896 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_153
timestamp 1698431365
transform 1 0 18480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_161
timestamp 1698431365
transform 1 0 19376 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_165
timestamp 1698431365
transform 1 0 19824 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698431365
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_197
timestamp 1698431365
transform 1 0 23408 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_201
timestamp 1698431365
transform 1 0 23856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_217
timestamp 1698431365
transform 1 0 25648 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_225
timestamp 1698431365
transform 1 0 26544 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_234
timestamp 1698431365
transform 1 0 27552 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_251
timestamp 1698431365
transform 1 0 29456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_253
timestamp 1698431365
transform 1 0 29680 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_262
timestamp 1698431365
transform 1 0 30688 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_270
timestamp 1698431365
transform 1 0 31584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_280
timestamp 1698431365
transform 1 0 32704 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_296
timestamp 1698431365
transform 1 0 34496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_300
timestamp 1698431365
transform 1 0 34944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_349
timestamp 1698431365
transform 1 0 40432 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_357
timestamp 1698431365
transform 1 0 41328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_364
timestamp 1698431365
transform 1 0 42112 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_380
timestamp 1698431365
transform 1 0 43904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_34
timestamp 1698431365
transform 1 0 5152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_38
timestamp 1698431365
transform 1 0 5600 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_120
timestamp 1698431365
transform 1 0 14784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_122
timestamp 1698431365
transform 1 0 15008 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_132
timestamp 1698431365
transform 1 0 16128 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_174
timestamp 1698431365
transform 1 0 20832 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_182
timestamp 1698431365
transform 1 0 21728 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_185
timestamp 1698431365
transform 1 0 22064 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_201
timestamp 1698431365
transform 1 0 23856 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_242
timestamp 1698431365
transform 1 0 28448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_246
timestamp 1698431365
transform 1 0 28896 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_286
timestamp 1698431365
transform 1 0 33376 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_306
timestamp 1698431365
transform 1 0 35616 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_338
timestamp 1698431365
transform 1 0 39200 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_18
timestamp 1698431365
transform 1 0 3360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_20
timestamp 1698431365
transform 1 0 3584 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_27
timestamp 1698431365
transform 1 0 4368 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_46
timestamp 1698431365
transform 1 0 6496 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_54
timestamp 1698431365
transform 1 0 7392 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_58
timestamp 1698431365
transform 1 0 7840 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_92
timestamp 1698431365
transform 1 0 11648 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_100
timestamp 1698431365
transform 1 0 12544 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698431365
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_139
timestamp 1698431365
transform 1 0 16912 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_143
timestamp 1698431365
transform 1 0 17360 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_155
timestamp 1698431365
transform 1 0 18704 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_168
timestamp 1698431365
transform 1 0 20160 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_184
timestamp 1698431365
transform 1 0 21952 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_235
timestamp 1698431365
transform 1 0 27664 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_279
timestamp 1698431365
transform 1 0 32592 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_283
timestamp 1698431365
transform 1 0 33040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_285
timestamp 1698431365
transform 1 0 33264 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_353
timestamp 1698431365
transform 1 0 40880 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_369
timestamp 1698431365
transform 1 0 42672 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_377
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_383
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_46
timestamp 1698431365
transform 1 0 6496 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_54
timestamp 1698431365
transform 1 0 7392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_56
timestamp 1698431365
transform 1 0 7616 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_63
timestamp 1698431365
transform 1 0 8400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_67
timestamp 1698431365
transform 1 0 8848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_100
timestamp 1698431365
transform 1 0 12544 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_132
timestamp 1698431365
transform 1 0 16128 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_165
timestamp 1698431365
transform 1 0 19824 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_197
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698431365
transform 1 0 24304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_228
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_232
timestamp 1698431365
transform 1 0 27328 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_245
timestamp 1698431365
transform 1 0 28784 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_261
timestamp 1698431365
transform 1 0 30576 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_274
timestamp 1698431365
transform 1 0 32032 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_298
timestamp 1698431365
transform 1 0 34720 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_302
timestamp 1698431365
transform 1 0 35168 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_315
timestamp 1698431365
transform 1 0 36624 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_331
timestamp 1698431365
transform 1 0 38416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_335
timestamp 1698431365
transform 1 0 38864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_337
timestamp 1698431365
transform 1 0 39088 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_18
timestamp 1698431365
transform 1 0 3360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_53
timestamp 1698431365
transform 1 0 7280 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_61
timestamp 1698431365
transform 1 0 8176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_65
timestamp 1698431365
transform 1 0 8624 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_73
timestamp 1698431365
transform 1 0 9520 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_77
timestamp 1698431365
transform 1 0 9968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_79
timestamp 1698431365
transform 1 0 10192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_92
timestamp 1698431365
transform 1 0 11648 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_100
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_113
timestamp 1698431365
transform 1 0 14000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_117
timestamp 1698431365
transform 1 0 14448 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_125
timestamp 1698431365
transform 1 0 15344 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_129
timestamp 1698431365
transform 1 0 15792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_144
timestamp 1698431365
transform 1 0 17472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_148
timestamp 1698431365
transform 1 0 17920 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_164
timestamp 1698431365
transform 1 0 19712 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_207
timestamp 1698431365
transform 1 0 24528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_211
timestamp 1698431365
transform 1 0 24976 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_331
timestamp 1698431365
transform 1 0 38416 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_368
timestamp 1698431365
transform 1 0 42560 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_34
timestamp 1698431365
transform 1 0 5152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_49
timestamp 1698431365
transform 1 0 6832 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_104
timestamp 1698431365
transform 1 0 12992 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_120
timestamp 1698431365
transform 1 0 14784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_122
timestamp 1698431365
transform 1 0 15008 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_236
timestamp 1698431365
transform 1 0 27776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_240
timestamp 1698431365
transform 1 0 28224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_253
timestamp 1698431365
transform 1 0 29680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_257
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_265
timestamp 1698431365
transform 1 0 31024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698431365
transform 1 0 31920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_298
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_302
timestamp 1698431365
transform 1 0 35168 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_304
timestamp 1698431365
transform 1 0 35392 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_317
timestamp 1698431365
transform 1 0 36848 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_333
timestamp 1698431365
transform 1 0 38640 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_356
timestamp 1698431365
transform 1 0 41216 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_366
timestamp 1698431365
transform 1 0 42336 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_382
timestamp 1698431365
transform 1 0 44128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_22
timestamp 1698431365
transform 1 0 3808 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_29
timestamp 1698431365
transform 1 0 4592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_33
timestamp 1698431365
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_46
timestamp 1698431365
transform 1 0 6496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_55
timestamp 1698431365
transform 1 0 7504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_59
timestamp 1698431365
transform 1 0 7952 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_75
timestamp 1698431365
transform 1 0 9744 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_83
timestamp 1698431365
transform 1 0 10640 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_87
timestamp 1698431365
transform 1 0 11088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_89
timestamp 1698431365
transform 1 0 11312 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_92
timestamp 1698431365
transform 1 0 11648 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_100
timestamp 1698431365
transform 1 0 12544 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_139
timestamp 1698431365
transform 1 0 16912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_147
timestamp 1698431365
transform 1 0 17808 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_163
timestamp 1698431365
transform 1 0 19600 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_251
timestamp 1698431365
transform 1 0 29456 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_265
timestamp 1698431365
transform 1 0 31024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_269
timestamp 1698431365
transform 1 0 31472 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_301
timestamp 1698431365
transform 1 0 35056 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_330
timestamp 1698431365
transform 1 0 38304 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_346
timestamp 1698431365
transform 1 0 40096 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_383
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_32
timestamp 1698431365
transform 1 0 4928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_36
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_44
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_64
timestamp 1698431365
transform 1 0 8512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_80
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_82
timestamp 1698431365
transform 1 0 10528 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_103
timestamp 1698431365
transform 1 0 12880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_107
timestamp 1698431365
transform 1 0 13328 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_123
timestamp 1698431365
transform 1 0 15120 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_128
timestamp 1698431365
transform 1 0 15680 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_132
timestamp 1698431365
transform 1 0 16128 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_150
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_161
timestamp 1698431365
transform 1 0 19376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_165
timestamp 1698431365
transform 1 0 19824 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_181
timestamp 1698431365
transform 1 0 21616 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_189
timestamp 1698431365
transform 1 0 22512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_193
timestamp 1698431365
transform 1 0 22960 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_202
timestamp 1698431365
transform 1 0 23968 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_224
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_226
timestamp 1698431365
transform 1 0 26656 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_264
timestamp 1698431365
transform 1 0 30912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_308
timestamp 1698431365
transform 1 0 35840 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_340
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_49
timestamp 1698431365
transform 1 0 6832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_51
timestamp 1698431365
transform 1 0 7056 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_54
timestamp 1698431365
transform 1 0 7392 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_86
timestamp 1698431365
transform 1 0 10976 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_94
timestamp 1698431365
transform 1 0 11872 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_98
timestamp 1698431365
transform 1 0 12320 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_118
timestamp 1698431365
transform 1 0 14560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_122
timestamp 1698431365
transform 1 0 15008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_126
timestamp 1698431365
transform 1 0 15456 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_158
timestamp 1698431365
transform 1 0 19040 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_162
timestamp 1698431365
transform 1 0 19488 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_165
timestamp 1698431365
transform 1 0 19824 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_189
timestamp 1698431365
transform 1 0 22512 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_205
timestamp 1698431365
transform 1 0 24304 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_213
timestamp 1698431365
transform 1 0 25200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_221
timestamp 1698431365
transform 1 0 26096 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_237
timestamp 1698431365
transform 1 0 27888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_275
timestamp 1698431365
transform 1 0 32144 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_291
timestamp 1698431365
transform 1 0 33936 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_299
timestamp 1698431365
transform 1 0 34832 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_303
timestamp 1698431365
transform 1 0 35280 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_305
timestamp 1698431365
transform 1 0 35504 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_381
timestamp 1698431365
transform 1 0 44016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_383
timestamp 1698431365
transform 1 0 44240 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_104
timestamp 1698431365
transform 1 0 12992 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_123
timestamp 1698431365
transform 1 0 15120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_125
timestamp 1698431365
transform 1 0 15344 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_135
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_154
timestamp 1698431365
transform 1 0 18592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_192
timestamp 1698431365
transform 1 0 22848 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_218
timestamp 1698431365
transform 1 0 25760 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_222
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_254
timestamp 1698431365
transform 1 0 29792 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_270
timestamp 1698431365
transform 1 0 31584 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_278
timestamp 1698431365
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_327
timestamp 1698431365
transform 1 0 37968 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_331
timestamp 1698431365
transform 1 0 38416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_341
timestamp 1698431365
transform 1 0 39536 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_50
timestamp 1698431365
transform 1 0 6944 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_66
timestamp 1698431365
transform 1 0 8736 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_86
timestamp 1698431365
transform 1 0 10976 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_102
timestamp 1698431365
transform 1 0 12768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_139
timestamp 1698431365
transform 1 0 16912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_143
timestamp 1698431365
transform 1 0 17360 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_159
timestamp 1698431365
transform 1 0 19152 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_163
timestamp 1698431365
transform 1 0 19600 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_279
timestamp 1698431365
transform 1 0 32592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_281
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_284
timestamp 1698431365
transform 1 0 33152 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_290
timestamp 1698431365
transform 1 0 33824 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_306
timestamp 1698431365
transform 1 0 35616 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_330
timestamp 1698431365
transform 1 0 38304 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_346
timestamp 1698431365
transform 1 0 40096 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_354
timestamp 1698431365
transform 1 0 40992 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_356
timestamp 1698431365
transform 1 0 41216 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_370
timestamp 1698431365
transform 1 0 42784 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_378
timestamp 1698431365
transform 1 0 43680 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_382
timestamp 1698431365
transform 1 0 44128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_32
timestamp 1698431365
transform 1 0 4928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_36
timestamp 1698431365
transform 1 0 5376 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_48
timestamp 1698431365
transform 1 0 6720 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_64
timestamp 1698431365
transform 1 0 8512 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_83
timestamp 1698431365
transform 1 0 10640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_90
timestamp 1698431365
transform 1 0 11424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_94
timestamp 1698431365
transform 1 0 11872 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_110
timestamp 1698431365
transform 1 0 13664 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_114
timestamp 1698431365
transform 1 0 14112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_137
timestamp 1698431365
transform 1 0 16688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_218
timestamp 1698431365
transform 1 0 25760 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_231
timestamp 1698431365
transform 1 0 27216 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_263
timestamp 1698431365
transform 1 0 30800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_340
timestamp 1698431365
transform 1 0 39424 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_381
timestamp 1698431365
transform 1 0 44016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_383
timestamp 1698431365
transform 1 0 44240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_93
timestamp 1698431365
transform 1 0 11760 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_97
timestamp 1698431365
transform 1 0 12208 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_109
timestamp 1698431365
transform 1 0 13552 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_114
timestamp 1698431365
transform 1 0 14112 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_135
timestamp 1698431365
transform 1 0 16464 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_168
timestamp 1698431365
transform 1 0 20160 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698431365
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_209
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_213
timestamp 1698431365
transform 1 0 25200 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_215
timestamp 1698431365
transform 1 0 25424 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_234
timestamp 1698431365
transform 1 0 27552 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_257
timestamp 1698431365
transform 1 0 30128 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_276
timestamp 1698431365
transform 1 0 32256 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_308
timestamp 1698431365
transform 1 0 35840 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_312
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_322
timestamp 1698431365
transform 1 0 37408 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_330
timestamp 1698431365
transform 1 0 38304 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_334
timestamp 1698431365
transform 1 0 38752 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_343
timestamp 1698431365
transform 1 0 39760 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_375
timestamp 1698431365
transform 1 0 43344 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_383
timestamp 1698431365
transform 1 0 44240 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_34
timestamp 1698431365
transform 1 0 5152 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_42
timestamp 1698431365
transform 1 0 6048 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_46
timestamp 1698431365
transform 1 0 6496 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_49
timestamp 1698431365
transform 1 0 6832 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_65
timestamp 1698431365
transform 1 0 8624 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_74
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_132
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_154
timestamp 1698431365
transform 1 0 18592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_170
timestamp 1698431365
transform 1 0 20384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_174
timestamp 1698431365
transform 1 0 20832 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_230
timestamp 1698431365
transform 1 0 27104 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_270
timestamp 1698431365
transform 1 0 31584 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_294
timestamp 1698431365
transform 1 0 34272 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_296
timestamp 1698431365
transform 1 0 34496 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_311
timestamp 1698431365
transform 1 0 36176 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_327
timestamp 1698431365
transform 1 0 37968 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_331
timestamp 1698431365
transform 1 0 38416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_341
timestamp 1698431365
transform 1 0 39536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_343
timestamp 1698431365
transform 1 0 39760 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_45
timestamp 1698431365
transform 1 0 6384 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_61
timestamp 1698431365
transform 1 0 8176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_73
timestamp 1698431365
transform 1 0 9520 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_81
timestamp 1698431365
transform 1 0 10416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_85
timestamp 1698431365
transform 1 0 10864 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_92
timestamp 1698431365
transform 1 0 11648 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_111
timestamp 1698431365
transform 1 0 13776 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_227
timestamp 1698431365
transform 1 0 26768 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_322
timestamp 1698431365
transform 1 0 37408 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_354
timestamp 1698431365
transform 1 0 40992 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_363
timestamp 1698431365
transform 1 0 42000 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_379
timestamp 1698431365
transform 1 0 43792 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_36
timestamp 1698431365
transform 1 0 5376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_40
timestamp 1698431365
transform 1 0 5824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_44
timestamp 1698431365
transform 1 0 6272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_62
timestamp 1698431365
transform 1 0 8288 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_92
timestamp 1698431365
transform 1 0 11648 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_106
timestamp 1698431365
transform 1 0 13216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_114
timestamp 1698431365
transform 1 0 14112 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_124
timestamp 1698431365
transform 1 0 15232 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_149
timestamp 1698431365
transform 1 0 18032 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_157
timestamp 1698431365
transform 1 0 18928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_159
timestamp 1698431365
transform 1 0 19152 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_170
timestamp 1698431365
transform 1 0 20384 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_178
timestamp 1698431365
transform 1 0 21280 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_192
timestamp 1698431365
transform 1 0 22848 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_208
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_222
timestamp 1698431365
transform 1 0 26208 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_254
timestamp 1698431365
transform 1 0 29792 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_258
timestamp 1698431365
transform 1 0 30240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_261
timestamp 1698431365
transform 1 0 30576 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_277
timestamp 1698431365
transform 1 0 32368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_286
timestamp 1698431365
transform 1 0 33376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_288
timestamp 1698431365
transform 1 0 33600 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_328
timestamp 1698431365
transform 1 0 38080 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_344
timestamp 1698431365
transform 1 0 39872 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_348
timestamp 1698431365
transform 1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_354
timestamp 1698431365
transform 1 0 40992 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_362
timestamp 1698431365
transform 1 0 41888 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_378
timestamp 1698431365
transform 1 0 43680 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_382
timestamp 1698431365
transform 1 0 44128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_59
timestamp 1698431365
transform 1 0 7952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_63
timestamp 1698431365
transform 1 0 8400 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_79
timestamp 1698431365
transform 1 0 10192 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_85
timestamp 1698431365
transform 1 0 10864 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_89
timestamp 1698431365
transform 1 0 11312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_91
timestamp 1698431365
transform 1 0 11536 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_100
timestamp 1698431365
transform 1 0 12544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_115
timestamp 1698431365
transform 1 0 14224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_128
timestamp 1698431365
transform 1 0 15680 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_136
timestamp 1698431365
transform 1 0 16576 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_142
timestamp 1698431365
transform 1 0 17248 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_209
timestamp 1698431365
transform 1 0 24752 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_213
timestamp 1698431365
transform 1 0 25200 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_227
timestamp 1698431365
transform 1 0 26768 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_243
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_279
timestamp 1698431365
transform 1 0 32592 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_295
timestamp 1698431365
transform 1 0 34384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_299
timestamp 1698431365
transform 1 0 34832 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_303
timestamp 1698431365
transform 1 0 35280 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_305
timestamp 1698431365
transform 1 0 35504 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_333
timestamp 1698431365
transform 1 0 38640 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_341
timestamp 1698431365
transform 1 0 39536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_383
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_34
timestamp 1698431365
transform 1 0 5152 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_50
timestamp 1698431365
transform 1 0 6944 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_58
timestamp 1698431365
transform 1 0 7840 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_62
timestamp 1698431365
transform 1 0 8288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_97
timestamp 1698431365
transform 1 0 12208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_101
timestamp 1698431365
transform 1 0 12656 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_117
timestamp 1698431365
transform 1 0 14448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_121
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_123
timestamp 1698431365
transform 1 0 15120 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_132
timestamp 1698431365
transform 1 0 16128 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_158
timestamp 1698431365
transform 1 0 19040 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_166
timestamp 1698431365
transform 1 0 19936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_170
timestamp 1698431365
transform 1 0 20384 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_179
timestamp 1698431365
transform 1 0 21392 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_183
timestamp 1698431365
transform 1 0 21840 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_204
timestamp 1698431365
transform 1 0 24192 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_220
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_252
timestamp 1698431365
transform 1 0 29568 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_255
timestamp 1698431365
transform 1 0 29904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_259
timestamp 1698431365
transform 1 0 30352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_275
timestamp 1698431365
transform 1 0 32144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_41
timestamp 1698431365
transform 1 0 5936 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_49
timestamp 1698431365
transform 1 0 6832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_80
timestamp 1698431365
transform 1 0 10304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_84
timestamp 1698431365
transform 1 0 10752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_88
timestamp 1698431365
transform 1 0 11200 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_109
timestamp 1698431365
transform 1 0 13552 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_139
timestamp 1698431365
transform 1 0 16912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_143
timestamp 1698431365
transform 1 0 17360 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_159
timestamp 1698431365
transform 1 0 19152 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_182
timestamp 1698431365
transform 1 0 21728 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_198
timestamp 1698431365
transform 1 0 23520 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_202
timestamp 1698431365
transform 1 0 23968 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_288
timestamp 1698431365
transform 1 0 33600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_292
timestamp 1698431365
transform 1 0 34048 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_308
timestamp 1698431365
transform 1 0 35840 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_322
timestamp 1698431365
transform 1 0 37408 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_338
timestamp 1698431365
transform 1 0 39200 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_346
timestamp 1698431365
transform 1 0 40096 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_353
timestamp 1698431365
transform 1 0 40880 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_369
timestamp 1698431365
transform 1 0 42672 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_377
timestamp 1698431365
transform 1 0 43568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_74
timestamp 1698431365
transform 1 0 9632 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_77
timestamp 1698431365
transform 1 0 9968 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_109
timestamp 1698431365
transform 1 0 13552 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_125
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_133
timestamp 1698431365
transform 1 0 16240 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_137
timestamp 1698431365
transform 1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_158
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_162
timestamp 1698431365
transform 1 0 19488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_170
timestamp 1698431365
transform 1 0 20384 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_186
timestamp 1698431365
transform 1 0 22176 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_194
timestamp 1698431365
transform 1 0 23072 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_196
timestamp 1698431365
transform 1 0 23296 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_228
timestamp 1698431365
transform 1 0 26880 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_232
timestamp 1698431365
transform 1 0 27328 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_262
timestamp 1698431365
transform 1 0 30688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_266
timestamp 1698431365
transform 1 0 31136 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_274
timestamp 1698431365
transform 1 0 32032 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_278
timestamp 1698431365
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_288
timestamp 1698431365
transform 1 0 33600 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_326
timestamp 1698431365
transform 1 0 37856 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_330
timestamp 1698431365
transform 1 0 38304 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_338
timestamp 1698431365
transform 1 0 39200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_381
timestamp 1698431365
transform 1 0 44016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_383
timestamp 1698431365
transform 1 0 44240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_49
timestamp 1698431365
transform 1 0 6832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_67
timestamp 1698431365
transform 1 0 8848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_99
timestamp 1698431365
transform 1 0 12432 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_103
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_139
timestamp 1698431365
transform 1 0 16912 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_155
timestamp 1698431365
transform 1 0 18704 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_163
timestamp 1698431365
transform 1 0 19600 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_217
timestamp 1698431365
transform 1 0 25648 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_233
timestamp 1698431365
transform 1 0 27440 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_328
timestamp 1698431365
transform 1 0 38080 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_344
timestamp 1698431365
transform 1 0 39872 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_348
timestamp 1698431365
transform 1 0 40320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_355
timestamp 1698431365
transform 1 0 41104 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_371
timestamp 1698431365
transform 1 0 42896 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_379
timestamp 1698431365
transform 1 0 43792 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_383
timestamp 1698431365
transform 1 0 44240 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_18
timestamp 1698431365
transform 1 0 3360 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_36
timestamp 1698431365
transform 1 0 5376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_40
timestamp 1698431365
transform 1 0 5824 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_56
timestamp 1698431365
transform 1 0 7616 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_64
timestamp 1698431365
transform 1 0 8512 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_80
timestamp 1698431365
transform 1 0 10304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_113
timestamp 1698431365
transform 1 0 14000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_117
timestamp 1698431365
transform 1 0 14448 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_133
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_158
timestamp 1698431365
transform 1 0 19040 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_166
timestamp 1698431365
transform 1 0 19936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698431365
transform 1 0 20160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_175
timestamp 1698431365
transform 1 0 20944 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_191
timestamp 1698431365
transform 1 0 22736 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_199
timestamp 1698431365
transform 1 0 23632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_201
timestamp 1698431365
transform 1 0 23856 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_204
timestamp 1698431365
transform 1 0 24192 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_220
timestamp 1698431365
transform 1 0 25984 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_252
timestamp 1698431365
transform 1 0 29568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_268
timestamp 1698431365
transform 1 0 31360 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_358
timestamp 1698431365
transform 1 0 41440 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_374
timestamp 1698431365
transform 1 0 43232 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_382
timestamp 1698431365
transform 1 0 44128 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_41
timestamp 1698431365
transform 1 0 5936 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_49
timestamp 1698431365
transform 1 0 6832 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_53
timestamp 1698431365
transform 1 0 7280 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_55
timestamp 1698431365
transform 1 0 7504 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_85
timestamp 1698431365
transform 1 0 10864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_89
timestamp 1698431365
transform 1 0 11312 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_123
timestamp 1698431365
transform 1 0 15120 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_127
timestamp 1698431365
transform 1 0 15568 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_157
timestamp 1698431365
transform 1 0 18928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_161
timestamp 1698431365
transform 1 0 19376 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_193
timestamp 1698431365
transform 1 0 22960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_195
timestamp 1698431365
transform 1 0 23184 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_223
timestamp 1698431365
transform 1 0 26320 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_227
timestamp 1698431365
transform 1 0 26768 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_243
timestamp 1698431365
transform 1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_323
timestamp 1698431365
transform 1 0 37520 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_339
timestamp 1698431365
transform 1 0 39312 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_343
timestamp 1698431365
transform 1 0 39760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_345
timestamp 1698431365
transform 1 0 39984 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_351
timestamp 1698431365
transform 1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_358
timestamp 1698431365
transform 1 0 41440 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_374
timestamp 1698431365
transform 1 0 43232 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_382
timestamp 1698431365
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_158
timestamp 1698431365
transform 1 0 19040 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_166
timestamp 1698431365
transform 1 0 19936 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_172
timestamp 1698431365
transform 1 0 20608 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_188
timestamp 1698431365
transform 1 0 22400 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_196
timestamp 1698431365
transform 1 0 23296 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_214
timestamp 1698431365
transform 1 0 25312 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_233
timestamp 1698431365
transform 1 0 27440 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_265
timestamp 1698431365
transform 1 0 31024 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_273
timestamp 1698431365
transform 1 0 31920 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_277
timestamp 1698431365
transform 1 0 32368 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_279
timestamp 1698431365
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_290
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_294
timestamp 1698431365
transform 1 0 34272 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_332
timestamp 1698431365
transform 1 0 38528 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_336
timestamp 1698431365
transform 1 0 38976 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_340
timestamp 1698431365
transform 1 0 39424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_347
timestamp 1698431365
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_349
timestamp 1698431365
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_366
timestamp 1698431365
transform 1 0 42336 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_382
timestamp 1698431365
transform 1 0 44128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698431365
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_41
timestamp 1698431365
transform 1 0 5936 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_57
timestamp 1698431365
transform 1 0 7728 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_69
timestamp 1698431365
transform 1 0 9072 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_123
timestamp 1698431365
transform 1 0 15120 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_131
timestamp 1698431365
transform 1 0 16016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_133
timestamp 1698431365
transform 1 0 16240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_136
timestamp 1698431365
transform 1 0 16576 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_144
timestamp 1698431365
transform 1 0 17472 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_193
timestamp 1698431365
transform 1 0 22960 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_226
timestamp 1698431365
transform 1 0 26656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_230
timestamp 1698431365
transform 1 0 27104 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_238
timestamp 1698431365
transform 1 0 28000 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_251
timestamp 1698431365
transform 1 0 29456 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_281
timestamp 1698431365
transform 1 0 32816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_285
timestamp 1698431365
transform 1 0 33264 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_301
timestamp 1698431365
transform 1 0 35056 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_309
timestamp 1698431365
transform 1 0 35952 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_313
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_333
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_366
timestamp 1698431365
transform 1 0 42336 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_18
timestamp 1698431365
transform 1 0 3360 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_26
timestamp 1698431365
transform 1 0 4256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_59
timestamp 1698431365
transform 1 0 7952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_63
timestamp 1698431365
transform 1 0 8400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_67
timestamp 1698431365
transform 1 0 8848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_69
timestamp 1698431365
transform 1 0 9072 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_103
timestamp 1698431365
transform 1 0 12880 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_134
timestamp 1698431365
transform 1 0 16352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_173
timestamp 1698431365
transform 1 0 20720 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_189
timestamp 1698431365
transform 1 0 22512 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_197
timestamp 1698431365
transform 1 0 23408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_207
timestamp 1698431365
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_232
timestamp 1698431365
transform 1 0 27328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_263
timestamp 1698431365
transform 1 0 30800 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_267
timestamp 1698431365
transform 1 0 31248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_275
timestamp 1698431365
transform 1 0 32144 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_311
timestamp 1698431365
transform 1 0 36176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_315
timestamp 1698431365
transform 1 0 36624 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_347
timestamp 1698431365
transform 1 0 40208 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_382
timestamp 1698431365
transform 1 0 44128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_349
timestamp 1698431365
transform 1 0 40432 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_357
timestamp 1698431365
transform 1 0 41328 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_26
timestamp 1698431365
transform 1 0 4256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_30
timestamp 1698431365
transform 1 0 4704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_36
timestamp 1698431365
transform 1 0 5376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_38
timestamp 1698431365
transform 1 0 5600 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_45
timestamp 1698431365
transform 1 0 6384 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_61
timestamp 1698431365
transform 1 0 8176 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_65
timestamp 1698431365
transform 1 0 8624 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_70
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_79
timestamp 1698431365
transform 1 0 10192 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_95
timestamp 1698431365
transform 1 0 11984 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_99
timestamp 1698431365
transform 1 0 12432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_101
timestamp 1698431365
transform 1 0 12656 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_106
timestamp 1698431365
transform 1 0 13216 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_133
timestamp 1698431365
transform 1 0 16240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_135
timestamp 1698431365
transform 1 0 16464 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_138
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_140
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_167
timestamp 1698431365
transform 1 0 20048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_169
timestamp 1698431365
transform 1 0 20272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_174
timestamp 1698431365
transform 1 0 20832 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_201
timestamp 1698431365
transform 1 0 23856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_203
timestamp 1698431365
transform 1 0 24080 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_208
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_235
timestamp 1698431365
transform 1 0 27664 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_237
timestamp 1698431365
transform 1 0 27888 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_240
timestamp 1698431365
transform 1 0 28224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_242
timestamp 1698431365
transform 1 0 28448 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_269
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_271
timestamp 1698431365
transform 1 0 31696 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_274
timestamp 1698431365
transform 1 0 32032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_303
timestamp 1698431365
transform 1 0 35280 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_305
timestamp 1698431365
transform 1 0 35504 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_308
timestamp 1698431365
transform 1 0 35840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_310
timestamp 1698431365
transform 1 0 36064 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_337
timestamp 1698431365
transform 1 0 39088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_339
timestamp 1698431365
transform 1 0 39312 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_342
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_344
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_371
timestamp 1698431365
transform 1 0 42896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_373
timestamp 1698431365
transform 1 0 43120 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_376
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 9520 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 5712 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698431365
transform 1 0 17136 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698431365
transform 1 0 20944 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698431365
transform -1 0 31472 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698431365
transform 1 0 36176 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698431365
transform 1 0 39984 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform 1 0 41440 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_50 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 44576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 44576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 44576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 44576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 44576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 44576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 44576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 44576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 44576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 44576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 44576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 44576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 44576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 44576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 44576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 44576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 44576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 44576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 44576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 44576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 44576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 44576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 44576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 44576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 44576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 44576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 44576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 44576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 44576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 44576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 44576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 44576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 44576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 44576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 44576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 44576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 44576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 44576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 44576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 44576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 44576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 44576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 44576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_112
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_113
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_114
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_115
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_118
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_119
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_120
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_121
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_122
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_123
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_124
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_125
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_126
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_127
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_128
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_129
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_130
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_131
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_132
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_133
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_134
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_135
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_136
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_137
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_138
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_139
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_140
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_141
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_142
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_143
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_144
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_145
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_146
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_147
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_148
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_149
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_150
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_151
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_152
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_153
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_154
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_155
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_156
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_157
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_158
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_159
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_160
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_161
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_162
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_163
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_164
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_165
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_166
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_167
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_168
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_169
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_170
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_171
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_172
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_173
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_174
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_175
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_176
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_177
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_178
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_179
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_180
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_181
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_182
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_183
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_184
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_185
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_186
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_187
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_188
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_189
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_190
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_191
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_192
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_193
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_194
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_195
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_196
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_197
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_198
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_199
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_200
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_201
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_202
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_209
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_210
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_212
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_213
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_214
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_215
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_216
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_217
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_218
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_219
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_220
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_221
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_222
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_223
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_224
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_225
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_226
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_227
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_228
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_229
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_230
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_231
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_232
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_233
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_234
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_235
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_236
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_237
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_238
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_239
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_240
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_241
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_242
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_243
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_244
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_245
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_246
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_247
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_248
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_249
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_250
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_251
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_252
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_253
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_254
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_255
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_256
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_257
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_258
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_259
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_260
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_261
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_262
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_263
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_264
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_265
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_266
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_267
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_268
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_269
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_270
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_271
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_272
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_273
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_274
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_275
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_276
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_277
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_278
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_279
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_280
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_281
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_282
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_283
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_284
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_285
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_286
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_287
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_288
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_289
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_290
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_291
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_292
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_293
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_294
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_295
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_296
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_297
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_298
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_299
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_300
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_301
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_302
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_303
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_304
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_305
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_306
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_307
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_308
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_309
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_310
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_311
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_312
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_313
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_314
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_315
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_316
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_317
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_318
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_319
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_320
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_321
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_322
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_323
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_324
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_325
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_326
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_327
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_328
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_329
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_330
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_331
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_332
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_333
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_334
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_335
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_336
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_337
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_338
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_339
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_340
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_341
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_342
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_343
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_344
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_345
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_346
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_347
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_348
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_349
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_350
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_351
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_352
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_353
timestamp 1698431365
transform 1 0 12768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_354
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_355
timestamp 1698431365
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_356
timestamp 1698431365
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_357
timestamp 1698431365
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_358
timestamp 1698431365
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_359
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_360
timestamp 1698431365
transform 1 0 39424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_361
timestamp 1698431365
transform 1 0 43232 0 -1 42336
box -86 -86 310 870
<< labels >>
flabel metal2 s 9408 45200 9520 46000 0 FreeSans 448 90 0 0 io_in
port 0 nsew signal input
flabel metal2 s 13216 45200 13328 46000 0 FreeSans 448 90 0 0 io_out[0]
port 1 nsew signal tristate
flabel metal2 s 17024 45200 17136 46000 0 FreeSans 448 90 0 0 io_out[1]
port 2 nsew signal tristate
flabel metal2 s 20832 45200 20944 46000 0 FreeSans 448 90 0 0 io_out[2]
port 3 nsew signal tristate
flabel metal2 s 24640 45200 24752 46000 0 FreeSans 448 90 0 0 io_out[3]
port 4 nsew signal tristate
flabel metal2 s 28448 45200 28560 46000 0 FreeSans 448 90 0 0 io_out[4]
port 5 nsew signal tristate
flabel metal2 s 32256 45200 32368 46000 0 FreeSans 448 90 0 0 io_out[5]
port 6 nsew signal tristate
flabel metal2 s 36064 45200 36176 46000 0 FreeSans 448 90 0 0 io_out[6]
port 7 nsew signal tristate
flabel metal2 s 39872 45200 39984 46000 0 FreeSans 448 90 0 0 io_out[7]
port 8 nsew signal tristate
flabel metal2 s 43680 45200 43792 46000 0 FreeSans 448 90 0 0 io_out[8]
port 9 nsew signal tristate
flabel metal2 s 5600 45200 5712 46000 0 FreeSans 448 90 0 0 rst_n
port 10 nsew signal input
flabel metal4 s 4448 3076 4768 42396 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 35168 3076 35488 42396 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 19808 3076 20128 42396 0 FreeSans 1280 90 0 0 vss
port 12 nsew ground bidirectional
flabel metal2 s 1792 45200 1904 46000 0 FreeSans 448 90 0 0 wb_clk_i
port 13 nsew signal input
rlabel metal1 22960 41552 22960 41552 0 vdd
rlabel metal1 22960 42336 22960 42336 0 vss
rlabel metal2 18984 39984 18984 39984 0 _000_
rlabel metal2 25704 39984 25704 39984 0 _001_
rlabel metal2 25816 39704 25816 39704 0 _002_
rlabel metal2 23632 38136 23632 38136 0 _003_
rlabel metal2 33880 39648 33880 39648 0 _004_
rlabel metal2 14616 39872 14616 39872 0 _005_
rlabel metal2 18424 39984 18424 39984 0 _006_
rlabel metal2 20664 14504 20664 14504 0 _007_
rlabel metal2 25032 13272 25032 13272 0 _008_
rlabel metal2 27832 4424 27832 4424 0 _009_
rlabel metal2 22456 4760 22456 4760 0 _010_
rlabel metal2 22848 8904 22848 8904 0 _011_
rlabel metal3 30800 8344 30800 8344 0 _012_
rlabel metal2 35224 12488 35224 12488 0 _013_
rlabel metal2 28840 12544 28840 12544 0 _014_
rlabel metal2 31304 17640 31304 17640 0 _015_
rlabel metal3 24640 17528 24640 17528 0 _016_
rlabel metal3 28504 38808 28504 38808 0 _017_
rlabel metal2 20216 38136 20216 38136 0 _018_
rlabel metal2 20440 38472 20440 38472 0 _019_
rlabel metal2 37072 27944 37072 27944 0 _020_
rlabel metal2 35896 31388 35896 31388 0 _021_
rlabel metal3 36624 35560 36624 35560 0 _022_
rlabel metal2 41832 39480 41832 39480 0 _023_
rlabel metal2 41496 39256 41496 39256 0 _024_
rlabel metal3 40992 35560 40992 35560 0 _025_
rlabel metal2 36792 38640 36792 38640 0 _026_
rlabel metal2 41832 32984 41832 32984 0 _027_
rlabel metal2 41944 29008 41944 29008 0 _028_
rlabel metal2 41888 19320 41888 19320 0 _029_
rlabel metal2 34328 16800 34328 16800 0 _030_
rlabel metal2 41272 16800 41272 16800 0 _031_
rlabel metal2 38136 14840 38136 14840 0 _032_
rlabel metal3 34832 21784 34832 21784 0 _033_
rlabel metal2 41888 24920 41888 24920 0 _034_
rlabel metal2 39648 23352 39648 23352 0 _035_
rlabel metal2 15960 15624 15960 15624 0 _036_
rlabel metal3 21728 18424 21728 18424 0 _037_
rlabel metal2 21784 23184 21784 23184 0 _038_
rlabel metal2 14392 20496 14392 20496 0 _039_
rlabel metal2 10584 20496 10584 20496 0 _040_
rlabel metal3 3192 26936 3192 26936 0 _041_
rlabel metal2 2632 21896 2632 21896 0 _042_
rlabel metal2 4088 25928 4088 25928 0 _043_
rlabel metal2 2632 17976 2632 17976 0 _044_
rlabel metal2 2744 15624 2744 15624 0 _045_
rlabel metal2 4536 9352 4536 9352 0 _046_
rlabel metal3 5152 12264 5152 12264 0 _047_
rlabel metal2 10752 6776 10752 6776 0 _048_
rlabel metal2 12768 5992 12768 5992 0 _049_
rlabel metal2 17976 11760 17976 11760 0 _050_
rlabel metal2 19544 7784 19544 7784 0 _051_
rlabel metal3 3640 37464 3640 37464 0 _052_
rlabel metal2 5096 37688 5096 37688 0 _053_
rlabel metal3 19768 27720 19768 27720 0 _054_
rlabel metal2 15624 34384 15624 34384 0 _055_
rlabel metal2 11928 34384 11928 34384 0 _056_
rlabel metal2 7000 33656 7000 33656 0 _057_
rlabel metal2 10920 35112 10920 35112 0 _058_
rlabel metal3 5040 32424 5040 32424 0 _059_
rlabel metal2 30296 21168 30296 21168 0 _060_
rlabel metal3 28504 24920 28504 24920 0 _061_
rlabel metal2 27048 21224 27048 21224 0 _062_
rlabel metal2 32088 34552 32088 34552 0 _063_
rlabel metal2 30184 31528 30184 31528 0 _064_
rlabel metal2 29792 31528 29792 31528 0 _065_
rlabel metal2 31752 30968 31752 30968 0 _066_
rlabel metal2 29904 30968 29904 30968 0 _067_
rlabel metal3 26320 30968 26320 30968 0 _068_
rlabel metal2 26208 30184 26208 30184 0 _069_
rlabel metal3 24192 32424 24192 32424 0 _070_
rlabel metal2 19768 30576 19768 30576 0 _071_
rlabel metal3 18144 30968 18144 30968 0 _072_
rlabel metal3 6552 31864 6552 31864 0 _073_
rlabel metal2 7896 32816 7896 32816 0 _074_
rlabel metal2 19096 31248 19096 31248 0 _075_
rlabel metal2 26824 15904 26824 15904 0 _076_
rlabel metal3 25144 13496 25144 13496 0 _077_
rlabel metal2 27552 7672 27552 7672 0 _078_
rlabel metal2 25256 29344 25256 29344 0 _079_
rlabel metal2 19600 30184 19600 30184 0 _080_
rlabel metal3 15400 27832 15400 27832 0 _081_
rlabel metal2 14056 27776 14056 27776 0 _082_
rlabel metal2 9800 29120 9800 29120 0 _083_
rlabel metal2 9464 29120 9464 29120 0 _084_
rlabel metal2 10024 28616 10024 28616 0 _085_
rlabel metal2 13944 28504 13944 28504 0 _086_
rlabel metal2 15400 26656 15400 26656 0 _087_
rlabel metal2 13832 27216 13832 27216 0 _088_
rlabel metal2 15064 28784 15064 28784 0 _089_
rlabel metal3 13160 28616 13160 28616 0 _090_
rlabel metal2 21336 27832 21336 27832 0 _091_
rlabel metal2 15512 29120 15512 29120 0 _092_
rlabel metal2 16632 29512 16632 29512 0 _093_
rlabel metal2 17304 25984 17304 25984 0 _094_
rlabel metal2 14728 29848 14728 29848 0 _095_
rlabel metal2 15960 29680 15960 29680 0 _096_
rlabel metal2 15904 28056 15904 28056 0 _097_
rlabel metal3 16856 26488 16856 26488 0 _098_
rlabel metal2 15960 27776 15960 27776 0 _099_
rlabel metal2 6328 29288 6328 29288 0 _100_
rlabel metal3 11256 30128 11256 30128 0 _101_
rlabel metal3 7952 30184 7952 30184 0 _102_
rlabel metal2 16520 29680 16520 29680 0 _103_
rlabel metal2 15288 29960 15288 29960 0 _104_
rlabel metal2 21112 33432 21112 33432 0 _105_
rlabel metal2 31416 23968 31416 23968 0 _106_
rlabel metal2 27384 29624 27384 29624 0 _107_
rlabel metal2 25592 30576 25592 30576 0 _108_
rlabel metal2 26712 31360 26712 31360 0 _109_
rlabel metal3 24640 33880 24640 33880 0 _110_
rlabel metal2 21672 32760 21672 32760 0 _111_
rlabel metal2 20440 35000 20440 35000 0 _112_
rlabel metal2 20216 35168 20216 35168 0 _113_
rlabel metal2 21336 34944 21336 34944 0 _114_
rlabel metal3 21000 37912 21000 37912 0 _115_
rlabel metal2 20216 39256 20216 39256 0 _116_
rlabel metal2 26600 33432 26600 33432 0 _117_
rlabel metal2 25648 31976 25648 31976 0 _118_
rlabel metal2 26320 30968 26320 30968 0 _119_
rlabel metal2 25928 32256 25928 32256 0 _120_
rlabel metal2 26488 33992 26488 33992 0 _121_
rlabel metal2 25816 37016 25816 37016 0 _122_
rlabel metal2 26488 39200 26488 39200 0 _123_
rlabel metal2 23128 26488 23128 26488 0 _124_
rlabel metal3 21784 32872 21784 32872 0 _125_
rlabel metal2 23464 36008 23464 36008 0 _126_
rlabel metal2 21336 36960 21336 36960 0 _127_
rlabel metal2 19544 39648 19544 39648 0 _128_
rlabel metal2 23968 20888 23968 20888 0 _129_
rlabel metal3 22120 34104 22120 34104 0 _130_
rlabel metal2 25200 34216 25200 34216 0 _131_
rlabel metal3 25088 37016 25088 37016 0 _132_
rlabel metal2 24136 39648 24136 39648 0 _133_
rlabel metal2 23912 38080 23912 38080 0 _134_
rlabel metal3 22568 38920 22568 38920 0 _135_
rlabel metal2 14952 39032 14952 39032 0 _136_
rlabel metal2 22456 7840 22456 7840 0 _137_
rlabel metal2 21672 21140 21672 21140 0 _138_
rlabel metal2 25480 20496 25480 20496 0 _139_
rlabel metal2 25368 12432 25368 12432 0 _140_
rlabel metal2 27440 6664 27440 6664 0 _141_
rlabel metal2 28056 5936 28056 5936 0 _142_
rlabel metal2 25928 26992 25928 26992 0 _143_
rlabel metal2 25928 6720 25928 6720 0 _144_
rlabel metal3 27496 6552 27496 6552 0 _145_
rlabel metal3 27384 5656 27384 5656 0 _146_
rlabel metal2 26376 5544 26376 5544 0 _147_
rlabel metal2 25704 5824 25704 5824 0 _148_
rlabel metal2 27832 7560 27832 7560 0 _149_
rlabel metal2 22848 8232 22848 8232 0 _150_
rlabel metal2 23128 6944 23128 6944 0 _151_
rlabel metal2 22792 5040 22792 5040 0 _152_
rlabel metal2 23352 8316 23352 8316 0 _153_
rlabel metal3 24360 26152 24360 26152 0 _154_
rlabel metal3 23408 8232 23408 8232 0 _155_
rlabel metal3 29512 10584 29512 10584 0 _156_
rlabel metal2 29624 10360 29624 10360 0 _157_
rlabel metal2 27496 9520 27496 9520 0 _158_
rlabel metal2 30632 12600 30632 12600 0 _159_
rlabel metal2 32984 11592 32984 11592 0 _160_
rlabel metal3 30072 12936 30072 12936 0 _161_
rlabel metal2 29960 12264 29960 12264 0 _162_
rlabel metal2 29232 15064 29232 15064 0 _163_
rlabel metal2 25816 23912 25816 23912 0 _164_
rlabel metal2 30296 16072 30296 16072 0 _165_
rlabel metal2 24136 17248 24136 17248 0 _166_
rlabel metal2 25592 29456 25592 29456 0 _167_
rlabel metal2 31864 29120 31864 29120 0 _168_
rlabel metal3 34720 30184 34720 30184 0 _169_
rlabel metal2 37352 29288 37352 29288 0 _170_
rlabel metal2 36120 27664 36120 27664 0 _171_
rlabel metal2 26600 16352 26600 16352 0 _172_
rlabel metal2 38920 24584 38920 24584 0 _173_
rlabel metal3 38808 31864 38808 31864 0 _174_
rlabel metal2 37016 28560 37016 28560 0 _175_
rlabel metal2 39032 28392 39032 28392 0 _176_
rlabel metal2 7336 33264 7336 33264 0 _177_
rlabel metal2 39816 27832 39816 27832 0 _178_
rlabel metal2 35392 30744 35392 30744 0 _179_
rlabel metal3 35336 30968 35336 30968 0 _180_
rlabel metal2 39368 31416 39368 31416 0 _181_
rlabel metal2 36120 31248 36120 31248 0 _182_
rlabel metal2 37464 36008 37464 36008 0 _183_
rlabel metal2 37128 35392 37128 35392 0 _184_
rlabel metal3 39032 32760 39032 32760 0 _185_
rlabel metal3 41104 31640 41104 31640 0 _186_
rlabel metal2 41552 37912 41552 37912 0 _187_
rlabel metal3 41160 38808 41160 38808 0 _188_
rlabel metal2 41328 37464 41328 37464 0 _189_
rlabel metal2 40600 38416 40600 38416 0 _190_
rlabel metal2 40040 36008 40040 36008 0 _191_
rlabel metal2 40488 36176 40488 36176 0 _192_
rlabel metal3 39312 34664 39312 34664 0 _193_
rlabel metal2 37464 38192 37464 38192 0 _194_
rlabel metal2 41664 31976 41664 31976 0 _195_
rlabel metal2 41160 32592 41160 32592 0 _196_
rlabel metal2 42392 24360 42392 24360 0 _197_
rlabel metal2 41776 21000 41776 21000 0 _198_
rlabel metal2 40600 26992 40600 26992 0 _199_
rlabel metal2 42504 28784 42504 28784 0 _200_
rlabel metal2 41384 18648 41384 18648 0 _201_
rlabel metal2 42056 19096 42056 19096 0 _202_
rlabel metal2 39928 23688 39928 23688 0 _203_
rlabel metal2 13160 26040 13160 26040 0 _204_
rlabel metal2 35504 18424 35504 18424 0 _205_
rlabel metal2 35560 17920 35560 17920 0 _206_
rlabel metal2 35056 17752 35056 17752 0 _207_
rlabel metal2 41160 17416 41160 17416 0 _208_
rlabel metal2 41608 17920 41608 17920 0 _209_
rlabel metal2 36288 19208 36288 19208 0 _210_
rlabel metal2 37352 17584 37352 17584 0 _211_
rlabel metal2 37464 16128 37464 16128 0 _212_
rlabel metal2 36680 25088 36680 25088 0 _213_
rlabel metal2 36568 24080 36568 24080 0 _214_
rlabel metal2 35448 22120 35448 22120 0 _215_
rlabel metal2 42000 23912 42000 23912 0 _216_
rlabel metal2 41216 24696 41216 24696 0 _217_
rlabel metal3 19208 26376 19208 26376 0 _218_
rlabel metal3 39172 23128 39172 23128 0 _219_
rlabel metal2 39256 23800 39256 23800 0 _220_
rlabel metal2 17920 23128 17920 23128 0 _221_
rlabel metal2 18424 27160 18424 27160 0 _222_
rlabel metal2 12936 27552 12936 27552 0 _223_
rlabel metal2 13720 22792 13720 22792 0 _224_
rlabel metal3 17752 20216 17752 20216 0 _225_
rlabel metal2 12712 10640 12712 10640 0 _226_
rlabel metal2 11144 30632 11144 30632 0 _227_
rlabel metal2 11480 30912 11480 30912 0 _228_
rlabel metal2 17864 16464 17864 16464 0 _229_
rlabel metal2 17976 16744 17976 16744 0 _230_
rlabel metal2 17528 17304 17528 17304 0 _231_
rlabel metal2 18424 22680 18424 22680 0 _232_
rlabel metal2 11368 17136 11368 17136 0 _233_
rlabel metal2 19768 22120 19768 22120 0 _234_
rlabel metal2 10752 28840 10752 28840 0 _235_
rlabel metal3 20160 19880 20160 19880 0 _236_
rlabel metal2 19208 23464 19208 23464 0 _237_
rlabel metal2 18648 22512 18648 22512 0 _238_
rlabel metal2 19320 24584 19320 24584 0 _239_
rlabel metal3 20664 22456 20664 22456 0 _240_
rlabel metal2 3864 23016 3864 23016 0 _241_
rlabel metal2 16072 24024 16072 24024 0 _242_
rlabel metal2 16240 24584 16240 24584 0 _243_
rlabel metal2 14728 21224 14728 21224 0 _244_
rlabel metal2 9016 23912 9016 23912 0 _245_
rlabel metal3 9744 23352 9744 23352 0 _246_
rlabel metal2 11256 23968 11256 23968 0 _247_
rlabel metal2 11424 24024 11424 24024 0 _248_
rlabel metal2 10920 21392 10920 21392 0 _249_
rlabel metal2 6552 18480 6552 18480 0 _250_
rlabel metal2 8512 24920 8512 24920 0 _251_
rlabel metal2 6608 26264 6608 26264 0 _252_
rlabel metal2 4088 24360 4088 24360 0 _253_
rlabel metal2 9912 23072 9912 23072 0 _254_
rlabel metal2 10248 22568 10248 22568 0 _255_
rlabel metal3 4984 22456 4984 22456 0 _256_
rlabel metal2 4368 37240 4368 37240 0 _257_
rlabel metal2 6384 19096 6384 19096 0 _258_
rlabel metal2 6216 22792 6216 22792 0 _259_
rlabel metal2 6440 25368 6440 25368 0 _260_
rlabel metal3 5152 25592 5152 25592 0 _261_
rlabel metal2 6776 18368 6776 18368 0 _262_
rlabel metal2 5656 18704 5656 18704 0 _263_
rlabel metal3 7112 17416 7112 17416 0 _264_
rlabel metal3 5936 18424 5936 18424 0 _265_
rlabel metal2 5544 18200 5544 18200 0 _266_
rlabel metal2 7784 16016 7784 16016 0 _267_
rlabel metal3 9912 15288 9912 15288 0 _268_
rlabel metal2 7336 18032 7336 18032 0 _269_
rlabel metal2 8120 13440 8120 13440 0 _270_
rlabel metal2 7784 14168 7784 14168 0 _271_
rlabel metal2 10024 15008 10024 15008 0 _272_
rlabel metal2 9688 15792 9688 15792 0 _273_
rlabel metal2 24472 20720 24472 20720 0 _274_
rlabel metal2 7448 10304 7448 10304 0 _275_
rlabel metal2 7504 11368 7504 11368 0 _276_
rlabel metal3 29624 30688 29624 30688 0 _277_
rlabel metal2 19768 16240 19768 16240 0 _278_
rlabel metal3 11760 15176 11760 15176 0 _279_
rlabel metal2 6552 10416 6552 10416 0 _280_
rlabel metal2 6776 10080 6776 10080 0 _281_
rlabel metal2 7784 12880 7784 12880 0 _282_
rlabel metal3 8288 12152 8288 12152 0 _283_
rlabel metal2 8680 11088 8680 11088 0 _284_
rlabel metal2 8400 11480 8400 11480 0 _285_
rlabel metal2 11592 12432 11592 12432 0 _286_
rlabel metal3 13608 11256 13608 11256 0 _287_
rlabel metal3 11480 10584 11480 10584 0 _288_
rlabel metal2 11592 10304 11592 10304 0 _289_
rlabel metal2 11144 8792 11144 8792 0 _290_
rlabel metal2 14392 9912 14392 9912 0 _291_
rlabel metal2 12600 10864 12600 10864 0 _292_
rlabel metal2 12936 9800 12936 9800 0 _293_
rlabel metal2 12376 9016 12376 9016 0 _294_
rlabel metal2 15736 10472 15736 10472 0 _295_
rlabel metal2 16072 11816 16072 11816 0 _296_
rlabel metal2 13832 11760 13832 11760 0 _297_
rlabel metal3 16576 11368 16576 11368 0 _298_
rlabel metal2 16968 11368 16968 11368 0 _299_
rlabel metal2 19208 10472 19208 10472 0 _300_
rlabel metal2 16408 9912 16408 9912 0 _301_
rlabel metal2 19096 9912 19096 9912 0 _302_
rlabel metal2 18312 8316 18312 8316 0 _303_
rlabel metal2 11144 27048 11144 27048 0 _304_
rlabel metal2 11088 29176 11088 29176 0 _305_
rlabel metal2 7784 35672 7784 35672 0 _306_
rlabel metal3 6160 36680 6160 36680 0 _307_
rlabel metal3 7224 33096 7224 33096 0 _308_
rlabel metal2 5208 36232 5208 36232 0 _309_
rlabel metal3 17808 26264 17808 26264 0 _310_
rlabel metal2 19096 26992 19096 26992 0 _311_
rlabel metal2 30184 33544 30184 33544 0 _312_
rlabel metal3 16184 33208 16184 33208 0 _313_
rlabel metal2 18704 27832 18704 27832 0 _314_
rlabel metal2 25256 27552 25256 27552 0 _315_
rlabel metal2 16296 29960 16296 29960 0 _316_
rlabel metal2 15400 33768 15400 33768 0 _317_
rlabel metal2 12208 33208 12208 33208 0 _318_
rlabel metal2 11816 32984 11816 32984 0 _319_
rlabel metal3 7168 30632 7168 30632 0 _320_
rlabel metal2 10976 32984 10976 32984 0 _321_
rlabel metal2 10696 33992 10696 33992 0 _322_
rlabel metal2 7392 30408 7392 30408 0 _323_
rlabel metal2 30520 22008 30520 22008 0 _324_
rlabel metal2 29512 25424 29512 25424 0 _325_
rlabel metal2 28560 24696 28560 24696 0 _326_
rlabel metal2 29064 24696 29064 24696 0 _327_
rlabel metal2 27384 22008 27384 22008 0 _328_
rlabel metal2 31752 33992 31752 33992 0 _329_
rlabel metal2 27608 35168 27608 35168 0 bcd\[0\]
rlabel metal2 20608 31864 20608 31864 0 bcd\[1\]
rlabel metal2 7784 39984 7784 39984 0 bcd\[2\]
rlabel metal2 7000 38136 7000 38136 0 clkdiv\[0\]
rlabel metal2 7000 30688 7000 30688 0 clkdiv\[1\]
rlabel metal2 22680 27384 22680 27384 0 clkdiv\[2\]
rlabel metal2 16296 28560 16296 28560 0 clkdiv\[3\]
rlabel metal2 13832 31052 13832 31052 0 clkdiv\[4\]
rlabel metal3 6440 32648 6440 32648 0 clkdiv\[5\]
rlabel metal2 7784 37408 7784 37408 0 clkdiv\[6\]
rlabel metal2 6104 30912 6104 30912 0 clkdiv\[7\]
rlabel metal3 25592 30856 25592 30856 0 clknet_0_wb_clk_i
rlabel metal2 1960 18816 1960 18816 0 clknet_3_0__leaf_wb_clk_i
rlabel metal2 21280 5096 21280 5096 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 1848 27832 1848 27832 0 clknet_3_2__leaf_wb_clk_i
rlabel metal3 18872 28728 18872 28728 0 clknet_3_3__leaf_wb_clk_i
rlabel metal2 27048 5488 27048 5488 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 32704 8232 32704 8232 0 clknet_3_5__leaf_wb_clk_i
rlabel metal3 28560 26936 28560 26936 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 40656 29400 40656 29400 0 clknet_3_7__leaf_wb_clk_i
rlabel metal2 17640 24136 17640 24136 0 counter\[0\]
rlabel metal3 7672 15288 7672 15288 0 counter\[10\]
rlabel metal2 7784 15260 7784 15260 0 counter\[11\]
rlabel metal2 15176 10528 15176 10528 0 counter\[12\]
rlabel metal2 14616 7392 14616 7392 0 counter\[13\]
rlabel metal2 16688 11256 16688 11256 0 counter\[14\]
rlabel metal3 18536 9688 18536 9688 0 counter\[15\]
rlabel metal2 20216 19600 20216 19600 0 counter\[1\]
rlabel metal2 21448 25536 21448 25536 0 counter\[2\]
rlabel metal2 15624 26264 15624 26264 0 counter\[3\]
rlabel metal2 13664 26936 13664 26936 0 counter\[4\]
rlabel metal3 6328 29400 6328 29400 0 counter\[5\]
rlabel metal2 10304 23128 10304 23128 0 counter\[6\]
rlabel metal2 5880 28588 5880 28588 0 counter\[7\]
rlabel metal2 5768 16520 5768 16520 0 counter\[8\]
rlabel metal2 8680 15680 8680 15680 0 counter\[9\]
rlabel metal2 9464 44478 9464 44478 0 io_in
rlabel metal3 13888 41832 13888 41832 0 io_out[0]
rlabel metal2 17640 45304 17640 45304 0 io_out[1]
rlabel metal2 21448 45304 21448 45304 0 io_out[2]
rlabel metal3 25312 41832 25312 41832 0 io_out[3]
rlabel metal2 28728 41832 28728 41832 0 io_out[4]
rlabel metal2 32872 45304 32872 45304 0 io_out[5]
rlabel metal2 36680 45304 36680 45304 0 io_out[6]
rlabel metal3 40544 41832 40544 41832 0 io_out[7]
rlabel metal2 43736 43274 43736 43274 0 io_out[8]
rlabel metal2 31864 27384 31864 27384 0 lfsr\[0\]
rlabel metal2 35784 18032 35784 18032 0 lfsr\[10\]
rlabel metal2 41608 18480 41608 18480 0 lfsr\[11\]
rlabel metal2 40264 15736 40264 15736 0 lfsr\[12\]
rlabel metal2 36344 22456 36344 22456 0 lfsr\[13\]
rlabel metal3 43876 25592 43876 25592 0 lfsr\[14\]
rlabel metal2 41832 24360 41832 24360 0 lfsr\[15\]
rlabel metal3 30632 30128 30632 30128 0 lfsr\[1\]
rlabel metal2 35112 30968 35112 30968 0 lfsr\[2\]
rlabel metal3 39816 37912 39816 37912 0 lfsr\[4\]
rlabel metal2 43848 35896 43848 35896 0 lfsr\[5\]
rlabel metal3 35952 37912 35952 37912 0 lfsr\[6\]
rlabel metal2 40488 33320 40488 33320 0 lfsr\[7\]
rlabel metal2 42560 28504 42560 28504 0 lfsr\[8\]
rlabel metal2 42392 19488 42392 19488 0 lfsr\[9\]
rlabel metal3 22456 13608 22456 13608 0 m_clkdiv\[0\]
rlabel metal2 24752 13720 24752 13720 0 m_clkdiv\[1\]
rlabel metal2 27384 5096 27384 5096 0 m_clkdiv\[2\]
rlabel metal2 26488 6776 26488 6776 0 m_clkdiv\[3\]
rlabel metal3 27216 9016 27216 9016 0 m_clkdiv\[4\]
rlabel metal3 28896 8344 28896 8344 0 m_clkdiv\[5\]
rlabel metal2 33040 12040 33040 12040 0 m_clkdiv\[6\]
rlabel metal2 30856 13216 30856 13216 0 m_clkdiv\[7\]
rlabel metal2 29288 16352 29288 16352 0 m_clkdiv\[8\]
rlabel metal2 28392 16464 28392 16464 0 m_clkdiv\[9\]
rlabel metal2 10248 31556 10248 31556 0 net1
rlabel metal2 30856 34160 30856 34160 0 net10
rlabel metal3 38640 38920 38640 38920 0 net11
rlabel metal2 6216 39256 6216 39256 0 net2
rlabel metal2 12712 41104 12712 41104 0 net3
rlabel metal2 16184 41104 16184 41104 0 net4
rlabel metal2 20552 41104 20552 41104 0 net5
rlabel metal2 23576 40264 23576 40264 0 net6
rlabel metal2 30632 41104 30632 41104 0 net7
rlabel metal2 32648 40824 32648 40824 0 net8
rlabel metal2 36008 41104 36008 41104 0 net9
rlabel metal2 31640 24024 31640 24024 0 r_counter\[0\]
rlabel metal2 31248 30184 31248 30184 0 r_counter\[1\]
rlabel metal2 30856 28924 30856 28924 0 r_counter\[2\]
rlabel metal2 5656 44478 5656 44478 0 rst_n
rlabel metal2 22008 22064 22008 22064 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 46000 46000
<< end >>
