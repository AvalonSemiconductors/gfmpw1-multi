* NGSPICE file created from wrapped_ay8913.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

.subckt wrapped_ay8913 custom_settings[0] custom_settings[1] custom_settings[2] custom_settings[3]
+ io_in_1[0] io_in_1[1] io_in_1[2] io_in_1[3] io_in_1[4] io_in_1[5] io_in_1[6] io_in_1[7]
+ io_in_2[0] io_in_2[1] io_out[10] io_out[11] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[2]
+ io_out[3] io_out[4] io_out[5] io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i
+ io_out[16] io_out[15] io_out[0] io_out[14] io_out[13] io_out[12] io_out[22] io_out[6]
X_2106_ tt_um_rejunity_ay8913.tone_B_generator.counter\[3\] _0626_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2037_ _0529_ _0569_ _0526_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1445__A1 _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1693__A1 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1270_ blink.counter\[7\] _0897_ _0904_ _0911_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1389__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1606_ tt_um_rejunity_ay8913.pwm_A.accumulator\[2\] _0868_ _1156_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2586_ _0200_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1537_ _1003_ tt_um_rejunity_ay8913.tone_B_generator.period\[8\] _1111_ _1112_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1468_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\] _1062_ _1063_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\]
+ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1399_ tt_um_rejunity_ay8913.pwm_master.accumulator\[2\] net20 _1008_ _1009_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1675__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1969__A2 _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ _0054_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_11_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1253_ _0890_ _0899_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1322_ _0946_ _0945_ _0947_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2371_ _0991_ _1173_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1657__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1409__A1 _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2569_ _0183_ clknet_leaf_21_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2638_ _0252_ clknet_leaf_32_wb_clk_i tt_um_rejunity_ay8913.envelope_B vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1351__A3 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1871_ _0347_ _0429_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1940_ _0482_ _0483_ _0478_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2423_ _0037_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1236_ _0875_ _0886_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1305_ blink.counter\[20\] _0932_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2354_ _0828_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2285_ _0782_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1869__A1 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2070_ _0594_ _0595_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1785_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\] _0357_ _0360_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1854_ _0409_ _0418_ _0419_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_44_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_12_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1923_ tt_um_rejunity_ay8913.noise_generator.lfsr\[10\] _0464_ _0471_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2406_ _0020_ clknet_leaf_42_wb_clk_i blink.counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2268_ _0766_ _0769_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1219_ _0870_ _0868_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2337_ _0816_ tt_um_rejunity_ay8913.tone_A_generator.period\[8\] _0817_ _0818_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2199_ _0701_ tt_um_rejunity_ay8913.tone_A_generator.period\[8\] _0703_ _0705_ _0706_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_14_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1570_ _1132_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2122_ tt_um_rejunity_ay8913.tone_B_generator.period\[6\] _0642_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2053_ _0574_ _0582_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1768_ tt_um_rejunity_ay8913.envelope_generator.period\[10\] _0343_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1837_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\] _0401_ _0402_ _0407_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1906_ tt_um_rejunity_ay8913.noise_generator.lfsr\[4\] _0458_ _0459_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1699_ _0260_ _0283_ _0285_ tt_um_rejunity_ay8913.tone_disable_A _0286_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput20 net20 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1622_ _1166_ _1167_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1553_ _1122_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1484_ _1072_ _1073_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2105_ _0617_ _0624_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2036_ _0533_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1206__A2 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1693__A2 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2585_ _0199_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1605_ _1155_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1536_ _1109_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1372__A1 _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1398_ _1007_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1467_ _1057_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2019_ tt_um_rejunity_ay8913.tone_C_generator.period\[6\] _0552_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1363__A1 _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2091__A2 _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1252_ blink.counter\[4\] _0898_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1321_ _0946_ _0945_ _0892_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2370_ _1177_ _0836_ _0837_ _0854_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_46_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2499_ _0113_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1519_ _1091_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2568_ _0182_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2637_ _0251_ clknet_leaf_32_wb_clk_i tt_um_rejunity_ay8913.amplitude_B\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_39_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_39_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1351__A4 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1870_ _0347_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_54_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2422_ _0036_ clknet_leaf_21_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2353_ _0268_ _0823_ _0825_ tt_um_rejunity_ay8913.envelope_generator.period\[2\]
+ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1235_ _0881_ _0883_ _0884_ _0885_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1304_ blink.counter\[20\] _0932_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2284_ _0754_ _0780_ _0781_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1566__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1999_ tt_um_rejunity_ay8913.tone_C_generator.counter\[9\] _0532_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_3_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1922_ _0468_ _0470_ _0467_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1784_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\] _0343_ _0359_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1548__A1 _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1853_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\] _0332_ _0413_ _0411_
+ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2405_ _0019_ clknet_leaf_3_wb_clk_i blink.counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2336_ _0814_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2267_ _0767_ _0768_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1218_ _0863_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2198_ _0702_ tt_um_rejunity_ay8913.tone_A_generator.period\[11\] tt_um_rejunity_ay8913.tone_A_generator.period\[10\]
+ _0704_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2121_ tt_um_rejunity_ay8913.tone_B_generator.period\[7\] _0641_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2052_ tt_um_rejunity_ay8913.tone_C_generator.counter\[3\] _0581_ _0582_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1905_ _0443_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1767_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\] _0342_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1836_ _0315_ _0405_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1698_ _0284_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2319_ net13 net12 _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input11_I io_in_1[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput21 net21 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1552_ _0980_ _1118_ _1120_ tt_um_rejunity_ay8913.tone_B_generator.period\[1\] _1122_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1621_ tt_um_rejunity_ay8913.pwm_A.accumulator\[6\] _1163_ _1161_ _1167_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input3_I custom_settings[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2104_ _0619_ _0623_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1483_ tt_um_rejunity_ay8913.pwm_C.accumulator\[3\] _1070_ _1034_ _1073_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2035_ _0567_ _0556_ _0535_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_17_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1819_ _0386_ _0392_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2584_ _0198_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1535_ _1109_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1604_ _1021_ tt_um_rejunity_ay8913.pwm_B.accumulator\[7\] tt_um_rejunity_ay8913.pwm_B.accumulator\[8\]
+ _1150_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_1_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1466_ _1044_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1397_ _0994_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2018_ tt_um_rejunity_ay8913.tone_C_generator.period\[7\] _0551_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1320_ blink.counter\[25\] _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1251_ _0893_ _0896_ _0898_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_54_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_9_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2636_ _0250_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.envelope_C vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1518_ _1089_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2498_ _0112_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2567_ _0181_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1449_ net21 _1048_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2421_ _0035_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2352_ _0827_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1303_ _0888_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2283_ _0711_ _0779_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1234_ blink.counter\[30\] blink.counter\[29\] blink.counter\[28\] blink.counter\[27\]
+ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1998_ tt_um_rejunity_ay8913.tone_C_generator.period\[9\] _0531_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2619_ _0233_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.latched_register\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1852_ _0340_ _0417_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_44_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1921_ tt_um_rejunity_ay8913.noise_generator.lfsr\[8\] _0469_ _0470_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1783_ _0356_ _0357_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1548__A2 _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2404_ _0018_ clknet_leaf_2_wb_clk_i blink.counter\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2266_ tt_um_rejunity_ay8913.tone_A_generator.counter\[5\] _0722_ tt_um_rejunity_ay8913.tone_A_generator.counter\[3\]
+ _0760_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2335_ _0995_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1217_ _0869_ net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2197_ tt_um_rejunity_ay8913.tone_A_generator.counter\[10\] _0704_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2120_ _0629_ _0631_ _0639_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
Xclkbuf_leaf_23_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_23_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2051_ _0537_ _0576_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1835_ _0401_ _0402_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1904_ tt_um_rejunity_ay8913.noise_generator.lfsr\[5\] _0453_ _0457_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1766_ _0339_ tt_um_rejunity_ay8913.envelope_generator.period\[9\] tt_um_rejunity_ay8913.envelope_generator.period\[8\]
+ _0340_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1697_ _1010_ _0282_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2188__C _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2249__A3 _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2249_ tt_um_rejunity_ay8913.tone_A_generator.counter\[1\] tt_um_rejunity_ay8913.tone_A_generator.counter\[0\]
+ _0387_ _0388_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2318_ _0804_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput22 net22 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1551_ _1121_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _1165_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1482_ tt_um_rejunity_ay8913.pwm_C.accumulator\[3\] _1070_ _1072_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2103_ tt_um_rejunity_ay8913.tone_B_generator.counter\[10\] _0620_ _0621_ _0622_
+ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2034_ _0565_ _0566_ _0554_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1818_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\] _0391_ _0392_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1749_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\] _0324_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_7_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1669__A1 _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1534_ _1107_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1603_ _1012_ _1154_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1465_ _1056_ _1061_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2583_ _0197_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_C vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2017_ _0539_ _0541_ _0549_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1396_ _1005_ _0993_ _1006_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1250_ _0897_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_19_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2635_ _0249_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.amplitude_C\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1517_ _1096_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2497_ _0111_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2566_ _0180_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1448_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\] tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
+ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1379_ _0992_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2420_ _0034_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1302_ _0923_ _0932_ _0933_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1233_ blink.counter\[26\] blink.counter\[25\] blink.counter\[24\] blink.counter\[23\]
+ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_2351_ _0266_ _0823_ _0825_ tt_um_rejunity_ay8913.envelope_generator.period\[1\]
+ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2282_ _0711_ _0779_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1997_ tt_um_rejunity_ay8913.tone_C_generator.period\[10\] _0530_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2549_ _0163_ clknet_leaf_40_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2618_ _0232_ clknet_leaf_32_wb_clk_i tt_um_rejunity_ay8913.latched_register\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1851_ _0332_ _0413_ _0412_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1975__I _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1920_ _0443_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1782_ tt_um_rejunity_ay8913.envelope_generator.period\[11\] _0357_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2403_ _0017_ clknet_leaf_4_wb_clk_i blink.counter\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2265_ _0722_ _0763_ tt_um_rejunity_ay8913.tone_A_generator.counter\[5\] _0767_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1216_ _0860_ _0863_ _0868_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2196_ _0702_ tt_um_rejunity_ay8913.tone_A_generator.period\[11\] _0703_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2334_ _0814_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2050_ _0580_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_32_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1765_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\] _0340_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1834_ _0385_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1903_ _0454_ _0455_ _0456_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1696_ _0282_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2179_ tt_um_rejunity_ay8913.tone_B_generator.counter\[8\] _0684_ _0690_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2249__A4 _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2248_ _0752_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2317_ net13 net12 _0803_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_31_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput23 net23 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1550_ _0964_ _1118_ _1120_ tt_um_rejunity_ay8913.tone_B_generator.period\[0\] _1121_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1481_ _1070_ _1071_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1384__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2033_ _0555_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2102_ tt_um_rejunity_ay8913.tone_B_generator.counter\[9\] _0622_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1817_ _0390_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1748_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\] _0323_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_7_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1679_ _1176_ _0272_ _0273_ tt_um_rejunity_ay8913.tone_A_generator.period\[4\] _0274_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_51_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1366__A1 _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1294__B _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2582_ _0196_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1602_ tt_um_rejunity_ay8913.pwm_B.accumulator\[8\] _1153_ _1154_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1464_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\] _1047_ _1058_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\]
+ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1533_ _0968_ _0990_ _0970_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1395_ _1003_ tt_um_rejunity_ay8913.tone_C_generator.period\[11\] _0997_ _1006_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_22_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2016_ _0545_ _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_19_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1520__A1 _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1823__A2 _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1516_ _0984_ _1090_ _1092_ tt_um_rejunity_ay8913.tone_C_generator.period\[3\] _1096_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2565_ _0179_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2634_ _0248_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1447_ _1044_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2496_ _0110_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.envelope_A vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1378_ _0967_ _0991_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1569__A1 _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_17_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_17_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1301_ blink.counter\[19\] _0931_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2350_ _0826_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1232_ blink.counter\[19\] _0882_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2281_ tt_um_rejunity_ay8913.tone_A_generator.counter\[8\] _0773_ _0779_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1996_ _0528_ tt_um_rejunity_ay8913.tone_C_generator.period\[9\] tt_um_rejunity_ay8913.tone_C_generator.period\[8\]
+ _0522_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2617_ _0231_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.active vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2548_ _0162_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2479_ _0093_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1781_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\] _0356_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1850_ _0404_ _0416_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_44_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2402_ _0016_ clknet_leaf_5_wb_clk_i blink.counter\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1705__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2333_ _0991_ _1107_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1215_ _0867_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2264_ _0754_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2195_ tt_um_rejunity_ay8913.tone_A_generator.counter\[11\] _0702_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_35_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\] _0512_ _0516_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2188__A1 _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_32_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_32_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1902_ _0446_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1764_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\] _0339_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1833_ _0394_ _0403_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2316_ net8 net11 net10 net9 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__2351__A1 _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1695_ _0967_ _1108_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2178_ _0689_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2247_ _0700_ _0753_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1480_ tt_um_rejunity_ay8913.pwm_C.accumulator\[2\] _0860_ _1034_ _1071_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2032_ tt_um_rejunity_ay8913.tone_C_generator.counter\[5\] _0561_ _0545_ _0564_ _0565_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2101_ tt_um_rejunity_ay8913.tone_B_generator.period\[9\] _0621_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1747_ _0320_ tt_um_rejunity_ay8913.envelope_generator.period\[0\] _0321_ _0322_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1816_ _0389_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1678_ _0263_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_51_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2315__A1 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2581_ _0195_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1601_ tt_um_rejunity_ay8913.pwm_B.accumulator\[7\] _1149_ _1153_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1532_ _0965_ _1106_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input1_I custom_settings[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1394_ net7 _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1463_ _1056_ _1060_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2015_ tt_um_rejunity_ay8913.tone_C_generator.counter\[3\] _0546_ _0547_ tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
+ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_36_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1515_ _1095_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2633_ _0247_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2564_ _0178_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.noise_generator.signal_edge.signal
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2495_ _0109_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.amplitude_A\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1446_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\] _1046_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1377_ tt_um_rejunity_ay8913.latched_register\[1\] _0990_ _0970_ _0991_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_16_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1300_ blink.counter\[19\] _0931_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1231_ blink.counter\[22\] blink.counter\[21\] blink.counter\[20\] _0882_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_19_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2280_ _0778_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1995_ tt_um_rejunity_ay8913.tone_C_generator.counter\[9\] _0528_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2616_ _0230_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2478_ _0092_ clknet_leaf_30_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1429_ _0995_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2547_ _0161_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1780_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\] _0348_ _0354_
+ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1953__A2 _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2401_ _0015_ clknet_leaf_5_wb_clk_i blink.counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2332_ _0813_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2263_ _0765_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1469__A1 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1214_ _0864_ _0865_ _0857_ tt_um_rejunity_ay8913.envelope_A _0866_ _0867_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_2194_ tt_um_rejunity_ay8913.tone_A_generator.counter\[8\] _0701_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1641__A1 _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\] _0512_ _0515_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_2_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_11_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2188__A2 _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1699__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1832_ _0401_ _0402_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_32_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1901_ tt_um_rejunity_ay8913.noise_generator.lfsr\[3\] _0444_ _0455_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1763_ _0336_ tt_um_rejunity_ay8913.envelope_generator.period\[13\] tt_um_rejunity_ay8913.envelope_generator.period\[12\]
+ _0337_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1694_ _0281_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1507__I _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2246_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2315_ _1082_ _0801_ _0802_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2177_ _0677_ _0688_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_35_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2100_ tt_um_rejunity_ay8913.tone_B_generator.period\[10\] _0620_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2031_ _0539_ _0563_ _0548_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1997__I tt_um_rejunity_ay8913.tone_C_generator.period\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1815_ _0387_ _0388_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1946__B _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1746_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\] tt_um_rejunity_ay8913.envelope_generator.period\[1\]
+ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1677_ _0261_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2229_ _0733_ _0734_ _0735_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2580_ _0194_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1600_ tt_um_rejunity_ay8913.pwm_B.accumulator\[7\] _1150_ _1152_ _0098_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1462_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\] _1047_ _1058_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\]
+ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1531_ tt_um_rejunity_ay8913.latched_register\[2\] _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1393_ _1001_ _0993_ _1004_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2014_ tt_um_rejunity_ay8913.tone_C_generator.period\[4\] _0547_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1729_ _0294_ _0306_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_19_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _0246_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1514_ _0982_ _1090_ _1092_ tt_um_rejunity_ay8913.tone_C_generator.period\[2\] _1095_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2494_ _0108_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1445_ _1037_ _1045_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_10_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2563_ _0177_ clknet_leaf_40_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1376_ tt_um_rejunity_ay8913.latched_register\[0\] _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_2_2__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1230_ _0876_ _0880_ blink.counter\[18\] _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_26_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_26_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ _0522_ tt_um_rejunity_ay8913.tone_C_generator.period\[8\] _0524_ _0526_ _0527_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ _0229_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2477_ _0091_ clknet_leaf_30_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1428_ _1032_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2546_ _0160_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.invert_output
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1359_ _0977_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0014_ clknet_leaf_8_wb_clk_i blink.counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2262_ _0753_ _0764_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2331_ blink.LED _0889_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1213_ tt_um_rejunity_ay8913.amplitude_A\[0\] tt_um_rejunity_ay8913.envelope_A tt_um_rejunity_ay8913.tone_disable_A
+ tt_um_rejunity_ay8913.tone_A _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_47_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2193_ _0699_ _0391_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1641__A2 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ _0511_ _0512_ _0514_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_7_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2529_ _0143_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1396__A1 _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ _0324_ _0323_ _0320_ _0382_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_32_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1900_ tt_um_rejunity_ay8913.noise_generator.lfsr\[4\] _0453_ _0454_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1762_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\] _0337_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1387__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1693_ tt_um_rejunity_ay8913.noise_generator.signal_edge.signal _1086_ _0281_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_41_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_41_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2176_ tt_um_rejunity_ay8913.tone_B_generator.counter\[8\] _0684_ _0688_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2245_ _0390_ _0751_ _0975_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2314_ _0799_ tt_um_rejunity_ay8913.clk_counter\[6\] _0796_ _0802_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_7_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1550__A1 _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput15 net15 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1369__A1 _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ tt_um_rejunity_ay8913.tone_C_generator.counter\[2\] _0558_ _0562_ _0541_ _0563_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1518__I _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1745_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\] _0320_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1814_ _0381_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_40_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1676_ _0271_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2159_ _0633_ _0674_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2228_ tt_um_rejunity_ay8913.tone_A_generator.counter\[7\] _0730_ _0735_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1523__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ _1105_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1461_ _1056_ _1059_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1392_ _1003_ tt_um_rejunity_ay8913.tone_C_generator.period\[10\] _0997_ _1004_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2013_ tt_um_rejunity_ay8913.tone_C_generator.period\[3\] _0546_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1514__A1 _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1728_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\] _0305_ _0306_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_13_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1659_ _1104_ _1187_ _1188_ tt_um_rejunity_ay8913.envelope_generator.period\[15\]
+ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_36_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2631_ _0245_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2562_ _0176_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1513_ _1094_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1444_ net20 _1042_ _1044_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\] _1045_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2493_ _0107_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1375_ _0988_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_16_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1993_ _0523_ tt_um_rejunity_ay8913.tone_C_generator.period\[11\] tt_um_rejunity_ay8913.tone_C_generator.period\[10\]
+ _0525_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2545_ _0159_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2614_ _0228_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1358_ _0976_ _0972_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1427_ _1027_ _1031_ _1025_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2476_ _0090_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1289_ blink.counter\[15\] blink.counter\[14\] blink.counter\[13\] _0919_ _0925_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_18_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2192_ tt_um_rejunity_ay8913.tone_A_generator.counter\[0\] _0699_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2261_ _0722_ _0763_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1212_ tt_um_rejunity_ay8913.noise_disable_A _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2330_ _1172_ _0808_ _0812_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1976_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\] _0513_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
+ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2528_ _0142_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.stop
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2459_ _0073_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1761_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\] _0336_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\] _0401_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1692_ _1043_ _1133_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2313_ _0799_ _0797_ tt_um_rejunity_ay8913.clk_counter\[6\] _0801_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2175_ _0687_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_10_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_10_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2244_ _0714_ _0729_ _0739_ _0747_ _0750_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_43_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1959_ _0498_ tt_um_rejunity_ay8913.noise_generator.period\[1\] tt_um_rejunity_ay8913.noise_generator.period\[0\]
+ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput16 net16 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2327__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1744_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\] _0317_ _0318_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\]
+ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1813_ _0379_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_25_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1675_ _0270_ _0262_ _0264_ tt_um_rejunity_ay8913.tone_A_generator.period\[3\] _0271_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2158_ _0626_ _0627_ _0666_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2227_ tt_um_rejunity_ay8913.tone_A_generator.counter\[6\] _0731_ _0734_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2088__A3 _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2089_ _0608_ _0609_ _0278_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_48_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1460_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\] _1047_ _1058_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\]
+ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1391_ _1002_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2012_ _0542_ tt_um_rejunity_ay8913.tone_C_generator.period\[5\] tt_um_rejunity_ay8913.tone_C_generator.period\[4\]
+ _0544_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1658_ _0258_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1727_ _0302_ _0304_ _0305_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_13_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1589_ tt_um_rejunity_ay8913.pwm_B.accumulator\[4\] _1142_ _1078_ _1145_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1512_ _0980_ _1090_ _1092_ tt_um_rejunity_ay8913.tone_C_generator.period\[1\] _1094_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2630_ _0244_ clknet_leaf_21_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2492_ _0106_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2561_ _0175_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1443_ _1043_ _1041_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_4_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1374_ net4 _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1499__A1 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1653__A1 _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1992_ tt_um_rejunity_ay8913.tone_C_generator.counter\[10\] _0525_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_35_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_35_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2544_ _0158_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2475_ _0089_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2613_ _0227_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1288_ blink.counter\[14\] _0921_ blink.counter\[15\] _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1357_ _0975_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1426_ tt_um_rejunity_ay8913.pwm_master.accumulator\[7\] _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1362__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2260_ _0715_ _0716_ _0755_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1211_ tt_um_rejunity_ay8913.noise_generator.lfsr\[0\] _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2191_ _0697_ _0698_ _0278_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1975_ _0391_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2458_ _0072_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1409_ _1012_ _1016_ _1017_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2527_ _0141_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2389_ _0003_ clknet_leaf_6_wb_clk_i blink.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2290__A1 _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1891__B _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1760_ _0314_ _0331_ _0334_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1357__I _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1691_ _0279_ _1058_ _0280_ _1012_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_27_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2312_ _0799_ _0797_ _0800_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2174_ _0677_ _0686_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_11_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2243_ _0703_ _0749_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1958_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\] _0498_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput17 net17 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1889_ _1054_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1640__I _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1812_ _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1743_ tt_um_rejunity_ay8913.envelope_generator.period\[2\] _0318_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1674_ net7 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2226_ tt_um_rejunity_ay8913.tone_A_generator.counter\[7\] _0730_ _0731_ _0732_ _0733_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2157_ _0673_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2088_ tt_um_rejunity_ay8913.tone_C _0513_ _0572_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_16_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1390_ _0994_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ _0543_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1657_ _1102_ _1187_ _1188_ tt_um_rejunity_ay8913.envelope_generator.period\[14\]
+ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1588_ tt_um_rejunity_ay8913.pwm_B.accumulator\[4\] _1142_ _1144_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1726_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\] _0295_ _0303_
+ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2209_ tt_um_rejunity_ay8913.tone_A_generator.counter\[2\] _0716_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_14_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1455__I _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1511_ _1093_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1365__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1442_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\] _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2491_ _0105_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2560_ _0174_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1373_ _0987_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1709_ net9 _0282_ _0284_ tt_um_rejunity_ay8913.noise_disable_C _0291_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_5_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_5_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_1_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1894__B _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1991_ _0523_ tt_um_rejunity_ay8913.tone_C_generator.period\[11\] _0524_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2612_ _0226_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2543_ _0157_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2474_ _0088_ clknet_leaf_30_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1425_ _1028_ _1030_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1287_ _0888_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1356_ _0974_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_41_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_21_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1210_ tt_um_rejunity_ay8913.noise_generator.lfsr\[0\] _0861_ _0857_ tt_um_rejunity_ay8913.envelope_B
+ _0862_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2190_ tt_um_rejunity_ay8913.tone_B _0520_ _0662_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_47_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1974_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\] tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\]
+ _0390_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_11_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2388_ _0002_ clknet_leaf_6_wb_clk_i blink.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2457_ _0071_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1562__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1408_ tt_um_rejunity_ay8913.pwm_master.accumulator\[2\] _0869_ _1014_ _1015_ _1017_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2526_ _0140_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1339_ _0949_ _0959_ _0960_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2290__A2 _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1690_ net17 _1057_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2311_ _0799_ _0797_ _0790_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2242_ _0708_ _0748_ _0705_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2173_ _0684_ _0685_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1957_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\] _0497_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2509_ _0123_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput18 net18 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1888_ _0864_ _0444_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1526__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1811_ _0293_ _0383_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1368__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1673_ _0269_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1742_ tt_um_rejunity_ay8913.envelope_generator.period\[3\] _0317_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1214__B1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2225_ tt_um_rejunity_ay8913.tone_A_generator.counter\[6\] _0732_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2156_ _0664_ _0672_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2245__A2 _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2087_ _0607_ _0572_ tt_um_rejunity_ay8913.tone_C _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1508__A1 _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1897__B _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1651__I _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2010_ tt_um_rejunity_ay8913.tone_C_generator.counter\[4\] _0543_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_29_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1725_ _0295_ _0303_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\]
+ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1656_ _0257_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1587_ _1142_ _1143_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2139_ _0623_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2208_ tt_um_rejunity_ay8913.tone_A_generator.counter\[3\] _0715_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1510_ _0964_ _1090_ _1092_ tt_um_rejunity_ay8913.tone_C_generator.period\[0\] _1093_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1441_ _1041_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2490_ _0104_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1372_ _0986_ _0972_ _0977_ tt_um_rejunity_ay8913.noise_generator.period\[4\] _0987_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2384__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1708_ _0290_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1639_ _0965_ _1106_ _1088_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_1_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1990_ tt_um_rejunity_ay8913.tone_C_generator.counter\[11\] _0523_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_15_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2542_ _0156_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2611_ _0225_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2473_ _0087_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1355_ net14 _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1424_ _0996_ _1029_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1286_ _0906_ _0922_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_21_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1973_ _1052_ _0508_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2525_ _0139_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ _0001_ clknet_leaf_7_wb_clk_i blink.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2456_ _0070_ clknet_leaf_14_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1338_ _0958_ blink.counter\[28\] _0953_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1407_ tt_um_rejunity_ay8913.pwm_master.accumulator\[2\] _0869_ _1014_ _1015_ _1016_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1269_ blink.counter\[9\] blink.counter\[8\] _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2172_ _0643_ _0679_ tt_um_rejunity_ay8913.tone_B_generator.counter\[7\] _0685_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2310_ tt_um_rejunity_ay8913.clk_counter\[5\] _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2241_ _0712_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1956_ _0495_ _0496_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1887_ _0443_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2508_ _0122_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput19 net19 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2439_ _0053_ clknet_leaf_28_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1741_ _0315_ tt_um_rejunity_ay8913.envelope_generator.period\[4\] _0316_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1214__A1 _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1810_ _0311_ _0383_ _0384_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1672_ _0268_ _0262_ _0264_ tt_um_rejunity_ay8913.tone_A_generator.period\[2\] _0269_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2190__A2 _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2155_ tt_um_rejunity_ay8913.tone_B_generator.counter\[3\] _0671_ _0672_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2224_ tt_um_rejunity_ay8913.tone_A_generator.period\[6\] _0731_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_51_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2086_ _0607_ _0572_ _0605_ _0523_ _1082_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1939_ tt_um_rejunity_ay8913.noise_generator.lfsr\[13\] _0480_ _0483_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1508__A2 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1683__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1724_ _0300_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1655_ _1100_ _1187_ _1188_ tt_um_rejunity_ay8913.envelope_generator.period\[13\]
+ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1586_ tt_um_rejunity_ay8913.pwm_B.accumulator\[3\] _1140_ _1078_ _1143_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_53_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2138_ _0657_ _0646_ _0625_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2069_ _0553_ _0589_ tt_um_rejunity_ay8913.tone_C_generator.counter\[7\] _0595_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2207_ _0706_ _0713_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1371_ net8 _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1440_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\] tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
+ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_18_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1638_ _1177_ _1174_ _1178_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1707_ _1176_ _0282_ _0284_ tt_um_rejunity_ay8913.noise_disable_B _0290_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1569_ _1002_ _1048_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1647__A1 _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2541_ _0155_ clknet_leaf_18_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2472_ _0086_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2610_ _0224_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1285_ blink.counter\[14\] _0921_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1354_ _0972_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1423_ _1027_ _1025_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_13_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_13_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_38_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ _1086_ _0508_ _0510_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2455_ _0069_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2524_ _0138_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2386_ _0000_ clknet_leaf_7_wb_clk_i blink.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1268_ _0892_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1337_ _0955_ _0954_ _0958_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1406_ _1013_ _0871_ _0872_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1199_ _0848_ _0852_ _0849_ net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_46_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2171_ tt_um_rejunity_ay8913.tone_B_generator.counter\[7\] _0643_ _0679_ _0684_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_48_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2240_ _0746_ _0735_ _0714_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_31_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1955_ tt_um_rejunity_ay8913.noise_generator.lfsr\[16\] _0440_ _1161_ _0496_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1886_ _0442_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2507_ _0121_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2438_ _0052_ clknet_leaf_28_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2369_ _0988_ _0836_ _0837_ _0853_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_54_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1740_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\] _0315_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1671_ net6 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input8_I io_in_1[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2190__A3 _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2154_ _0627_ _0666_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2085_ _0391_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2223_ tt_um_rejunity_ay8913.tone_A_generator.period\[7\] _0730_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_51_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1869_ _0386_ _0428_ _0429_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1938_ tt_um_rejunity_ay8913.noise_generator.lfsr\[14\] _0475_ _0482_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1654_ _1189_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_38_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_38_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1723_ _0293_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1585_ tt_um_rejunity_ay8913.pwm_B.accumulator\[3\] _1140_ _1142_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2206_ _0708_ _0712_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2137_ _0655_ _0656_ _0644_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2068_ tt_um_rejunity_ay8913.tone_C_generator.counter\[7\] _0553_ _0589_ _0594_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_54_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1370_ _0985_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1637_ _1114_ tt_um_rejunity_ay8913.envelope_A _1174_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_18_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1706_ _0289_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1568_ _1050_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1499_ _1082_ _1083_ _1084_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2540_ _0154_ clknet_leaf_18_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2471_ _0085_ clknet_leaf_14_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1422_ _1027_ _1025_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1284_ _0910_ _0920_ _0921_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1353_ _0967_ _0971_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_38_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2045__A2 _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1556__A1 _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1971_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\] _0382_ _0510_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1668__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2454_ _0068_ clknet_leaf_14_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1405_ _0871_ _0872_ _1013_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2385_ _0846_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2523_ _0137_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.restart_envelope vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput1 custom_settings[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1267_ _0906_ _0909_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1336_ blink.counter\[29\] _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1198_ tt_um_rejunity_ay8913.pwm_master.accumulator\[10\] _0852_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1529__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2170_ _0683_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_48_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1701__A1 _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1954_ _0443_ _0494_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1885_ tt_um_rejunity_ay8913.noise_generator.signal_edge.signal _0438_ _0442_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2506_ _0120_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2437_ _0051_ clknet_leaf_28_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2368_ _1052_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1319_ _0934_ _0943_ _0945_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2299_ _0788_ _0789_ _0791_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1670_ _0267_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2222_ _0718_ _0720_ _0728_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2153_ _0670_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2084_ _0606_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1937_ _0479_ _0481_ _0478_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1868_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\] _0425_ _0356_
+ _0422_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1799_ _0320_ tt_um_rejunity_ay8913.envelope_generator.period\[0\] tt_um_rejunity_ay8913.envelope_generator.period\[2\]
+ _0324_ _0367_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_31_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_8_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_8_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_32_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ _0986_ _1187_ _1188_ tt_um_rejunity_ay8913.envelope_generator.period\[12\]
+ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1584_ _1140_ _1141_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1722_ _0294_ _0301_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2205_ tt_um_rejunity_ay8913.tone_A_generator.counter\[10\] _0709_ _0710_ _0711_
+ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2136_ _0645_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2067_ _0593_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2191__B _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2378__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2302__A1 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1705_ _0270_ _0283_ _0285_ tt_um_rejunity_ay8913.noise_disable_A _0289_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1567_ _1130_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1636_ _1176_ _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2119_ _0635_ _0638_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1498_ tt_um_rejunity_ay8913.pwm_C.accumulator\[6\] tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
+ _1076_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1804__B1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2470_ _0084_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1421_ tt_um_rejunity_ay8913.pwm_master.accumulator\[6\] _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1283_ blink.counter\[13\] _0919_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1352_ _0968_ tt_um_rejunity_ay8913.latched_register\[0\] _0970_ _0971_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xclkbuf_leaf_22_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_22_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2599_ _0213_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1619_ tt_um_rejunity_ay8913.pwm_A.accumulator\[6\] _1163_ _1165_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_52_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1970_ _0278_ _0509_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2522_ _0136_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.noise_disable_C vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1335_ _0949_ _0956_ _0957_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2453_ _0067_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1404_ tt_um_rejunity_ay8913.pwm_master.accumulator\[3\] _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2384_ _0270_ _0292_ _0842_ tt_um_rejunity_ay8913.envelope_continue _0846_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput2 custom_settings[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1266_ blink.counter\[8\] _0908_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1197_ _0848_ _0851_ _0849_ net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_34_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1465__A1 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1953_ tt_um_rejunity_ay8913.noise_generator.lfsr\[3\] _0864_ _0493_ _0494_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1884_ tt_um_rejunity_ay8913.noise_generator.lfsr\[1\] _0440_ _0441_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2193__A2 _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2505_ _0119_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1318_ _0944_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2436_ _0050_ clknet_leaf_28_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2298_ _0788_ _0789_ _0790_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2367_ _0971_ _1173_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1249_ blink.counter\[3\] blink.counter\[2\] blink.counter\[1\] blink.counter\[0\]
+ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_19_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2152_ _0664_ _0669_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2221_ _0724_ _0727_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2083_ _0575_ _0604_ _0605_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_33_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1438__A1 _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1867_ _0425_ _0424_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
+ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_51_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1936_ tt_um_rejunity_ay8913.noise_generator.lfsr\[12\] _0480_ _0481_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1798_ _0314_ _0330_ _0319_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2419_ _0033_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1721_ _0295_ _0300_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1652_ _1181_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2148__A2 _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1583_ tt_um_rejunity_ay8913.pwm_B.accumulator\[2\] _0870_ _1078_ _1141_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1659__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2135_ tt_um_rejunity_ay8913.tone_B_generator.counter\[5\] _0651_ _0635_ _0654_ _0655_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2204_ tt_um_rejunity_ay8913.tone_A_generator.counter\[9\] _0711_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2066_ _0587_ _0592_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1919_ tt_um_rejunity_ay8913.noise_generator.lfsr\[9\] _0464_ _0468_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1704_ _0288_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1566_ _1104_ _1125_ _1126_ tt_um_rejunity_ay8913.tone_B_generator.period\[7\] _1130_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1635_ net8 _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1497_ tt_um_rejunity_ay8913.pwm_C.accumulator\[6\] _1077_ tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
+ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2118_ tt_um_rejunity_ay8913.tone_B_generator.counter\[3\] _0636_ _0637_ tt_um_rejunity_ay8913.tone_B_generator.counter\[4\]
+ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2049_ _0574_ _0579_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_32_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ _1024_ _1022_ _1026_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1351_ tt_um_rejunity_ay8913.active _0969_ net12 net14 _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1282_ blink.counter\[13\] _0919_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1618_ _1163_ _1164_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1549_ _1119_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2598_ _0212_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ _0135_ clknet_leaf_32_wb_clk_i tt_um_rejunity_ay8913.noise_disable_B vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1265_ _0893_ _0907_ _0908_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1334_ _0955_ _0953_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1403_ _1011_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2452_ _0066_ clknet_leaf_37_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2383_ _0845_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput3 custom_settings[3] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1196_ tt_um_rejunity_ay8913.pwm_C.accumulator\[9\] _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1883_ _0439_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1952_ _0488_ _0492_ tt_um_rejunity_ay8913.noise_generator.lfsr\[3\] _0864_ _0493_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2504_ _0118_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2435_ _0049_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1248_ blink.counter\[3\] _0894_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1317_ blink.counter\[24\] _0942_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2366_ _0835_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2297_ _1051_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_54_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2151_ _0627_ _0666_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2082_ tt_um_rejunity_ay8913.tone_C_generator.counter\[10\] _0532_ _0600_ _0605_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2220_ tt_um_rejunity_ay8913.tone_A_generator.counter\[3\] _0725_ _0726_ tt_um_rejunity_ay8913.tone_A_generator.counter\[4\]
+ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1866_ _0386_ _0426_ _0427_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1797_ _0335_ _0366_ _0367_ _0371_ _0353_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1935_ _0442_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2418_ _0032_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input14_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2349_ _0260_ _0823_ _0825_ tt_um_rejunity_ay8913.envelope_generator.period\[0\]
+ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ _1179_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_13_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1720_ _0297_ _0299_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1582_ tt_um_rejunity_ay8913.pwm_B.accumulator\[2\] _0870_ _1140_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2134_ _0629_ _0653_ _0638_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2065_ _0553_ _0589_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input6_I io_in_1[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2203_ tt_um_rejunity_ay8913.tone_A_generator.period\[9\] _0710_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_16_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_16_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1849_ _0332_ _0415_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1918_ _0465_ _0466_ _0467_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_4_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1510__A1 _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1634_ _0989_ _1174_ _1175_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1703_ _0268_ _0283_ _0285_ tt_um_rejunity_ay8913.tone_disable_C _0288_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1565_ _1129_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1496_ _1011_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2117_ tt_um_rejunity_ay8913.tone_B_generator.period\[4\] _0637_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2048_ _0537_ _0576_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1281_ _0910_ _0918_ _0919_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1350_ net13 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_46_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2597_ _0211_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1617_ tt_um_rejunity_ay8913.pwm_A.accumulator\[5\] _1160_ _1161_ _1164_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1970__A1 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1548_ _1054_ _1117_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1479_ tt_um_rejunity_ay8913.pwm_C.accumulator\[2\] _0860_ _1070_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_31_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_31_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1713__A1 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1477__B1 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2451_ _0065_ clknet_leaf_37_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2520_ _0134_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.noise_disable_A vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1402_ _1010_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1264_ blink.counter\[7\] _0905_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1333_ _0955_ _0954_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput4 io_in_1[0] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2382_ _0268_ _0137_ _0842_ tt_um_rejunity_ay8913.envelope_attack _0845_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1195_ _0848_ _0850_ _0849_ net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1882_ tt_um_rejunity_ay8913.noise_generator.signal_edge.signal _0438_ _0439_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1951_ tt_um_rejunity_ay8913.noise_generator.lfsr\[4\] tt_um_rejunity_ay8913.noise_generator.lfsr\[2\]
+ tt_um_rejunity_ay8913.noise_generator.lfsr\[1\] _0491_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_2503_ _0117_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2365_ net11 _0830_ _0831_ tt_um_rejunity_ay8913.envelope_generator.period\[7\] _0835_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2434_ _0048_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1247_ _0893_ _0894_ _0895_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_47_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1316_ blink.counter\[24\] _0942_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2296_ tt_um_rejunity_ay8913.clk_counter\[1\] _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1392__A2 tt_um_rejunity_ay8913.tone_C_generator.period\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2150_ _0668_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2081_ _0525_ _0602_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1934_ tt_um_rejunity_ay8913.noise_generator.lfsr\[13\] _0475_ _0479_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1865_ _0425_ _0424_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1796_ _0370_ _0350_ _0355_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2417_ _0031_ clknet_leaf_4_wb_clk_i blink.counter\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2348_ _0824_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2323__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2279_ _0766_ _0777_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_50_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1650_ _1186_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1581_ _1133_ _1139_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_13_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2202_ tt_um_rejunity_ay8913.tone_A_generator.period\[10\] _0709_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2133_ tt_um_rejunity_ay8913.tone_B_generator.counter\[2\] _0648_ _0652_ _0631_ _0653_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2064_ _0591_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1917_ _0446_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1779_ _0352_ tt_um_rejunity_ay8913.envelope_generator.period\[15\] _0354_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1848_ _0413_ _0412_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1564_ _1102_ _1125_ _1126_ tt_um_rejunity_ay8913.tone_B_generator.period\[6\] _1129_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ _1114_ tt_um_rejunity_ay8913.amplitude_A\[0\] _1174_ _1175_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1702_ _0287_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1495_ tt_um_rejunity_ay8913.pwm_C.accumulator\[6\] _1077_ _1081_ _0064_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2116_ tt_um_rejunity_ay8913.tone_B_generator.period\[3\] _0636_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2047_ _0578_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_1_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1280_ blink.counter\[12\] blink.counter\[11\] blink.counter\[10\] _0912_ _0919_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_46_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ _1117_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1616_ tt_um_rejunity_ay8913.pwm_A.accumulator\[5\] _1160_ _1163_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2596_ _0210_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.tone_B vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1478_ _1065_ _1069_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1889__I _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_39_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1401_ _0974_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2450_ _0064_ clknet_leaf_37_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2381_ _0844_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1263_ blink.counter\[7\] _0905_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1332_ blink.counter\[28\] _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 io_in_1[1] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1194_ tt_um_rejunity_ay8913.pwm_B.accumulator\[9\] _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2579_ _0193_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1950_ _0489_ _0490_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2502_ _0116_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1881_ tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0
+ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2364_ _0834_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1315_ _0934_ _0941_ _0942_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2433_ _0047_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1246_ blink.counter\[1\] _0874_ blink.counter\[2\] _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2295_ _0788_ _0447_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1604__A1 _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2080_ _0603_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1933_ _0476_ _0477_ _0478_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1864_ _0425_ _0424_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1795_ _0369_ _0358_ _0361_ _0338_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_3_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2416_ _0030_ clknet_leaf_4_wb_clk_i blink.counter\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2347_ _0976_ _0822_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2278_ tt_um_rejunity_ay8913.tone_A_generator.counter\[8\] _0773_ _0777_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1229_ _0878_ _0879_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2087__A1 _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1580_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\] _1137_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
+ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2132_ _0630_ tt_um_rejunity_ay8913.tone_B_generator.period\[1\] _0652_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2201_ _0707_ tt_um_rejunity_ay8913.tone_A_generator.period\[9\] tt_um_rejunity_ay8913.tone_A_generator.period\[8\]
+ _0701_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_21_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2063_ _0587_ _0590_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_44_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1847_ _0404_ _0414_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1916_ tt_um_rejunity_ay8913.noise_generator.lfsr\[7\] _0458_ _0466_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1778_ _0352_ tt_um_rejunity_ay8913.envelope_generator.period\[15\] _0353_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_25_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_25_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_4_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_3__f_wb_clk_i clknet_0_wb_clk_i clknet_2_3__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1701_ _0266_ _0283_ _0285_ tt_um_rejunity_ay8913.tone_disable_B _0287_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1563_ _1128_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1494_ tt_um_rejunity_ay8913.pwm_C.accumulator\[6\] _1077_ _1080_ _1081_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1632_ _1088_ _1173_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2115_ _0632_ tt_um_rejunity_ay8913.tone_B_generator.period\[5\] tt_um_rejunity_ay8913.tone_B_generator.period\[4\]
+ _0634_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_1_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2046_ _0575_ _0576_ _0577_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_13_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1192__A1 blink.LED vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2595_ _0209_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1477_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\] _1044_ _1057_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\]
+ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1615_ _1160_ _1162_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1546_ _0971_ _1107_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_37_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2029_ _0540_ tt_um_rejunity_ay8913.tone_C_generator.period\[1\] _0562_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_40_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_40_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1331_ _0949_ _0952_ _0954_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1400_ tt_um_rejunity_ay8913.pwm_master.accumulator\[2\] net20 _1009_ _0041_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2380_ _0266_ _0137_ _0842_ tt_um_rejunity_ay8913.envelope_alternate _0844_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1262_ _0902_ _0903_ _0905_ _0906_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1193_ _0847_ _0848_ _0849_ net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput6 io_in_1[2] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1529_ _1104_ _1097_ _1098_ tt_um_rejunity_ay8913.tone_C_generator.period\[7\] _1105_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2578_ _0192_ clknet_leaf_8_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_40_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ tt_um_rejunity_ay8913.envelope_attack _0302_ _0436_ _0437_ _0160_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2501_ _0115_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_47_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1314_ blink.counter\[23\] blink.counter\[19\] _0882_ _0931_ _0942_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2363_ net10 _0830_ _0831_ tt_um_rejunity_ay8913.envelope_generator.period\[6\] _0834_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2432_ _0046_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2294_ tt_um_rejunity_ay8913.clk_counter\[0\] _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_56_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1245_ blink.counter\[2\] blink.counter\[1\] _0874_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1863_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\] _0425_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1932_ _0446_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1794_ _0368_ _0359_ _0360_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2415_ _0029_ clknet_leaf_4_wb_clk_i blink.counter\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1228_ blink.counter\[16\] blink.counter\[15\] blink.counter\[14\] blink.counter\[13\]
+ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_2346_ _0822_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2277_ _0776_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_2_2__f_wb_clk_i clknet_0_wb_clk_i clknet_2_2__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2087__A2 _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1399__B _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2250__A2 _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1210__B1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2131_ tt_um_rejunity_ay8913.tone_B_generator.period\[5\] _0651_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2062_ _0588_ _0589_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2200_ tt_um_rejunity_ay8913.tone_A_generator.counter\[9\] _0707_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1777_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\] _0352_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1846_ _0413_ _0412_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1915_ tt_um_rejunity_ay8913.noise_generator.lfsr\[8\] _0464_ _0465_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input12_I io_in_2[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2329_ net7 _0804_ _1134_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1700_ _0286_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1631_ _1172_ _1106_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1562_ _1100_ _1125_ _1126_ tt_um_rejunity_ay8913.tone_B_generator.period\[5\] _1128_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1493_ _1007_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2114_ _0633_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2045_ _0519_ _0395_ _0540_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input4_I io_in_1[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1829_ _0394_ _0400_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1192__A2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2594_ _0208_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1614_ tt_um_rejunity_ay8913.pwm_A.accumulator\[4\] _1158_ _1161_ _1162_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1707__A1 _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1545_ _1005_ _1110_ _1116_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1476_ _1065_ _1068_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2380__A1 _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2028_ tt_um_rejunity_ay8913.tone_C_generator.period\[5\] _0561_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_37_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1261_ _0892_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1330_ _0953_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1192_ blink.LED net3 _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput7 io_in_1[3] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2577_ _0191_ clknet_leaf_8_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2353__A1 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1528_ net11 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1459_ _1057_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2344__A1 _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2500_ _0114_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2431_ _0045_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1244_ _0892_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_2_1__f_wb_clk_i clknet_0_wb_clk_i clknet_2_1__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2362_ _0833_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1313_ blink.counter\[23\] _0940_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2293_ _0786_ _0787_ _1086_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_19_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_19_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2629_ _0243_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2317__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1862_ _0409_ _0423_ _0424_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1793_ _0342_ _0343_ _0344_ _0345_ _0341_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xinput10 io_in_1[6] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1931_ tt_um_rejunity_ay8913.noise_generator.lfsr\[11\] _0469_ _0477_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2414_ _0028_ clknet_leaf_6_wb_clk_i blink.counter\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1952__C _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1227_ blink.counter\[11\] _0877_ blink.counter\[9\] blink.counter\[12\] _0878_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2276_ _0766_ _0775_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2345_ _1108_ _1173_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_50_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2304__B _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1210__A1 tt_um_rejunity_ay8913.noise_generator.lfsr\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2061_ tt_um_rejunity_ay8913.tone_C_generator.counter\[5\] _0543_ tt_um_rejunity_ay8913.tone_C_generator.counter\[3\]
+ _0581_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2130_ _0632_ tt_um_rejunity_ay8913.tone_B_generator.period\[5\] _0647_ _0649_ _0650_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_28_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1914_ _0452_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1776_ _0338_ _0341_ _0346_ _0350_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1845_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\] _0413_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2328_ _0966_ _0808_ _0811_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2085__I _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2259_ _0762_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_34_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_34_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1630_ tt_um_rejunity_ay8913.latched_register\[3\] _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1561_ _1127_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1492_ _1077_ _1079_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2113_ tt_um_rejunity_ay8913.tone_B_generator.counter\[4\] _0633_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2044_ tt_um_rejunity_ay8913.tone_C_generator.counter\[1\] tt_um_rejunity_ay8913.tone_C_generator.counter\[0\]
+ _0387_ _0388_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_1_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\] _0398_ _0400_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1759_ _0332_ _0333_ _0312_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\]
+ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1973__A2 _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2593_ _0207_ clknet_leaf_11_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1544_ _1114_ tt_um_rejunity_ay8913.tone_B_generator.period\[11\] _1111_ _1116_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1613_ _1007_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1475_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\] _1062_ _1063_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\]
+ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1643__A1 _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ _0542_ tt_um_rejunity_ay8913.tone_C_generator.period\[5\] _0557_ _0559_ _0560_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_37_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1882__A1 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1260_ _0897_ _0904_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1191_ net3 _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput8 io_in_1[4] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_2_0__f_wb_clk_i clknet_0_wb_clk_i clknet_2_0__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_34_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1527_ _1103_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2576_ _0190_ clknet_leaf_8_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_2_1__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1458_ _1050_ _1042_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1389_ net6 _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_56_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2361_ net9 _0830_ _0831_ tt_um_rejunity_ay8913.envelope_generator.period\[5\] _0833_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2430_ _0044_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1243_ _0887_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1312_ _0934_ _0939_ _0940_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2292_ tt_um_rejunity_ay8913.tone_A _0520_ _0751_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2628_ _0242_ clknet_leaf_21_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2559_ _0173_ clknet_leaf_41_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2317__A2 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ tt_um_rejunity_ay8913.noise_generator.lfsr\[12\] _0475_ _0476_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1861_ _0356_ _0422_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1792_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\] _0333_ _0367_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput11 io_in_1[7] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2413_ _0027_ clknet_leaf_4_wb_clk_i blink.counter\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2344_ _1005_ _0815_ _0821_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1226_ blink.counter\[10\] _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1819__A1 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2275_ _0773_ _0774_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_50_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_4_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2060_ _0543_ _0584_ tt_um_rejunity_ay8913.tone_C_generator.counter\[5\] _0588_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1913_ _0462_ _0463_ _0456_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1775_ _0347_ _0348_ _0349_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
+ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1844_ _0409_ _0410_ _0412_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_8_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2258_ _0753_ _0761_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_4_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2327_ net6 _0805_ _1134_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1209_ tt_um_rejunity_ay8913.amplitude_B\[0\] tt_um_rejunity_ay8913.envelope_B tt_um_rejunity_ay8913.tone_disable_B
+ tt_um_rejunity_ay8913.tone_B _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2189_ _0513_ _0662_ tt_um_rejunity_ay8913.tone_B _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1560_ _0986_ _1125_ _1126_ tt_um_rejunity_ay8913.tone_B_generator.period\[4\] _1127_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2112_ tt_um_rejunity_ay8913.tone_B_generator.counter\[5\] _0632_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1491_ tt_um_rejunity_ay8913.pwm_C.accumulator\[5\] _1074_ _1078_ _1079_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1355__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2043_ _0573_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1827_ _0394_ _0399_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1758_ tt_um_rejunity_ay8913.envelope_generator.period\[7\] _0333_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1689_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\] _0279_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2592_ _0206_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1543_ _1001_ _1110_ _1115_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1612_ tt_um_rejunity_ay8913.pwm_A.accumulator\[4\] _1158_ _1160_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1474_ _1065_ _1067_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2026_ _0519_ tt_um_rejunity_ay8913.tone_C_generator.period\[0\] tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
+ _0540_ tt_um_rejunity_ay8913.tone_C_generator.counter\[2\] _0558_ _0559_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_37_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 io_in_1[5] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1190_ tt_um_rejunity_ay8913.pwm_A.accumulator\[9\] _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_34_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1526_ _1102_ _1097_ _1098_ tt_um_rejunity_ay8913.tone_C_generator.period\[6\] _1103_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2575_ _0189_ clknet_leaf_9_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1457_ _1055_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1388_ _0999_ _0993_ _1000_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2009_ tt_um_rejunity_ay8913.tone_C_generator.counter\[5\] _0542_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1552__A1 _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1607__A2 _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_ay8913_40 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _0832_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1311_ _0882_ _0932_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2291_ _0513_ _0751_ tt_um_rejunity_ay8913.tone_A _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1242_ _0890_ _0891_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2143__B _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2627_ _0241_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_28_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_28_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1509_ _1091_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2489_ _0103_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2558_ _0172_ clknet_leaf_41_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_43_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1860_ _0356_ _0422_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 io_in_2[0] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1791_ _0365_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1516__A1 _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2412_ _0026_ clknet_leaf_4_wb_clk_i blink.counter\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1307__B _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2274_ _0732_ _0768_ tt_um_rejunity_ay8913.tone_A_generator.counter\[7\] _0774_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2343_ _0816_ tt_um_rejunity_ay8913.tone_A_generator.period\[11\] _0817_ _0821_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1225_ blink.counter\[17\] _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1989_ tt_um_rejunity_ay8913.tone_C_generator.counter\[8\] _0522_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ _0411_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1912_ tt_um_rejunity_ay8913.noise_generator.lfsr\[6\] _0458_ _0463_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1774_ tt_um_rejunity_ay8913.envelope_generator.period\[13\] _0349_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2257_ tt_um_rejunity_ay8913.tone_A_generator.counter\[3\] _0760_ _0761_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1208_ tt_um_rejunity_ay8913.noise_disable_B _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2326_ _0968_ _0808_ _0810_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2188_ _0607_ _0662_ _0695_ _0613_ _1055_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_31_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1490_ _0995_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1636__I _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2111_ _0610_ tt_um_rejunity_ay8913.tone_B_generator.period\[0\] tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
+ _0630_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2042_ _0521_ _0574_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1826_ _0396_ _0398_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1757_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\] _0332_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1688_ _0278_ _1042_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input10_I io_in_1[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2309_ _0797_ _0798_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_0_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1456__I _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1191__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1611_ _1158_ _1159_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2591_ _0205_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1542_ _1114_ tt_um_rejunity_ay8913.tone_B_generator.period\[10\] _1111_ _1115_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1473_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\] _1062_ _1063_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\]
+ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input2_I custom_settings[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2025_ tt_um_rejunity_ay8913.tone_C_generator.period\[2\] _0558_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_37_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1809_ _0311_ _0383_ _0302_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2347__A1 _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_34_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2574_ _0188_ clknet_leaf_8_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1525_ net10 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1387_ _0996_ tt_um_rejunity_ay8913.tone_C_generator.period\[9\] _0997_ _1000_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1456_ _1054_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2008_ _0519_ tt_um_rejunity_ay8913.tone_C_generator.period\[0\] tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
+ _0540_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_37_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2329__A1 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_ay8913_30 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_41 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_36_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1241_ blink.counter\[1\] _0874_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1310_ blink.counter\[21\] _0936_ blink.counter\[22\] _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2290_ _0607_ _0751_ _0784_ _0702_ _1055_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _0171_ clknet_leaf_41_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2626_ _0240_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1508_ _1054_ _1089_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2488_ _0102_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1439_ _1040_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 io_in_2[1] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ _0351_ _0364_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1461__A1 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2411_ _0025_ clknet_leaf_3_wb_clk_i blink.counter\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1374__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1224_ blink.counter\[31\] _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2273_ tt_um_rejunity_ay8913.tone_A_generator.counter\[7\] _0732_ _0768_ _0773_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2342_ _1001_ _0815_ _0820_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1988_ _0519_ _0520_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2609_ _0223_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_A vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1459__I _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1773_ tt_um_rejunity_ay8913.envelope_generator.period\[14\] _0348_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1842_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\] tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\]
+ _0401_ _0402_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_12_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1911_ tt_um_rejunity_ay8913.noise_generator.lfsr\[7\] _0453_ _0462_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2187_ _0696_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2256_ _0716_ _0755_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1207_ _0856_ _0859_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2325_ net5 _0805_ _0790_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_12_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_12_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1664__A1 _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2110_ tt_um_rejunity_ay8913.tone_B_generator.counter\[1\] _0630_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2041_ _0573_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1655__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1825_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\] tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\]
+ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1756_ _0316_ _0328_ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2308_ tt_um_rejunity_ay8913.clk_counter\[4\] _0794_ _1008_ _0798_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1687_ _1134_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2239_ _0744_ _0745_ _0733_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1885__A1 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2590_ _0204_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1610_ tt_um_rejunity_ay8913.pwm_A.accumulator\[3\] _1156_ _1147_ _1159_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1472_ _1065_ _1066_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1541_ _1002_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2024_ _0554_ _0555_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1628__A1 _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1739_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\] _0312_ _0313_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\]
+ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1808_ _0372_ _0377_ _0382_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_51_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1467__I _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1524_ _1101_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2573_ _0187_ clknet_leaf_11_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2642_ _0256_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.envelope_continue vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1455_ _0975_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1386_ net5 _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2007_ tt_um_rejunity_ay8913.tone_C_generator.counter\[1\] _0540_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_9_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_ay8913_42 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_31 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_51_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1240_ _0874_ _0890_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1507_ _1089_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2487_ _0101_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _0239_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2556_ _0170_ clknet_leaf_41_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1369_ _0984_ _0973_ _0978_ tt_um_rejunity_ay8913.noise_generator.period\[3\] _0985_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1438_ _1021_ tt_um_rejunity_ay8913.pwm_master.accumulator\[8\] tt_um_rejunity_ay8913.pwm_master.accumulator\[9\]
+ _1033_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xclkbuf_leaf_37_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_37_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 rst_n net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2410_ _0024_ clknet_leaf_3_wb_clk_i blink.counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2341_ _0816_ tt_um_rejunity_ay8913.tone_A_generator.period\[10\] _0817_ _0820_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1223_ blink.counter\[0\] _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2272_ _0772_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1987_ _0397_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2539_ _0153_ clknet_leaf_18_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2608_ _0222_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1910_ _0460_ _0461_ _0456_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1772_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\] _0347_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1841_ _0329_ _0407_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_8_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2324_ _0990_ _0808_ _0809_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2186_ _0665_ _0694_ _0695_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2255_ _0759_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1206_ tt_um_rejunity_ay8913.envelope_C _0857_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2040_ _0397_ _0572_ _1010_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1755_ _0329_ tt_um_rejunity_ay8913.envelope_generator.period\[5\] tt_um_rejunity_ay8913.envelope_generator.period\[4\]
+ _0315_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1824_ _0389_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1686_ _0277_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2238_ _0734_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2307_ _0796_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2169_ _0677_ _0682_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1540_ _0999_ _1110_ _1113_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1471_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\] _1062_ _1063_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\]
+ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2023_ tt_um_rejunity_ay8913.tone_C_generator.counter\[7\] _0551_ _0556_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1807_ _0379_ _0381_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1564__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1738_ tt_um_rejunity_ay8913.envelope_generator.period\[5\] _0313_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1669_ _0266_ _0262_ _0264_ tt_um_rejunity_ay8913.tone_A_generator.period\[1\] _0267_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2292__A2 _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1432__B _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1523_ _1100_ _1097_ _1098_ tt_um_rejunity_ay8913.tone_C_generator.period\[5\] _1101_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2572_ _0186_ clknet_leaf_11_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1454_ _1046_ _1047_ _1049_ _1053_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2641_ _0255_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.envelope_attack vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1385_ _0989_ _0993_ _0998_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2006_ _0538_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_ay8913_32 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_leaf_7_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_7_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_30_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2624_ _0238_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1506_ _0967_ _1088_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2486_ _0100_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1437_ _1037_ _1039_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2555_ _0169_ clknet_leaf_42_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1299_ _0923_ _0930_ _0931_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1368_ net7 _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2271_ _0766_ _0771_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1671__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2340_ _0999_ _0815_ _0819_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1222_ _0873_ net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1986_ tt_um_rejunity_ay8913.tone_C_generator.counter\[0\] _0519_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_30_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2607_ _0221_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2469_ _0083_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2538_ _0152_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_6_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1840_ _0385_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_29_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1771_ _0342_ _0343_ _0344_ _0345_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2254_ _0753_ _0758_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2323_ net4 _0805_ _0790_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2185_ tt_um_rejunity_ay8913.tone_B_generator.counter\[10\] _0622_ _0690_ _0695_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1205_ tt_um_rejunity_ay8913.tone_C tt_um_rejunity_ay8913.tone_disable_C _0858_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ tt_um_rejunity_ay8913.noise_generator.signal_edge.signal _0508_ _0509_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_21_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_21_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1823_ _0320_ _0395_ _0323_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1754_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\] _0329_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1685_ _1104_ _0272_ _0273_ tt_um_rejunity_ay8913.tone_A_generator.period\[7\] _0277_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2237_ tt_um_rejunity_ay8913.tone_A_generator.counter\[5\] _0740_ _0724_ _0743_ _0744_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2306_ tt_um_rejunity_ay8913.clk_counter\[4\] _0794_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2168_ _0643_ _0679_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2099_ _0618_ tt_um_rejunity_ay8913.tone_B_generator.period\[9\] tt_um_rejunity_ay8913.tone_B_generator.period\[8\]
+ _0612_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_0_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2359__A1 _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1470_ _1055_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2022_ tt_um_rejunity_ay8913.tone_C_generator.counter\[6\] _0552_ _0555_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1806_ net2 _0378_ _0380_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1737_ tt_um_rejunity_ay8913.envelope_generator.period\[6\] _0312_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1668_ net5 _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1599_ tt_um_rejunity_ay8913.pwm_B.accumulator\[7\] _1150_ _1080_ _1152_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2044__A3 _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2292__A3 _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2640_ _0254_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.envelope_alternate vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2571_ _0185_ clknet_leaf_11_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1522_ net9 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1453_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\] _1050_ _1042_ _1052_ _1053_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1674__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2005_ _0536_ tt_um_rejunity_ay8913.tone_C_generator.period\[3\] tt_um_rejunity_ay8913.tone_C_generator.period\[2\]
+ _0537_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1384_ _0996_ tt_um_rejunity_ay8913.tone_C_generator.period\[8\] _0997_ _0998_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_33_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_ay8913_33 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_47_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_22_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2623_ _0237_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2554_ _0168_ clknet_leaf_42_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1367_ _0983_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1436_ tt_um_rejunity_ay8913.pwm_master.accumulator\[9\] _1038_ _1039_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2485_ _0099_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1505_ tt_um_rejunity_ay8913.latched_register\[1\] tt_um_rejunity_ay8913.latched_register\[0\]
+ _0970_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1298_ blink.counter\[18\] blink.counter\[17\] blink.counter\[16\] _0925_ _0931_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2270_ _0732_ _0768_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1221_ _0871_ _0872_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1685__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1437__A1 _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1988__A2 _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1985_ _0311_ _0294_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2537_ _0151_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2606_ _0220_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2468_ _0082_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2399_ _0013_ clknet_leaf_5_wb_clk_i blink.counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1419_ _0996_ _1025_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2089__B _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1419__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1770_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\] _0345_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2184_ _0615_ _0692_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2253_ _0716_ _0755_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2322_ _0804_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_25_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1204_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\] tt_um_rejunity_ay8913.envelope_generator.invert_output
+ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1968_ _0504_ _0506_ _0507_ _0397_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1899_ _0452_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1649__A1 _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1888__A1 _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1822_ _0382_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1753_ _0319_ _0326_ _0327_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1684_ _0276_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2167_ _0681_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2236_ _0718_ _0742_ _0727_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2305_ _0794_ _0795_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2098_ tt_um_rejunity_ay8913.tone_B_generator.counter\[9\] _0618_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2086__C _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2021_ tt_um_rejunity_ay8913.tone_C_generator.counter\[7\] _0551_ _0552_ _0553_ _0554_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1805_ tt_um_rejunity_ay8913.clk_counter\[3\] tt_um_rejunity_ay8913.clk_counter\[5\]
+ tt_um_rejunity_ay8913.clk_counter\[4\] tt_um_rejunity_ay8913.clk_counter\[6\] _0380_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_1736_ _0296_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1667_ _0265_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1598_ _1150_ _1151_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2219_ tt_um_rejunity_ay8913.tone_A_generator.period\[4\] _0726_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2044__A4 _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2570_ _0184_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1521_ _1099_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1452_ _1051_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1383_ _0992_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ tt_um_rejunity_ay8913.tone_C_generator.counter\[2\] _0537_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_45_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1719_ _0298_ tt_um_rejunity_ay8913.envelope_generator.hold tt_um_rejunity_ay8913.envelope_generator.stop
+ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_56_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_ay8913_34 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_51_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2622_ _0236_ clknet_leaf_42_wb_clk_i blink.LED vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1504_ _1087_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2553_ _0167_ clknet_leaf_42_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1366_ _0982_ _0973_ _0978_ tt_um_rejunity_ay8913.noise_generator.period\[2\] _0983_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2484_ _0098_ clknet_leaf_37_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1435_ tt_um_rejunity_ay8913.pwm_master.accumulator\[8\] _1032_ _1038_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1297_ _0876_ _0927_ blink.counter\[18\] _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_15_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_15_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1220_ _0856_ _0859_ _0870_ _0867_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_1984_ _0505_ _0518_ _0511_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2467_ _0081_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2536_ _0150_ clknet_leaf_18_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2605_ _0219_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2398_ _0012_ clknet_leaf_8_wb_clk_i blink.counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1418_ _1018_ _1017_ tt_um_rejunity_ay8913.pwm_master.accumulator\[4\] tt_um_rejunity_ay8913.pwm_master.accumulator\[5\]
+ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1349_ tt_um_rejunity_ay8913.latched_register\[1\] _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_29_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2147__A3 _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2321_ _0805_ _0807_ _1037_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2183_ _0693_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2252_ _0757_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1203_ _0853_ _0854_ _0855_ tt_um_rejunity_ay8913.noise_generator.lfsr\[0\] _0856_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_18_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _0505_ tt_um_rejunity_ay8913.noise_generator.period\[4\] _0507_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1898_ _0439_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2519_ _0133_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_disable_C vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_30_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_30_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_29_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1821_ _0385_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1752_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\] _0317_ _0327_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1683_ _1102_ _0272_ _0273_ tt_um_rejunity_ay8913.tone_A_generator.period\[6\] _0276_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2304_ tt_um_rejunity_ay8913.clk_counter\[3\] _0793_ _1008_ _0795_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2166_ _0677_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2097_ _0612_ tt_um_rejunity_ay8913.tone_B_generator.period\[8\] _0614_ _0616_ _0617_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2235_ tt_um_rejunity_ay8913.tone_A_generator.counter\[2\] _0737_ _0741_ _0720_ _0742_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_0_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2295__A2 _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2020_ tt_um_rejunity_ay8913.tone_C_generator.counter\[6\] _0553_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2293__B _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1666_ _0260_ _0262_ _0264_ tt_um_rejunity_ay8913.tone_A_generator.period\[0\] _0265_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1804_ tt_um_rejunity_ay8913.clk_counter\[0\] tt_um_rejunity_ay8913.clk_counter\[1\]
+ tt_um_rejunity_ay8913.clk_counter\[2\] net2 _0378_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_13_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1735_ _0302_ _0310_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1597_ tt_um_rejunity_ay8913.pwm_B.accumulator\[6\] _1146_ _1147_ _1151_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2149_ _0665_ _0666_ _0667_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_36_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2218_ tt_um_rejunity_ay8913.tone_A_generator.period\[3\] _0725_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1520_ _0986_ _1097_ _1098_ tt_um_rejunity_ay8913.tone_C_generator.period\[4\] _1099_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1451_ _0994_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1382_ _0995_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1703__A1 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2003_ tt_um_rejunity_ay8913.tone_C_generator.counter\[3\] _0536_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1211__I tt_um_rejunity_ay8913.noise_generator.lfsr\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_1649_ _0984_ _1180_ _1182_ tt_um_rejunity_ay8913.envelope_generator.period\[11\]
+ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1718_ tt_um_rejunity_ay8913.envelope_continue _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_56_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_ay8913_24 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_35 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_51_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1216__A3 _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2290__C _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2483_ _0097_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1503_ _1086_ tt_um_rejunity_ay8913.pwm_C.accumulator\[8\] _1084_ _1087_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_10_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2552_ _0166_ clknet_leaf_42_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2621_ _0235_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.latched_register\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1296_ _0929_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1365_ net6 _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1434_ _1011_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2331__A1 blink.LED vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2604_ _0218_ clknet_leaf_42_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1983_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\] _0515_ _0518_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2466_ _0080_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2535_ _0149_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1417_ tt_um_rejunity_ay8913.pwm_master.accumulator\[5\] _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2397_ _0011_ clknet_leaf_8_wb_clk_i blink.counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1279_ blink.counter\[12\] _0917_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1348_ _0965_ _0966_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2147__A4 _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2251_ _0754_ _0755_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2320_ tt_um_rejunity_ay8913.active _0806_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2182_ _0665_ _0691_ _0692_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1202_ tt_um_rejunity_ay8913.noise_disable_C _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1966_ _0497_ tt_um_rejunity_ay8913.noise_generator.period\[3\] tt_um_rejunity_ay8913.noise_generator.period\[4\]
+ _0505_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_34_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_0_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_0_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1897_ _0450_ _0451_ _0447_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2449_ _0063_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2518_ _0132_ clknet_leaf_32_wb_clk_i tt_um_rejunity_ay8913.tone_disable_B vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1820_ _0393_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_17_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1751_ _0322_ _0325_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1682_ _0275_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2234_ _0719_ tt_um_rejunity_ay8913.tone_A_generator.period\[1\] _0741_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2303_ tt_um_rejunity_ay8913.clk_counter\[3\] _0793_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2165_ _0678_ _0679_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2096_ _0613_ tt_um_rejunity_ay8913.tone_B_generator.period\[11\] tt_um_rejunity_ay8913.tone_B_generator.period\[10\]
+ _0615_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1949_ tt_um_rejunity_ay8913.noise_generator.lfsr\[16\] tt_um_rejunity_ay8913.noise_generator.lfsr\[15\]
+ tt_um_rejunity_ay8913.noise_generator.lfsr\[14\] tt_um_rejunity_ay8913.noise_generator.lfsr\[13\]
+ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_31_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1803_ net1 _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1665_ _0263_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1596_ _1149_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1734_ tt_um_rejunity_ay8913.envelope_generator.stop _0297_ _0300_ _0309_ _0310_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2217_ _0721_ tt_um_rejunity_ay8913.tone_A_generator.period\[5\] tt_um_rejunity_ay8913.tone_A_generator.period\[4\]
+ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_46_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2148_ _0610_ _0395_ _0630_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2079_ _0575_ _0601_ _0602_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1450_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\] _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1381_ _0994_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2002_ _0527_ _0534_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_33_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1648_ _1185_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1579_ _1133_ _1138_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1717_ _0296_ tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
+ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_56_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_ay8913_25 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_36 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1402__I _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1697__A1 _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2620_ _0234_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.latched_register\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1433_ tt_um_rejunity_ay8913.pwm_master.accumulator\[8\] _1033_ _1036_ _0047_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2482_ _0096_ clknet_leaf_37_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1502_ _1051_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2551_ _0165_ clknet_leaf_40_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1364_ _0981_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1295_ _0876_ _0927_ _0928_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1688__A1 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1679__A1 _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1603__A1 _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_24_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2331__A2 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1982_ _0511_ _0517_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2534_ _0148_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2603_ _0217_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2396_ _0010_ clknet_leaf_6_wb_clk_i blink.counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2465_ _0079_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1416_ _1020_ _1023_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1347_ tt_um_rejunity_ay8913.latched_register\[2\] _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1278_ _0910_ _0916_ _0917_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2086__A1 _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2250_ _0699_ _0395_ _0719_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1201_ tt_um_rejunity_ay8913.envelope_C _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2181_ _0622_ _0690_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1815__A1 _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1965_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[4\] _0505_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_43_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1896_ tt_um_rejunity_ay8913.noise_generator.lfsr\[2\] _0444_ _0451_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2517_ _0131_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_disable_A vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2448_ _0062_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2379_ _0843_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1806__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1750_ _0323_ tt_um_rejunity_ay8913.envelope_generator.period\[1\] tt_um_rejunity_ay8913.envelope_generator.period\[2\]
+ _0324_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_25_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1681_ _1100_ _0272_ _0273_ tt_um_rejunity_ay8913.tone_A_generator.period\[5\] _0275_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2164_ tt_um_rejunity_ay8913.tone_B_generator.counter\[5\] _0633_ tt_um_rejunity_ay8913.tone_B_generator.counter\[3\]
+ _0671_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_input9_I io_in_1[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2233_ tt_um_rejunity_ay8913.tone_A_generator.period\[5\] _0740_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2302_ _1082_ _0792_ _0793_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_45_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2095_ tt_um_rejunity_ay8913.tone_B_generator.counter\[10\] _0615_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1879_ tt_um_rejunity_ay8913.envelope_generator.invert_output _0435_ _0293_ _0437_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1948_ tt_um_rejunity_ay8913.noise_generator.lfsr\[12\] tt_um_rejunity_ay8913.noise_generator.lfsr\[11\]
+ tt_um_rejunity_ay8913.noise_generator.lfsr\[10\] tt_um_rejunity_ay8913.noise_generator.lfsr\[9\]
+ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_14_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1802_ _0322_ _0366_ _0373_ _0376_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1733_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\] tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\]
+ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\] _0295_ _0309_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_40_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1664_ _0976_ _0261_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1595_ tt_um_rejunity_ay8913.pwm_B.accumulator\[6\] _1146_ _1149_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_56_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2147_ tt_um_rejunity_ay8913.tone_B_generator.counter\[1\] tt_um_rejunity_ay8913.tone_B_generator.counter\[0\]
+ _0387_ _0388_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_2216_ _0722_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2078_ _0532_ _0600_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1380_ net14 _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2001_ _0529_ _0533_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1219__A2 _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1716_ tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal _0296_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1647_ _0982_ _1180_ _1182_ tt_um_rejunity_ay8913.envelope_generator.period\[10\]
+ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1578_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\] _1137_ _1138_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_16_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_ay8913_37 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_26 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_47_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2550_ _0164_ clknet_leaf_40_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1363_ _0980_ _0973_ _0978_ tt_um_rejunity_ay8913.noise_generator.period\[1\] _0981_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1432_ tt_um_rejunity_ay8913.pwm_master.accumulator\[8\] _1033_ _1008_ _1036_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2481_ _0095_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1501_ tt_um_rejunity_ay8913.pwm_C.accumulator\[8\] _1084_ _1085_ _0066_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1294_ _0876_ _0927_ _0889_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1413__I _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1981_ _0497_ _0515_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2533_ _0147_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1358__A1 _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2602_ _0216_ clknet_leaf_3_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2395_ _0009_ clknet_leaf_6_wb_clk_i blink.counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2464_ _0078_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1346_ tt_um_rejunity_ay8913.latched_register\[3\] _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1415_ _1021_ _1022_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1277_ blink.counter\[11\] _0877_ _0913_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2086__A2 _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_3__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1512__A1 _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2180_ _0622_ _0690_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1200_ tt_um_rejunity_ay8913.amplitude_C\[0\] _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1815__A2 _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1964_ _0497_ tt_um_rejunity_ay8913.noise_generator.period\[3\] tt_um_rejunity_ay8913.noise_generator.period\[2\]
+ _0502_ _0503_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1895_ tt_um_rejunity_ay8913.noise_generator.lfsr\[3\] _0440_ _0450_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2447_ _0061_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2516_ _0130_ clknet_leaf_40_wb_clk_i tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_11_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1329_ blink.counter\[27\] blink.counter\[26\] blink.counter\[25\] _0944_ _0953_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1503__A1 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2378_ _0260_ _0137_ _0842_ tt_um_rejunity_ay8913.envelope_generator.hold _0843_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1680_ _0274_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2301_ tt_um_rejunity_ay8913.clk_counter\[0\] _0789_ tt_um_rejunity_ay8913.clk_counter\[2\]
+ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_20_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2163_ _0633_ _0674_ tt_um_rejunity_ay8913.tone_B_generator.counter\[5\] _0678_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2232_ _0721_ tt_um_rejunity_ay8913.tone_A_generator.period\[5\] _0736_ _0738_ _0739_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_0_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2094_ _0613_ tt_um_rejunity_ay8913.tone_B_generator.period\[11\] _0614_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_0_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1972__A1 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1947_ tt_um_rejunity_ay8913.noise_generator.lfsr\[8\] tt_um_rejunity_ay8913.noise_generator.lfsr\[7\]
+ tt_um_rejunity_ay8913.noise_generator.lfsr\[6\] tt_um_rejunity_ay8913.noise_generator.lfsr\[5\]
+ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_1878_ tt_um_rejunity_ay8913.envelope_generator.invert_output _0435_ _0436_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_14_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1801_ _0374_ _0375_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1663_ _0261_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1732_ _0294_ _0308_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1594_ _1146_ _1148_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2146_ _0663_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2077_ _0532_ _0600_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2215_ tt_um_rejunity_ay8913.tone_A_generator.counter\[4\] _0722_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_18_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_18_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2361__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ tt_um_rejunity_ay8913.tone_C_generator.counter\[10\] _0530_ _0531_ _0532_
+ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1646_ _1184_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1715_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\] _0295_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1577_ _1132_ _1136_ _1137_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2129_ _0610_ tt_um_rejunity_ay8913.tone_B_generator.period\[0\] tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
+ _0630_ tt_um_rejunity_ay8913.tone_B_generator.counter\[2\] _0648_ _0649_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_51_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_ay8913_38 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_27 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_47_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1500_ tt_um_rejunity_ay8913.pwm_C.accumulator\[8\] _1084_ _1080_ _1085_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2480_ _0094_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1293_ _0923_ _0926_ _0927_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1362_ net5 _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1431_ _1033_ _1035_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1629_ _1171_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2325__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_33_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_33_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1980_ _0511_ _0515_ _0516_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2532_ _0146_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2601_ _0215_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2463_ _0077_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2394_ _0008_ clknet_leaf_6_wb_clk_i blink.counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1276_ _0877_ _0913_ blink.counter\[11\] _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1345_ net4 _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1414_ tt_um_rejunity_ay8913.pwm_master.accumulator\[4\] _1019_ _1022_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\] _0501_ _0503_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_11_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1894_ _0448_ _0449_ _0447_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2515_ _0129_ clknet_leaf_30_wb_clk_i net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2446_ _0060_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1259_ blink.counter\[6\] blink.counter\[5\] blink.counter\[4\] _0904_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1328_ blink.counter\[27\] _0951_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2377_ _1011_ _0292_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_46_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2231_ _0699_ tt_um_rejunity_ay8913.tone_A_generator.period\[0\] tt_um_rejunity_ay8913.tone_A_generator.period\[1\]
+ _0719_ tt_um_rejunity_ay8913.tone_A_generator.counter\[2\] _0737_ _0738_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_2300_ _0788_ _0789_ tt_um_rejunity_ay8913.clk_counter\[2\] _0792_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2162_ _0665_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2093_ tt_um_rejunity_ay8913.tone_B_generator.counter\[11\] _0613_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1239__I _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1972__A2 _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1946_ _0486_ _0487_ _1037_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1877_ _0298_ _0433_ _0434_ _0309_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2429_ _0043_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1800_ _0334_ _0316_ _0327_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_40_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1662_ _1088_ _1107_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1731_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\] _0307_ _0308_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2214_ tt_um_rejunity_ay8913.tone_A_generator.counter\[5\] _0721_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1593_ tt_um_rejunity_ay8913.pwm_B.accumulator\[5\] _1144_ _1147_ _1148_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2145_ _0611_ _0664_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2076_ tt_um_rejunity_ay8913.tone_C_generator.counter\[8\] _0594_ _0600_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1522__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1929_ _0452_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2189__A2 _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1872__A1 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1645_ _0980_ _1180_ _1182_ tt_um_rejunity_ay8913.envelope_generator.period\[9\]
+ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1576_ _1050_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\] tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
+ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_13_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1714_ _0293_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2128_ tt_um_rejunity_ay8913.tone_B_generator.period\[2\] _0648_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2059_ _0575_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xwrapped_ay8913_39 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_28 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1430_ tt_um_rejunity_ay8913.pwm_master.accumulator\[7\] _1028_ _1034_ _1035_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1292_ blink.counter\[16\] _0925_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1361_ _0979_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_3_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_3_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1559_ _1119_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1628_ _1021_ tt_um_rejunity_ay8913.pwm_A.accumulator\[7\] tt_um_rejunity_ay8913.pwm_A.accumulator\[8\]
+ _1166_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_52_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2600_ _0214_ clknet_leaf_3_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2393_ _0007_ clknet_leaf_6_wb_clk_i blink.counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2531_ _0145_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2462_ _0076_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1413_ _1002_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1275_ _0906_ _0915_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1344_ _0875_ _0963_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1993__B1 tt_um_rejunity_ay8913.tone_C_generator.period\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1350__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1962_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\] _0501_ _0502_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_28_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ tt_um_rejunity_ay8913.noise_generator.lfsr\[1\] _0444_ _0449_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2445_ _0059_ clknet_leaf_28_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2514_ _0128_ clknet_leaf_28_wb_clk_i net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2376_ _1177_ _0838_ _0839_ _0841_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1258_ blink.counter\[5\] blink.counter\[4\] _0898_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1327_ _0949_ _0950_ _0951_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_3_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2040__B _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2230_ tt_um_rejunity_ay8913.tone_A_generator.period\[2\] _0737_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1345__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2161_ _0676_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2092_ tt_um_rejunity_ay8913.tone_B_generator.counter\[8\] _0612_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1945_ tt_um_rejunity_ay8913.noise_generator.lfsr\[15\] _0480_ _0487_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1876_ _0298_ tt_um_rejunity_ay8913.envelope_attack _0311_ tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
+ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2359_ _1176_ _0830_ _0831_ tt_um_rejunity_ay8913.envelope_generator.period\[4\]
+ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2428_ _0042_ clknet_leaf_30_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1661_ net4 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1592_ _1007_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1730_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\] _0305_ _0307_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2144_ _0663_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2213_ _0699_ tt_um_rejunity_ay8913.tone_A_generator.period\[0\] tt_um_rejunity_ay8913.tone_A_generator.period\[1\]
+ _0719_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1803__I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I io_in_1[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2075_ _0599_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1859_ _0409_ _0421_ _0422_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1928_ _0473_ _0474_ _0467_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_27_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_27_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_41_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1713_ _0975_ tt_um_rejunity_ay8913.restart_envelope _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1644_ _1183_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1575_ _1131_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\] tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
+ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1560__A1 _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2127_ _0644_ _0645_ _0646_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2058_ _0586_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xwrapped_ay8913_29 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2040__A2 _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1606__A2 _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1360_ _0964_ _0973_ _0978_ tt_um_rejunity_ay8913.noise_generator.period\[0\] _0979_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1291_ blink.counter\[16\] _0925_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_52_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1558_ _1117_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1691__C _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1627_ _1012_ _1170_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1489_ _1076_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2308__B _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_42_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_42_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2530_ _0144_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2461_ _0075_ clknet_leaf_9_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2392_ _0006_ clknet_leaf_8_wb_clk_i blink.counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1343_ _0961_ _0962_ _0963_ _0893_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1412_ tt_um_rejunity_ay8913.pwm_master.accumulator\[4\] _1019_ _1020_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1818__A2 _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1274_ _0877_ _0913_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_3_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ _0498_ tt_um_rejunity_ay8913.noise_generator.period\[1\] _0500_ _0501_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_28_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1892_ tt_um_rejunity_ay8913.noise_generator.lfsr\[2\] _0440_ _0448_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2513_ _0127_ clknet_leaf_30_wb_clk_i net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1326_ blink.counter\[26\] _0946_ _0944_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2444_ _0058_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_3_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2375_ tt_um_rejunity_ay8913.envelope_B _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1257_ blink.counter\[6\] _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1541__I _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2321__B _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ _0664_ _0675_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2091_ _0610_ _0520_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1944_ tt_um_rejunity_ay8913.noise_generator.lfsr\[16\] _0452_ _0486_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1875_ tt_um_rejunity_ay8913.envelope_generator.hold tt_um_rejunity_ay8913.envelope_alternate
+ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2427_ _0041_ clknet_leaf_30_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1709__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2382__A1 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2358_ _0824_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2289_ _0785_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1309_ _0938_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_22_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1660_ _0259_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1591_ tt_um_rejunity_ay8913.pwm_B.accumulator\[5\] _1144_ _1146_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2143_ _0390_ _0662_ _1010_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2212_ tt_um_rejunity_ay8913.tone_A_generator.counter\[1\] _0719_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2074_ _0587_ _0598_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_36_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1858_ _0342_ _0345_ _0419_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_31_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1927_ tt_um_rejunity_ay8913.noise_generator.lfsr\[10\] _0469_ _0474_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1789_ _0353_ _0355_ _0358_ _0363_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__2355__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1643_ _0964_ _1180_ _1182_ tt_um_rejunity_ay8913.envelope_generator.period\[8\]
+ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1712_ _0292_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1574_ _1131_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\] _1135_ _0089_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2126_ tt_um_rejunity_ay8913.tone_B_generator.counter\[7\] _0641_ _0646_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2057_ _0574_ _0585_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_8_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2319__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1290_ _0923_ _0924_ _0925_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_53_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1626_ tt_um_rejunity_ay8913.pwm_A.accumulator\[8\] _1169_ _1170_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1557_ _1124_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1488_ tt_um_rejunity_ay8913.pwm_C.accumulator\[5\] _1074_ _1076_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_52_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2109_ _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2316__A4 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_11_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_11_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_37_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_2_0__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2460_ _0074_ clknet_leaf_9_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2391_ _0005_ clknet_leaf_7_wb_clk_i blink.counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1273_ _0910_ _0913_ _0914_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1342_ blink.counter\[30\] _0958_ blink.counter\[28\] _0953_ _0963_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1411_ _1018_ _1017_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_54_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2589_ _0203_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1609_ tt_um_rejunity_ay8913.pwm_A.accumulator\[3\] _1156_ _1158_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1203__B2 tt_um_rejunity_ay8913.noise_generator.lfsr\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1681__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1960_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\] _0499_ _0500_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1891_ _0441_ _0445_ _0447_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2512_ _0126_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2443_ _0057_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1256_ _0890_ _0901_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1325_ _0946_ _0945_ blink.counter\[26\] _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2374_ _0988_ _0838_ _0839_ _0840_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1672__A1 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1424__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1415__A1 _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ tt_um_rejunity_ay8913.tone_B_generator.counter\[0\] _0610_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__2143__A2 _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1874_ _0352_ _0432_ _0394_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1943_ _0484_ _0485_ _0478_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_24_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2426_ _0040_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1239_ _0889_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1645__A1 _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2357_ _0822_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1308_ blink.counter\[21\] _0936_ _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2288_ _0754_ _0783_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_22_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1590_ _1144_ _1145_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2142_ _0625_ _0640_ _0650_ _0658_ _0661_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_2073_ tt_um_rejunity_ay8913.tone_C_generator.counter\[8\] _0594_ _0598_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2211_ _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1627__A1 _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1788_ _0359_ _0360_ _0361_ _0362_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__1547__I _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1857_ _0345_ _0419_ _0342_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1926_ tt_um_rejunity_ay8913.noise_generator.lfsr\[11\] _0464_ _0473_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1866__A1 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2409_ _0023_ clknet_leaf_3_wb_clk_i blink.counter\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1457__I _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_36_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_33_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1642_ _1181_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1711_ _0965_ _1106_ _0991_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1573_ _1131_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\] _1048_ _1134_ _1135_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2125_ tt_um_rejunity_ay8913.tone_B_generator.counter\[6\] _0642_ _0645_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2056_ _0543_ _0584_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1909_ tt_um_rejunity_ay8913.noise_generator.lfsr\[5\] _0458_ _0461_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2319__A2 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1556_ _0984_ _1118_ _1120_ tt_um_rejunity_ay8913.tone_B_generator.period\[3\] _1124_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1625_ tt_um_rejunity_ay8913.pwm_A.accumulator\[7\] _1165_ _1169_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1487_ _1074_ _1075_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2108_ _0626_ tt_um_rejunity_ay8913.tone_B_generator.period\[3\] tt_um_rejunity_ay8913.tone_B_generator.period\[2\]
+ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2039_ _0535_ _0550_ _0560_ _0568_ _0571_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1470__I _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1410_ _1013_ _0871_ _0872_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2390_ _0004_ clknet_leaf_7_wb_clk_i blink.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1272_ blink.counter\[8\] _0908_ blink.counter\[9\] _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1341_ _0958_ _0955_ _0954_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1380__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2588_ _0202_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1539_ _1003_ tt_um_rejunity_ay8913.tone_B_generator.period\[9\] _1111_ _1113_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1608_ _1156_ _1157_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1690__A2 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2245__B _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1890_ _0446_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2511_ _0125_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2442_ _0056_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2373_ tt_um_rejunity_ay8913.amplitude_B\[0\] _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1255_ blink.counter\[5\] _0900_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1324_ _0888_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_49_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1360__A1 _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1942_ tt_um_rejunity_ay8913.noise_generator.lfsr\[14\] _0480_ _0485_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1873_ _0347_ _0429_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2356_ _0829_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2425_ _0039_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1238_ _0888_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1307_ blink.counter\[21\] _0936_ _0889_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2287_ tt_um_rejunity_ay8913.tone_A_generator.counter\[10\] _0711_ _0779_ _0784_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _0715_ tt_um_rejunity_ay8913.tone_A_generator.period\[3\] tt_um_rejunity_ay8913.tone_A_generator.period\[2\]
+ _0716_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2072_ _0597_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2141_ _0614_ _0660_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_36_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_6_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_6_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1925_ _0471_ _0472_ _0467_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1856_ _0404_ _0420_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1787_ _0340_ tt_um_rejunity_ay8913.envelope_generator.period\[8\] _0362_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2408_ _0022_ clknet_leaf_42_wb_clk_i blink.counter\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2339_ _0816_ tt_um_rejunity_ay8913.tone_A_generator.period\[9\] _0817_ _0819_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input13_I io_in_2[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2291__A2 _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1554__A1 _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1641_ _0976_ _1179_ _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1545__A1 _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1572_ _1051_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1710_ _0291_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2124_ tt_um_rejunity_ay8913.tone_B_generator.counter\[7\] _0641_ _0642_ _0643_ _0644_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input5_I io_in_1[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2055_ _0536_ _0537_ _0576_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1558__I _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1839_ _0404_ _0408_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1908_ tt_um_rejunity_ay8913.noise_generator.lfsr\[6\] _0453_ _0460_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1555_ _1123_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1624_ tt_um_rejunity_ay8913.pwm_A.accumulator\[7\] _1166_ _1168_ _0106_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2107_ tt_um_rejunity_ay8913.tone_B_generator.counter\[2\] _0627_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1486_ tt_um_rejunity_ay8913.pwm_C.accumulator\[4\] _1072_ _1034_ _1075_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_52_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2038_ _0524_ _0570_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1340_ blink.counter\[30\] _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1271_ _0912_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_20_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_20_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1661__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2587_ _0201_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1538_ _0989_ _1110_ _1112_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1469_ _1056_ _1064_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1607_ tt_um_rejunity_ay8913.pwm_A.accumulator\[2\] _0868_ _1147_ _1157_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1969__A1 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2510_ _0124_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1323_ _0948_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2441_ _0055_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2372_ _1052_ _0838_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1391__I _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1254_ blink.counter\[4\] _0898_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2639_ _0253_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.hold
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1872_ _0386_ _0430_ _0431_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1941_ tt_um_rejunity_ay8913.noise_generator.lfsr\[15\] _0475_ _0484_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1386__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2355_ _0270_ _0823_ _0825_ tt_um_rejunity_ay8913.envelope_generator.period\[3\]
+ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1306_ _0934_ _0935_ _0936_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2286_ _0704_ _0781_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2424_ _0038_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1237_ _0887_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2349__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2140_ _0619_ _0659_ _0616_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2071_ _0587_ _0596_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_36_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1855_ _0339_ _0419_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1924_ tt_um_rejunity_ay8913.noise_generator.lfsr\[9\] _0469_ _0472_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1786_ _0337_ tt_um_rejunity_ay8913.envelope_generator.period\[12\] _0361_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2269_ _0770_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2338_ _0989_ _0815_ _0818_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2407_ _0021_ clknet_leaf_42_wb_clk_i blink.counter\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ _1179_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1571_ _1131_ _1133_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2123_ tt_um_rejunity_ay8913.tone_B_generator.counter\[6\] _0643_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2054_ _0583_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1838_ _0406_ _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1907_ _0457_ _0459_ _0456_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1769_ tt_um_rejunity_ay8913.envelope_generator.period\[9\] _0344_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1463__A1 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1554_ _0982_ _1118_ _1120_ tt_um_rejunity_ay8913.tone_B_generator.period\[2\] _1123_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1394__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1623_ tt_um_rejunity_ay8913.pwm_A.accumulator\[7\] _1166_ _1080_ _1168_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1485_ tt_um_rejunity_ay8913.pwm_C.accumulator\[4\] _1072_ _1074_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
.ends

