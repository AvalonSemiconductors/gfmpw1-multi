magic
tech gf180mcuD
magscale 1 10
timestamp 1699037300
<< metal1 >>
rect 466 31502 478 31554
rect 530 31551 542 31554
rect 2258 31551 2270 31554
rect 530 31505 2270 31551
rect 530 31502 542 31505
rect 2258 31502 2270 31505
rect 2322 31502 2334 31554
rect 1344 31386 33760 31420
rect 1344 31334 9278 31386
rect 9330 31334 9382 31386
rect 9434 31334 9486 31386
rect 9538 31334 17342 31386
rect 17394 31334 17446 31386
rect 17498 31334 17550 31386
rect 17602 31334 25406 31386
rect 25458 31334 25510 31386
rect 25562 31334 25614 31386
rect 25666 31334 33470 31386
rect 33522 31334 33574 31386
rect 33626 31334 33678 31386
rect 33730 31334 33760 31386
rect 1344 31300 33760 31334
rect 1822 31218 1874 31230
rect 1822 31154 1874 31166
rect 2270 31218 2322 31230
rect 2270 31154 2322 31166
rect 2942 31218 2994 31230
rect 2942 31154 2994 31166
rect 3950 31218 4002 31230
rect 3950 31154 4002 31166
rect 4510 31218 4562 31230
rect 4510 31154 4562 31166
rect 4958 31218 5010 31230
rect 4958 31154 5010 31166
rect 5854 31218 5906 31230
rect 5854 31154 5906 31166
rect 18622 31218 18674 31230
rect 18622 31154 18674 31166
rect 21758 31218 21810 31230
rect 21758 31154 21810 31166
rect 24558 31218 24610 31230
rect 24558 31154 24610 31166
rect 26238 31218 26290 31230
rect 26238 31154 26290 31166
rect 3726 31106 3778 31118
rect 23662 31106 23714 31118
rect 7970 31054 7982 31106
rect 8034 31054 8046 31106
rect 16930 31054 16942 31106
rect 16994 31054 17006 31106
rect 24882 31054 24894 31106
rect 24946 31054 24958 31106
rect 29138 31054 29150 31106
rect 29202 31054 29214 31106
rect 3726 31042 3778 31054
rect 23662 31042 23714 31054
rect 17278 30994 17330 31006
rect 32286 30994 32338 31006
rect 6626 30942 6638 30994
rect 6690 30942 6702 30994
rect 9426 30942 9438 30994
rect 9490 30942 9502 30994
rect 13794 30942 13806 30994
rect 13858 30942 13870 30994
rect 17938 30942 17950 30994
rect 18002 30942 18014 30994
rect 20738 30942 20750 30994
rect 20802 30942 20814 30994
rect 23874 30942 23886 30994
rect 23938 30942 23950 30994
rect 25330 30942 25342 30994
rect 25394 30942 25406 30994
rect 28354 30942 28366 30994
rect 28418 30942 28430 30994
rect 17278 30930 17330 30942
rect 32286 30930 32338 30942
rect 32734 30994 32786 31006
rect 32734 30930 32786 30942
rect 12238 30882 12290 30894
rect 10098 30830 10110 30882
rect 10162 30830 10174 30882
rect 12238 30818 12290 30830
rect 13358 30882 13410 30894
rect 13358 30818 13410 30830
rect 16158 30882 16210 30894
rect 32174 30882 32226 30894
rect 31266 30830 31278 30882
rect 31330 30830 31342 30882
rect 16158 30818 16210 30830
rect 32174 30818 32226 30830
rect 13470 30770 13522 30782
rect 13470 30706 13522 30718
rect 32286 30770 32338 30782
rect 32286 30706 32338 30718
rect 32958 30770 33010 30782
rect 32958 30706 33010 30718
rect 1344 30602 33600 30636
rect 1344 30550 5246 30602
rect 5298 30550 5350 30602
rect 5402 30550 5454 30602
rect 5506 30550 13310 30602
rect 13362 30550 13414 30602
rect 13466 30550 13518 30602
rect 13570 30550 21374 30602
rect 21426 30550 21478 30602
rect 21530 30550 21582 30602
rect 21634 30550 29438 30602
rect 29490 30550 29542 30602
rect 29594 30550 29646 30602
rect 29698 30550 33600 30602
rect 1344 30516 33600 30550
rect 20638 30322 20690 30334
rect 5058 30270 5070 30322
rect 5122 30270 5134 30322
rect 8530 30270 8542 30322
rect 8594 30270 8606 30322
rect 18610 30270 18622 30322
rect 18674 30270 18686 30322
rect 27682 30270 27694 30322
rect 27746 30270 27758 30322
rect 32498 30270 32510 30322
rect 32562 30270 32574 30322
rect 20638 30258 20690 30270
rect 14814 30210 14866 30222
rect 2258 30158 2270 30210
rect 2322 30158 2334 30210
rect 5618 30158 5630 30210
rect 5682 30158 5694 30210
rect 9762 30158 9774 30210
rect 9826 30158 9838 30210
rect 13794 30158 13806 30210
rect 13858 30158 13870 30210
rect 14814 30146 14866 30158
rect 14926 30210 14978 30222
rect 19070 30210 19122 30222
rect 15698 30158 15710 30210
rect 15762 30158 15774 30210
rect 16482 30158 16494 30210
rect 16546 30158 16558 30210
rect 14926 30146 14978 30158
rect 19070 30146 19122 30158
rect 19630 30210 19682 30222
rect 29262 30210 29314 30222
rect 21298 30158 21310 30210
rect 21362 30158 21374 30210
rect 24882 30158 24894 30210
rect 24946 30158 24958 30210
rect 29586 30158 29598 30210
rect 29650 30158 29662 30210
rect 33058 30158 33070 30210
rect 33122 30158 33134 30210
rect 19630 30146 19682 30158
rect 29262 30146 29314 30158
rect 9326 30098 9378 30110
rect 15038 30098 15090 30110
rect 20414 30098 20466 30110
rect 2930 30046 2942 30098
rect 2994 30046 3006 30098
rect 6402 30046 6414 30098
rect 6466 30046 6478 30098
rect 10546 30046 10558 30098
rect 10610 30046 10622 30098
rect 20290 30046 20302 30098
rect 20354 30046 20366 30098
rect 22082 30046 22094 30098
rect 22146 30046 22158 30098
rect 25554 30046 25566 30098
rect 25618 30046 25630 30098
rect 30370 30046 30382 30098
rect 30434 30046 30446 30098
rect 32834 30046 32846 30098
rect 32898 30046 32910 30098
rect 9326 30034 9378 30046
rect 15038 30034 15090 30046
rect 20414 30034 20466 30046
rect 8878 29986 8930 29998
rect 8878 29922 8930 29934
rect 9438 29986 9490 29998
rect 14030 29986 14082 29998
rect 20526 29986 20578 29998
rect 12786 29934 12798 29986
rect 12850 29934 12862 29986
rect 14354 29934 14366 29986
rect 14418 29934 14430 29986
rect 9438 29922 9490 29934
rect 14030 29922 14082 29934
rect 20526 29922 20578 29934
rect 20750 29986 20802 29998
rect 28366 29986 28418 29998
rect 24322 29934 24334 29986
rect 24386 29934 24398 29986
rect 28018 29934 28030 29986
rect 28082 29934 28094 29986
rect 20750 29922 20802 29934
rect 28366 29922 28418 29934
rect 1344 29818 33760 29852
rect 1344 29766 9278 29818
rect 9330 29766 9382 29818
rect 9434 29766 9486 29818
rect 9538 29766 17342 29818
rect 17394 29766 17446 29818
rect 17498 29766 17550 29818
rect 17602 29766 25406 29818
rect 25458 29766 25510 29818
rect 25562 29766 25614 29818
rect 25666 29766 33470 29818
rect 33522 29766 33574 29818
rect 33626 29766 33678 29818
rect 33730 29766 33760 29818
rect 1344 29732 33760 29766
rect 3950 29650 4002 29662
rect 3950 29586 4002 29598
rect 5070 29650 5122 29662
rect 5070 29586 5122 29598
rect 5518 29650 5570 29662
rect 5518 29586 5570 29598
rect 7198 29650 7250 29662
rect 7198 29586 7250 29598
rect 9102 29650 9154 29662
rect 9102 29586 9154 29598
rect 10110 29650 10162 29662
rect 10110 29586 10162 29598
rect 11678 29650 11730 29662
rect 11678 29586 11730 29598
rect 18398 29650 18450 29662
rect 18398 29586 18450 29598
rect 22318 29650 22370 29662
rect 22318 29586 22370 29598
rect 22542 29650 22594 29662
rect 22542 29586 22594 29598
rect 10222 29538 10274 29550
rect 15934 29538 15986 29550
rect 6066 29486 6078 29538
rect 6130 29486 6142 29538
rect 7410 29486 7422 29538
rect 7474 29486 7486 29538
rect 8194 29486 8206 29538
rect 8258 29486 8270 29538
rect 8530 29486 8542 29538
rect 8594 29486 8606 29538
rect 11330 29486 11342 29538
rect 11394 29486 11406 29538
rect 12786 29486 12798 29538
rect 12850 29486 12862 29538
rect 10222 29474 10274 29486
rect 15934 29474 15986 29486
rect 22990 29538 23042 29550
rect 22990 29474 23042 29486
rect 23102 29538 23154 29550
rect 30594 29486 30606 29538
rect 30658 29486 30670 29538
rect 23102 29474 23154 29486
rect 7758 29426 7810 29438
rect 15710 29426 15762 29438
rect 5842 29374 5854 29426
rect 5906 29374 5918 29426
rect 8642 29374 8654 29426
rect 8706 29374 8718 29426
rect 12114 29374 12126 29426
rect 12178 29374 12190 29426
rect 7758 29362 7810 29374
rect 15710 29362 15762 29374
rect 15822 29426 15874 29438
rect 17726 29426 17778 29438
rect 16146 29374 16158 29426
rect 16210 29374 16222 29426
rect 15822 29362 15874 29374
rect 17726 29362 17778 29374
rect 18174 29426 18226 29438
rect 22206 29426 22258 29438
rect 18834 29374 18846 29426
rect 18898 29374 18910 29426
rect 18174 29362 18226 29374
rect 22206 29362 22258 29374
rect 22766 29426 22818 29438
rect 22766 29362 22818 29374
rect 22878 29426 22930 29438
rect 24110 29426 24162 29438
rect 25454 29426 25506 29438
rect 23426 29374 23438 29426
rect 23490 29374 23502 29426
rect 24434 29374 24446 29426
rect 24498 29374 24510 29426
rect 22878 29362 22930 29374
rect 24110 29362 24162 29374
rect 25454 29362 25506 29374
rect 26126 29426 26178 29438
rect 26562 29374 26574 29426
rect 26626 29374 26638 29426
rect 31938 29374 31950 29426
rect 32002 29374 32014 29426
rect 26126 29362 26178 29374
rect 4062 29314 4114 29326
rect 4062 29250 4114 29262
rect 4510 29314 4562 29326
rect 4510 29250 4562 29262
rect 6750 29314 6802 29326
rect 6750 29250 6802 29262
rect 8094 29314 8146 29326
rect 8094 29250 8146 29262
rect 9662 29314 9714 29326
rect 9662 29250 9714 29262
rect 10894 29314 10946 29326
rect 17390 29314 17442 29326
rect 14914 29262 14926 29314
rect 14978 29262 14990 29314
rect 10894 29250 10946 29262
rect 17390 29250 17442 29262
rect 18286 29314 18338 29326
rect 23886 29314 23938 29326
rect 33182 29314 33234 29326
rect 19506 29262 19518 29314
rect 19570 29262 19582 29314
rect 21746 29262 21758 29314
rect 21810 29262 21822 29314
rect 27346 29262 27358 29314
rect 27410 29262 27422 29314
rect 29474 29262 29486 29314
rect 29538 29262 29550 29314
rect 18286 29250 18338 29262
rect 23886 29250 23938 29262
rect 33182 29250 33234 29262
rect 9998 29202 10050 29214
rect 9998 29138 10050 29150
rect 11006 29202 11058 29214
rect 11006 29138 11058 29150
rect 16606 29202 16658 29214
rect 16606 29138 16658 29150
rect 17502 29202 17554 29214
rect 17502 29138 17554 29150
rect 25678 29202 25730 29214
rect 25678 29138 25730 29150
rect 26126 29202 26178 29214
rect 26126 29138 26178 29150
rect 26238 29202 26290 29214
rect 26238 29138 26290 29150
rect 1344 29034 33600 29068
rect 1344 28982 5246 29034
rect 5298 28982 5350 29034
rect 5402 28982 5454 29034
rect 5506 28982 13310 29034
rect 13362 28982 13414 29034
rect 13466 28982 13518 29034
rect 13570 28982 21374 29034
rect 21426 28982 21478 29034
rect 21530 28982 21582 29034
rect 21634 28982 29438 29034
rect 29490 28982 29542 29034
rect 29594 28982 29646 29034
rect 29698 28982 33600 29034
rect 1344 28948 33600 28982
rect 9662 28866 9714 28878
rect 8418 28814 8430 28866
rect 8482 28863 8494 28866
rect 9314 28863 9326 28866
rect 8482 28817 9326 28863
rect 8482 28814 8494 28817
rect 9314 28814 9326 28817
rect 9378 28814 9390 28866
rect 9662 28802 9714 28814
rect 11342 28866 11394 28878
rect 11342 28802 11394 28814
rect 18734 28866 18786 28878
rect 18734 28802 18786 28814
rect 26910 28866 26962 28878
rect 26910 28802 26962 28814
rect 7646 28754 7698 28766
rect 4610 28702 4622 28754
rect 4674 28702 4686 28754
rect 6066 28702 6078 28754
rect 6130 28702 6142 28754
rect 7646 28690 7698 28702
rect 8430 28754 8482 28766
rect 8430 28690 8482 28702
rect 9326 28754 9378 28766
rect 9326 28690 9378 28702
rect 13470 28754 13522 28766
rect 18274 28702 18286 28754
rect 18338 28702 18350 28754
rect 21858 28702 21870 28754
rect 21922 28702 21934 28754
rect 23426 28702 23438 28754
rect 23490 28702 23502 28754
rect 25554 28702 25566 28754
rect 25618 28702 25630 28754
rect 29922 28702 29934 28754
rect 29986 28702 29998 28754
rect 31042 28702 31054 28754
rect 31106 28702 31118 28754
rect 33170 28702 33182 28754
rect 33234 28702 33246 28754
rect 13470 28690 13522 28702
rect 5182 28642 5234 28654
rect 14478 28642 14530 28654
rect 1698 28590 1710 28642
rect 1762 28590 1774 28642
rect 6402 28590 6414 28642
rect 6466 28590 6478 28642
rect 7858 28590 7870 28642
rect 7922 28590 7934 28642
rect 10322 28590 10334 28642
rect 10386 28590 10398 28642
rect 14130 28590 14142 28642
rect 14194 28590 14206 28642
rect 5182 28578 5234 28590
rect 14478 28578 14530 28590
rect 15038 28642 15090 28654
rect 19294 28642 19346 28654
rect 15474 28590 15486 28642
rect 15538 28590 15550 28642
rect 15038 28578 15090 28590
rect 19294 28578 19346 28590
rect 19966 28642 20018 28654
rect 19966 28578 20018 28590
rect 20302 28642 20354 28654
rect 22194 28590 22206 28642
rect 22258 28590 22270 28642
rect 22642 28590 22654 28642
rect 22706 28590 22718 28642
rect 25890 28590 25902 28642
rect 25954 28590 25966 28642
rect 30258 28590 30270 28642
rect 30322 28590 30334 28642
rect 20302 28578 20354 28590
rect 6638 28530 6690 28542
rect 2482 28478 2494 28530
rect 2546 28478 2558 28530
rect 6290 28478 6302 28530
rect 6354 28478 6366 28530
rect 6638 28466 6690 28478
rect 7534 28530 7586 28542
rect 7534 28466 7586 28478
rect 9998 28530 10050 28542
rect 9998 28466 10050 28478
rect 13694 28530 13746 28542
rect 13694 28466 13746 28478
rect 13806 28530 13858 28542
rect 18734 28530 18786 28542
rect 14690 28478 14702 28530
rect 14754 28478 14766 28530
rect 16146 28478 16158 28530
rect 16210 28478 16222 28530
rect 13806 28466 13858 28478
rect 18734 28466 18786 28478
rect 18846 28530 18898 28542
rect 18846 28466 18898 28478
rect 20638 28530 20690 28542
rect 20638 28466 20690 28478
rect 21534 28530 21586 28542
rect 21534 28466 21586 28478
rect 21870 28530 21922 28542
rect 21870 28466 21922 28478
rect 29374 28530 29426 28542
rect 29374 28466 29426 28478
rect 29486 28530 29538 28542
rect 29586 28478 29598 28530
rect 29650 28478 29662 28530
rect 29486 28466 29538 28478
rect 5742 28418 5794 28430
rect 5742 28354 5794 28366
rect 6862 28418 6914 28430
rect 6862 28354 6914 28366
rect 8990 28418 9042 28430
rect 8990 28354 9042 28366
rect 9774 28418 9826 28430
rect 9774 28354 9826 28366
rect 19182 28418 19234 28430
rect 19182 28354 19234 28366
rect 19406 28418 19458 28430
rect 19406 28354 19458 28366
rect 19630 28418 19682 28430
rect 19630 28354 19682 28366
rect 20190 28418 20242 28430
rect 20190 28354 20242 28366
rect 21758 28418 21810 28430
rect 21758 28354 21810 28366
rect 29150 28418 29202 28430
rect 29150 28354 29202 28366
rect 1344 28250 33760 28284
rect 1344 28198 9278 28250
rect 9330 28198 9382 28250
rect 9434 28198 9486 28250
rect 9538 28198 17342 28250
rect 17394 28198 17446 28250
rect 17498 28198 17550 28250
rect 17602 28198 25406 28250
rect 25458 28198 25510 28250
rect 25562 28198 25614 28250
rect 25666 28198 33470 28250
rect 33522 28198 33574 28250
rect 33626 28198 33678 28250
rect 33730 28198 33760 28250
rect 1344 28164 33760 28198
rect 5070 28082 5122 28094
rect 5070 28018 5122 28030
rect 5518 28082 5570 28094
rect 5518 28018 5570 28030
rect 8094 28082 8146 28094
rect 8094 28018 8146 28030
rect 12238 28082 12290 28094
rect 12238 28018 12290 28030
rect 15150 28082 15202 28094
rect 15150 28018 15202 28030
rect 18510 28082 18562 28094
rect 18510 28018 18562 28030
rect 20526 28082 20578 28094
rect 20526 28018 20578 28030
rect 24334 28082 24386 28094
rect 24334 28018 24386 28030
rect 24558 28082 24610 28094
rect 26126 28082 26178 28094
rect 25778 28030 25790 28082
rect 25842 28030 25854 28082
rect 24558 28018 24610 28030
rect 26126 28018 26178 28030
rect 26238 28082 26290 28094
rect 26238 28018 26290 28030
rect 26350 28082 26402 28094
rect 26350 28018 26402 28030
rect 7758 27970 7810 27982
rect 7758 27906 7810 27918
rect 9662 27970 9714 27982
rect 9662 27906 9714 27918
rect 9886 27970 9938 27982
rect 9886 27906 9938 27918
rect 10782 27970 10834 27982
rect 10782 27906 10834 27918
rect 24670 27970 24722 27982
rect 24670 27906 24722 27918
rect 26462 27970 26514 27982
rect 30258 27918 30270 27970
rect 30322 27918 30334 27970
rect 26462 27906 26514 27918
rect 7198 27858 7250 27870
rect 1698 27806 1710 27858
rect 1762 27806 1774 27858
rect 6290 27806 6302 27858
rect 6354 27806 6366 27858
rect 7198 27794 7250 27806
rect 9774 27858 9826 27870
rect 9774 27794 9826 27806
rect 10670 27858 10722 27870
rect 20414 27858 20466 27870
rect 25454 27858 25506 27870
rect 11218 27806 11230 27858
rect 11282 27806 11294 27858
rect 14130 27806 14142 27858
rect 14194 27806 14206 27858
rect 17714 27806 17726 27858
rect 17778 27806 17790 27858
rect 20962 27806 20974 27858
rect 21026 27806 21038 27858
rect 26898 27806 26910 27858
rect 26962 27806 26974 27858
rect 27234 27806 27246 27858
rect 27298 27806 27310 27858
rect 10670 27794 10722 27806
rect 20414 27794 20466 27806
rect 25454 27794 25506 27806
rect 8542 27746 8594 27758
rect 2482 27694 2494 27746
rect 2546 27694 2558 27746
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 6738 27694 6750 27746
rect 6802 27694 6814 27746
rect 8542 27682 8594 27694
rect 9102 27746 9154 27758
rect 25230 27746 25282 27758
rect 21746 27694 21758 27746
rect 21810 27694 21822 27746
rect 23986 27694 23998 27746
rect 24050 27694 24062 27746
rect 9102 27682 9154 27694
rect 25230 27682 25282 27694
rect 33182 27746 33234 27758
rect 33182 27682 33234 27694
rect 10782 27634 10834 27646
rect 7298 27582 7310 27634
rect 7362 27631 7374 27634
rect 7522 27631 7534 27634
rect 7362 27585 7534 27631
rect 7362 27582 7374 27585
rect 7522 27582 7534 27585
rect 7586 27582 7598 27634
rect 10322 27582 10334 27634
rect 10386 27582 10398 27634
rect 10782 27570 10834 27582
rect 20526 27634 20578 27646
rect 20526 27570 20578 27582
rect 1344 27466 33600 27500
rect 1344 27414 5246 27466
rect 5298 27414 5350 27466
rect 5402 27414 5454 27466
rect 5506 27414 13310 27466
rect 13362 27414 13414 27466
rect 13466 27414 13518 27466
rect 13570 27414 21374 27466
rect 21426 27414 21478 27466
rect 21530 27414 21582 27466
rect 21634 27414 29438 27466
rect 29490 27414 29542 27466
rect 29594 27414 29646 27466
rect 29698 27414 33600 27466
rect 1344 27380 33600 27414
rect 2830 27298 2882 27310
rect 2830 27234 2882 27246
rect 3278 27298 3330 27310
rect 3278 27234 3330 27246
rect 12574 27298 12626 27310
rect 14142 27298 14194 27310
rect 28478 27298 28530 27310
rect 12898 27246 12910 27298
rect 12962 27246 12974 27298
rect 18722 27246 18734 27298
rect 18786 27246 18798 27298
rect 12574 27234 12626 27246
rect 14142 27234 14194 27246
rect 28478 27234 28530 27246
rect 2942 27186 2994 27198
rect 2942 27122 2994 27134
rect 6302 27186 6354 27198
rect 7982 27186 8034 27198
rect 6738 27134 6750 27186
rect 6802 27134 6814 27186
rect 6302 27122 6354 27134
rect 7982 27122 8034 27134
rect 9214 27186 9266 27198
rect 12350 27186 12402 27198
rect 28590 27186 28642 27198
rect 9986 27134 9998 27186
rect 10050 27134 10062 27186
rect 10658 27134 10670 27186
rect 10722 27134 10734 27186
rect 16818 27134 16830 27186
rect 16882 27134 16894 27186
rect 22306 27134 22318 27186
rect 22370 27134 22382 27186
rect 26002 27134 26014 27186
rect 26066 27134 26078 27186
rect 28130 27134 28142 27186
rect 28194 27134 28206 27186
rect 31042 27134 31054 27186
rect 31106 27134 31118 27186
rect 33170 27134 33182 27186
rect 33234 27134 33246 27186
rect 9214 27122 9266 27134
rect 12350 27122 12402 27134
rect 28590 27122 28642 27134
rect 4846 27074 4898 27086
rect 4846 27010 4898 27022
rect 7534 27074 7586 27086
rect 10782 27074 10834 27086
rect 8530 27022 8542 27074
rect 8594 27022 8606 27074
rect 9538 27022 9550 27074
rect 9602 27022 9614 27074
rect 10210 27022 10222 27074
rect 10274 27022 10286 27074
rect 7534 27010 7586 27022
rect 10782 27010 10834 27022
rect 11790 27074 11842 27086
rect 14590 27074 14642 27086
rect 19294 27074 19346 27086
rect 14466 27022 14478 27074
rect 14530 27022 14542 27074
rect 15698 27022 15710 27074
rect 15762 27022 15774 27074
rect 18722 27022 18734 27074
rect 18786 27022 18798 27074
rect 19954 27022 19966 27074
rect 20018 27022 20030 27074
rect 20514 27022 20526 27074
rect 20578 27022 20590 27074
rect 24098 27022 24110 27074
rect 24162 27022 24174 27074
rect 25330 27022 25342 27074
rect 25394 27022 25406 27074
rect 29586 27022 29598 27074
rect 29650 27022 29662 27074
rect 29922 27022 29934 27074
rect 29986 27022 29998 27074
rect 30258 27022 30270 27074
rect 30322 27022 30334 27074
rect 11790 27010 11842 27022
rect 14590 27010 14642 27022
rect 19294 27010 19346 27022
rect 3390 26962 3442 26974
rect 3390 26898 3442 26910
rect 5182 26962 5234 26974
rect 6078 26962 6130 26974
rect 5954 26910 5966 26962
rect 6018 26910 6030 26962
rect 5182 26898 5234 26910
rect 6078 26898 6130 26910
rect 6190 26962 6242 26974
rect 7198 26962 7250 26974
rect 6962 26910 6974 26962
rect 7026 26910 7038 26962
rect 6190 26898 6242 26910
rect 7198 26898 7250 26910
rect 8094 26962 8146 26974
rect 8094 26898 8146 26910
rect 8206 26962 8258 26974
rect 8206 26898 8258 26910
rect 10670 26962 10722 26974
rect 10670 26898 10722 26910
rect 11006 26962 11058 26974
rect 11006 26898 11058 26910
rect 11230 26962 11282 26974
rect 11230 26898 11282 26910
rect 11902 26962 11954 26974
rect 14814 26962 14866 26974
rect 13458 26910 13470 26962
rect 13522 26910 13534 26962
rect 11902 26898 11954 26910
rect 14814 26898 14866 26910
rect 18174 26962 18226 26974
rect 21310 26962 21362 26974
rect 18386 26910 18398 26962
rect 18450 26910 18462 26962
rect 20626 26910 20638 26962
rect 20690 26910 20702 26962
rect 18174 26898 18226 26910
rect 21310 26898 21362 26910
rect 29262 26962 29314 26974
rect 29262 26898 29314 26910
rect 29374 26962 29426 26974
rect 29374 26898 29426 26910
rect 4958 26850 5010 26862
rect 4958 26786 5010 26798
rect 6414 26850 6466 26862
rect 6414 26786 6466 26798
rect 7310 26850 7362 26862
rect 7310 26786 7362 26798
rect 7870 26850 7922 26862
rect 7870 26786 7922 26798
rect 9774 26850 9826 26862
rect 9774 26786 9826 26798
rect 9998 26850 10050 26862
rect 9998 26786 10050 26798
rect 12126 26850 12178 26862
rect 12126 26786 12178 26798
rect 13806 26850 13858 26862
rect 13806 26786 13858 26798
rect 14702 26850 14754 26862
rect 14702 26786 14754 26798
rect 18958 26850 19010 26862
rect 18958 26786 19010 26798
rect 19406 26850 19458 26862
rect 29150 26850 29202 26862
rect 21634 26798 21646 26850
rect 21698 26798 21710 26850
rect 19406 26786 19458 26798
rect 29150 26786 29202 26798
rect 1344 26682 33760 26716
rect 1344 26630 9278 26682
rect 9330 26630 9382 26682
rect 9434 26630 9486 26682
rect 9538 26630 17342 26682
rect 17394 26630 17446 26682
rect 17498 26630 17550 26682
rect 17602 26630 25406 26682
rect 25458 26630 25510 26682
rect 25562 26630 25614 26682
rect 25666 26630 33470 26682
rect 33522 26630 33574 26682
rect 33626 26630 33678 26682
rect 33730 26630 33760 26682
rect 1344 26596 33760 26630
rect 7758 26514 7810 26526
rect 7758 26450 7810 26462
rect 12462 26514 12514 26526
rect 12462 26450 12514 26462
rect 12574 26514 12626 26526
rect 12574 26450 12626 26462
rect 14030 26514 14082 26526
rect 17726 26514 17778 26526
rect 16258 26462 16270 26514
rect 16322 26462 16334 26514
rect 14030 26450 14082 26462
rect 17726 26450 17778 26462
rect 18398 26514 18450 26526
rect 18398 26450 18450 26462
rect 18622 26514 18674 26526
rect 18622 26450 18674 26462
rect 19966 26514 20018 26526
rect 19966 26450 20018 26462
rect 6526 26402 6578 26414
rect 8542 26402 8594 26414
rect 11118 26402 11170 26414
rect 7410 26350 7422 26402
rect 7474 26350 7486 26402
rect 9762 26350 9774 26402
rect 9826 26350 9838 26402
rect 6526 26338 6578 26350
rect 8542 26338 8594 26350
rect 11118 26338 11170 26350
rect 15934 26402 15986 26414
rect 29598 26402 29650 26414
rect 26898 26350 26910 26402
rect 26962 26350 26974 26402
rect 30706 26350 30718 26402
rect 30770 26350 30782 26402
rect 15934 26338 15986 26350
rect 29598 26338 29650 26350
rect 6302 26290 6354 26302
rect 8430 26290 8482 26302
rect 5058 26238 5070 26290
rect 5122 26238 5134 26290
rect 6738 26238 6750 26290
rect 6802 26238 6814 26290
rect 6962 26238 6974 26290
rect 7026 26238 7038 26290
rect 6302 26226 6354 26238
rect 8430 26226 8482 26238
rect 8990 26290 9042 26302
rect 10558 26290 10610 26302
rect 12686 26290 12738 26302
rect 16830 26290 16882 26302
rect 19182 26290 19234 26302
rect 9986 26238 9998 26290
rect 10050 26238 10062 26290
rect 11890 26238 11902 26290
rect 11954 26238 11966 26290
rect 12226 26238 12238 26290
rect 12290 26238 12302 26290
rect 13010 26238 13022 26290
rect 13074 26238 13086 26290
rect 16146 26238 16158 26290
rect 16210 26238 16222 26290
rect 18162 26238 18174 26290
rect 18226 26238 18238 26290
rect 18834 26238 18846 26290
rect 18898 26238 18910 26290
rect 8990 26226 9042 26238
rect 10558 26226 10610 26238
rect 12686 26226 12738 26238
rect 16830 26226 16882 26238
rect 19182 26226 19234 26238
rect 19518 26290 19570 26302
rect 20190 26290 20242 26302
rect 19730 26238 19742 26290
rect 19794 26238 19806 26290
rect 19518 26226 19570 26238
rect 20190 26226 20242 26238
rect 20638 26290 20690 26302
rect 20638 26226 20690 26238
rect 20750 26290 20802 26302
rect 28814 26290 28866 26302
rect 21634 26238 21646 26290
rect 21698 26238 21710 26290
rect 25330 26238 25342 26290
rect 25394 26238 25406 26290
rect 20750 26226 20802 26238
rect 28814 26226 28866 26238
rect 29038 26290 29090 26302
rect 29038 26226 29090 26238
rect 29486 26290 29538 26302
rect 32162 26238 32174 26290
rect 32226 26238 32238 26290
rect 29486 26226 29538 26238
rect 5518 26178 5570 26190
rect 8766 26178 8818 26190
rect 5170 26126 5182 26178
rect 5234 26126 5246 26178
rect 7074 26126 7086 26178
rect 7138 26126 7150 26178
rect 5518 26114 5570 26126
rect 8766 26114 8818 26126
rect 16606 26178 16658 26190
rect 19630 26178 19682 26190
rect 17826 26126 17838 26178
rect 17890 26126 17902 26178
rect 18722 26126 18734 26178
rect 18786 26126 18798 26178
rect 16606 26114 16658 26126
rect 19630 26114 19682 26126
rect 20414 26178 20466 26190
rect 24446 26178 24498 26190
rect 22306 26126 22318 26178
rect 22370 26126 22382 26178
rect 20414 26114 20466 26126
rect 24446 26114 24498 26126
rect 28478 26178 28530 26190
rect 28478 26114 28530 26126
rect 33182 26178 33234 26190
rect 33182 26114 33234 26126
rect 10782 26066 10834 26078
rect 10782 26002 10834 26014
rect 11230 26066 11282 26078
rect 11230 26002 11282 26014
rect 11342 26066 11394 26078
rect 11342 26002 11394 26014
rect 16382 26066 16434 26078
rect 16382 26002 16434 26014
rect 17502 26066 17554 26078
rect 17502 26002 17554 26014
rect 29486 26066 29538 26078
rect 29486 26002 29538 26014
rect 1344 25898 33600 25932
rect 1344 25846 5246 25898
rect 5298 25846 5350 25898
rect 5402 25846 5454 25898
rect 5506 25846 13310 25898
rect 13362 25846 13414 25898
rect 13466 25846 13518 25898
rect 13570 25846 21374 25898
rect 21426 25846 21478 25898
rect 21530 25846 21582 25898
rect 21634 25846 29438 25898
rect 29490 25846 29542 25898
rect 29594 25846 29646 25898
rect 29698 25846 33600 25898
rect 1344 25812 33600 25846
rect 9550 25730 9602 25742
rect 9550 25666 9602 25678
rect 9886 25730 9938 25742
rect 9886 25666 9938 25678
rect 16830 25730 16882 25742
rect 16830 25666 16882 25678
rect 27806 25730 27858 25742
rect 27806 25666 27858 25678
rect 4174 25618 4226 25630
rect 4174 25554 4226 25566
rect 4622 25618 4674 25630
rect 4622 25554 4674 25566
rect 5742 25618 5794 25630
rect 9214 25618 9266 25630
rect 16942 25618 16994 25630
rect 6514 25566 6526 25618
rect 6578 25566 6590 25618
rect 12114 25566 12126 25618
rect 12178 25566 12190 25618
rect 15474 25566 15486 25618
rect 15538 25566 15550 25618
rect 5742 25554 5794 25566
rect 9214 25554 9266 25566
rect 16942 25554 16994 25566
rect 17726 25618 17778 25630
rect 17726 25554 17778 25566
rect 18958 25618 19010 25630
rect 28254 25618 28306 25630
rect 27458 25566 27470 25618
rect 27522 25566 27534 25618
rect 31042 25566 31054 25618
rect 31106 25566 31118 25618
rect 33170 25566 33182 25618
rect 33234 25566 33246 25618
rect 18958 25554 19010 25566
rect 28254 25554 28306 25566
rect 4734 25506 4786 25518
rect 4734 25442 4786 25454
rect 5182 25506 5234 25518
rect 7758 25506 7810 25518
rect 10558 25506 10610 25518
rect 5182 25442 5234 25454
rect 6526 25450 6578 25462
rect 7410 25454 7422 25506
rect 7474 25454 7486 25506
rect 10210 25454 10222 25506
rect 10274 25454 10286 25506
rect 7758 25442 7810 25454
rect 10558 25442 10610 25454
rect 11006 25506 11058 25518
rect 11006 25442 11058 25454
rect 11342 25506 11394 25518
rect 13918 25506 13970 25518
rect 11342 25442 11394 25454
rect 12686 25450 12738 25462
rect 6290 25342 6302 25394
rect 6354 25342 6366 25394
rect 6526 25386 6578 25398
rect 6638 25394 6690 25406
rect 6638 25330 6690 25342
rect 7198 25394 7250 25406
rect 7198 25330 7250 25342
rect 9662 25394 9714 25406
rect 11678 25394 11730 25406
rect 12574 25394 12626 25406
rect 9662 25330 9714 25342
rect 11454 25338 11506 25350
rect 3950 25282 4002 25294
rect 3950 25218 4002 25230
rect 4062 25282 4114 25294
rect 4062 25218 4114 25230
rect 4510 25282 4562 25294
rect 4510 25218 4562 25230
rect 6862 25282 6914 25294
rect 6862 25218 6914 25230
rect 7086 25282 7138 25294
rect 7086 25218 7138 25230
rect 9550 25282 9602 25294
rect 9550 25218 9602 25230
rect 9998 25282 10050 25294
rect 9998 25218 10050 25230
rect 10670 25282 10722 25294
rect 10670 25218 10722 25230
rect 10894 25282 10946 25294
rect 12338 25342 12350 25394
rect 12402 25342 12414 25394
rect 13918 25442 13970 25454
rect 14254 25506 14306 25518
rect 14254 25442 14306 25454
rect 14478 25506 14530 25518
rect 14478 25442 14530 25454
rect 15374 25506 15426 25518
rect 15374 25442 15426 25454
rect 15822 25506 15874 25518
rect 15822 25442 15874 25454
rect 16270 25506 16322 25518
rect 18510 25506 18562 25518
rect 17490 25454 17502 25506
rect 17554 25454 17566 25506
rect 17826 25454 17838 25506
rect 17890 25454 17902 25506
rect 16270 25442 16322 25454
rect 18510 25442 18562 25454
rect 18846 25506 18898 25518
rect 18846 25442 18898 25454
rect 19182 25506 19234 25518
rect 27022 25506 27074 25518
rect 26562 25454 26574 25506
rect 26626 25454 26638 25506
rect 19182 25442 19234 25454
rect 27022 25442 27074 25454
rect 27246 25506 27298 25518
rect 29374 25506 29426 25518
rect 28130 25454 28142 25506
rect 28194 25454 28206 25506
rect 29698 25454 29710 25506
rect 29762 25454 29774 25506
rect 30258 25454 30270 25506
rect 30322 25454 30334 25506
rect 27246 25442 27298 25454
rect 29374 25442 29426 25454
rect 12686 25386 12738 25398
rect 12910 25394 12962 25406
rect 11678 25330 11730 25342
rect 12574 25330 12626 25342
rect 12910 25330 12962 25342
rect 13694 25394 13746 25406
rect 13694 25330 13746 25342
rect 14926 25394 14978 25406
rect 14926 25330 14978 25342
rect 15150 25394 15202 25406
rect 15150 25330 15202 25342
rect 16494 25394 16546 25406
rect 16494 25330 16546 25342
rect 17278 25394 17330 25406
rect 17278 25330 17330 25342
rect 20526 25394 20578 25406
rect 20526 25330 20578 25342
rect 20638 25394 20690 25406
rect 27582 25394 27634 25406
rect 21970 25342 21982 25394
rect 22034 25342 22046 25394
rect 20638 25330 20690 25342
rect 27582 25330 27634 25342
rect 28590 25394 28642 25406
rect 28590 25330 28642 25342
rect 11454 25274 11506 25286
rect 14590 25282 14642 25294
rect 10894 25218 10946 25230
rect 14590 25218 14642 25230
rect 15486 25282 15538 25294
rect 15486 25218 15538 25230
rect 16046 25282 16098 25294
rect 16046 25218 16098 25230
rect 18062 25282 18114 25294
rect 18062 25218 18114 25230
rect 19406 25282 19458 25294
rect 19406 25218 19458 25230
rect 19518 25282 19570 25294
rect 19518 25218 19570 25230
rect 19630 25282 19682 25294
rect 19630 25218 19682 25230
rect 19854 25282 19906 25294
rect 19854 25218 19906 25230
rect 20302 25282 20354 25294
rect 20302 25218 20354 25230
rect 28366 25282 28418 25294
rect 28366 25218 28418 25230
rect 29822 25282 29874 25294
rect 29822 25218 29874 25230
rect 1344 25114 33760 25148
rect 1344 25062 9278 25114
rect 9330 25062 9382 25114
rect 9434 25062 9486 25114
rect 9538 25062 17342 25114
rect 17394 25062 17446 25114
rect 17498 25062 17550 25114
rect 17602 25062 25406 25114
rect 25458 25062 25510 25114
rect 25562 25062 25614 25114
rect 25666 25062 33470 25114
rect 33522 25062 33574 25114
rect 33626 25062 33678 25114
rect 33730 25062 33760 25114
rect 1344 25028 33760 25062
rect 6862 24946 6914 24958
rect 6862 24882 6914 24894
rect 7646 24946 7698 24958
rect 7646 24882 7698 24894
rect 7758 24946 7810 24958
rect 7758 24882 7810 24894
rect 8318 24946 8370 24958
rect 8318 24882 8370 24894
rect 8542 24946 8594 24958
rect 11678 24946 11730 24958
rect 10546 24894 10558 24946
rect 10610 24894 10622 24946
rect 8542 24882 8594 24894
rect 11678 24882 11730 24894
rect 12574 24946 12626 24958
rect 12574 24882 12626 24894
rect 12686 24946 12738 24958
rect 12686 24882 12738 24894
rect 13246 24946 13298 24958
rect 13246 24882 13298 24894
rect 13358 24946 13410 24958
rect 13358 24882 13410 24894
rect 15486 24946 15538 24958
rect 15486 24882 15538 24894
rect 16494 24946 16546 24958
rect 16494 24882 16546 24894
rect 18398 24946 18450 24958
rect 18398 24882 18450 24894
rect 18846 24946 18898 24958
rect 24658 24894 24670 24946
rect 24722 24894 24734 24946
rect 25554 24894 25566 24946
rect 25618 24894 25630 24946
rect 18846 24882 18898 24894
rect 5294 24834 5346 24846
rect 2482 24782 2494 24834
rect 2546 24782 2558 24834
rect 5294 24770 5346 24782
rect 12798 24834 12850 24846
rect 12798 24770 12850 24782
rect 13470 24834 13522 24846
rect 16718 24834 16770 24846
rect 14354 24782 14366 24834
rect 14418 24782 14430 24834
rect 16258 24782 16270 24834
rect 16322 24782 16334 24834
rect 13470 24770 13522 24782
rect 16718 24770 16770 24782
rect 16830 24834 16882 24846
rect 16830 24770 16882 24782
rect 17390 24834 17442 24846
rect 17390 24770 17442 24782
rect 17502 24834 17554 24846
rect 17502 24770 17554 24782
rect 18286 24834 18338 24846
rect 18286 24770 18338 24782
rect 18734 24834 18786 24846
rect 18734 24770 18786 24782
rect 20190 24834 20242 24846
rect 33182 24834 33234 24846
rect 30706 24782 30718 24834
rect 30770 24782 30782 24834
rect 20190 24770 20242 24782
rect 33182 24770 33234 24782
rect 5518 24722 5570 24734
rect 1810 24670 1822 24722
rect 1874 24670 1886 24722
rect 5518 24658 5570 24670
rect 5966 24722 6018 24734
rect 5966 24658 6018 24670
rect 6414 24722 6466 24734
rect 6414 24658 6466 24670
rect 6750 24722 6802 24734
rect 6750 24658 6802 24670
rect 6974 24722 7026 24734
rect 7534 24722 7586 24734
rect 9774 24722 9826 24734
rect 7298 24670 7310 24722
rect 7362 24670 7374 24722
rect 7970 24670 7982 24722
rect 8034 24670 8046 24722
rect 8866 24670 8878 24722
rect 8930 24670 8942 24722
rect 9538 24670 9550 24722
rect 9602 24670 9614 24722
rect 6974 24658 7026 24670
rect 7534 24658 7586 24670
rect 9774 24658 9826 24670
rect 10894 24722 10946 24734
rect 10894 24658 10946 24670
rect 13134 24722 13186 24734
rect 14926 24722 14978 24734
rect 13906 24670 13918 24722
rect 13970 24670 13982 24722
rect 14578 24670 14590 24722
rect 14642 24670 14654 24722
rect 13134 24658 13186 24670
rect 14926 24658 14978 24670
rect 15374 24722 15426 24734
rect 15374 24658 15426 24670
rect 15598 24722 15650 24734
rect 15598 24658 15650 24670
rect 15934 24722 15986 24734
rect 15934 24658 15986 24670
rect 19294 24722 19346 24734
rect 19294 24658 19346 24670
rect 19518 24722 19570 24734
rect 20414 24722 20466 24734
rect 19842 24670 19854 24722
rect 19906 24670 19918 24722
rect 19518 24658 19570 24670
rect 20414 24658 20466 24670
rect 20638 24722 20690 24734
rect 24334 24722 24386 24734
rect 21186 24670 21198 24722
rect 21250 24670 21262 24722
rect 20638 24658 20690 24670
rect 24334 24658 24386 24670
rect 25230 24722 25282 24734
rect 32510 24722 32562 24734
rect 28130 24670 28142 24722
rect 28194 24670 28206 24722
rect 28914 24670 28926 24722
rect 28978 24670 28990 24722
rect 25230 24658 25282 24670
rect 32510 24658 32562 24670
rect 5406 24610 5458 24622
rect 4610 24558 4622 24610
rect 4674 24558 4686 24610
rect 5406 24546 5458 24558
rect 8430 24610 8482 24622
rect 8430 24546 8482 24558
rect 12238 24610 12290 24622
rect 12238 24546 12290 24558
rect 19406 24610 19458 24622
rect 19406 24546 19458 24558
rect 20302 24610 20354 24622
rect 31950 24610 32002 24622
rect 21858 24558 21870 24610
rect 21922 24558 21934 24610
rect 23986 24558 23998 24610
rect 24050 24558 24062 24610
rect 27346 24558 27358 24610
rect 27410 24558 27422 24610
rect 20302 24546 20354 24558
rect 31950 24546 32002 24558
rect 9998 24498 10050 24510
rect 9998 24434 10050 24446
rect 10110 24498 10162 24510
rect 10110 24434 10162 24446
rect 17502 24498 17554 24510
rect 17502 24434 17554 24446
rect 18846 24498 18898 24510
rect 18846 24434 18898 24446
rect 33070 24498 33122 24510
rect 33070 24434 33122 24446
rect 1344 24330 33600 24364
rect 1344 24278 5246 24330
rect 5298 24278 5350 24330
rect 5402 24278 5454 24330
rect 5506 24278 13310 24330
rect 13362 24278 13414 24330
rect 13466 24278 13518 24330
rect 13570 24278 21374 24330
rect 21426 24278 21478 24330
rect 21530 24278 21582 24330
rect 21634 24278 29438 24330
rect 29490 24278 29542 24330
rect 29594 24278 29646 24330
rect 29698 24278 33600 24330
rect 1344 24244 33600 24278
rect 23102 24162 23154 24174
rect 6402 24110 6414 24162
rect 6466 24110 6478 24162
rect 19058 24110 19070 24162
rect 19122 24110 19134 24162
rect 23102 24098 23154 24110
rect 26798 24162 26850 24174
rect 26798 24098 26850 24110
rect 30830 24162 30882 24174
rect 30830 24098 30882 24110
rect 5966 24050 6018 24062
rect 4722 23998 4734 24050
rect 4786 23998 4798 24050
rect 5966 23986 6018 23998
rect 7758 24050 7810 24062
rect 27022 24050 27074 24062
rect 26338 23998 26350 24050
rect 26402 23998 26414 24050
rect 7758 23986 7810 23998
rect 27022 23986 27074 23998
rect 6190 23938 6242 23950
rect 7870 23938 7922 23950
rect 8766 23938 8818 23950
rect 1810 23886 1822 23938
rect 1874 23886 1886 23938
rect 6626 23886 6638 23938
rect 6690 23886 6702 23938
rect 7186 23886 7198 23938
rect 7250 23886 7262 23938
rect 8194 23886 8206 23938
rect 8258 23886 8270 23938
rect 6190 23874 6242 23886
rect 7870 23874 7922 23886
rect 8766 23874 8818 23886
rect 10110 23938 10162 23950
rect 10110 23874 10162 23886
rect 10446 23938 10498 23950
rect 10446 23874 10498 23886
rect 11006 23938 11058 23950
rect 15598 23938 15650 23950
rect 15250 23886 15262 23938
rect 15314 23886 15326 23938
rect 11006 23874 11058 23886
rect 15598 23874 15650 23886
rect 16270 23938 16322 23950
rect 16270 23874 16322 23886
rect 18174 23938 18226 23950
rect 18174 23874 18226 23886
rect 18510 23938 18562 23950
rect 20078 23938 20130 23950
rect 27358 23938 27410 23950
rect 18722 23886 18734 23938
rect 18786 23886 18798 23938
rect 19170 23886 19182 23938
rect 19234 23886 19246 23938
rect 19842 23886 19854 23938
rect 19906 23886 19918 23938
rect 20402 23886 20414 23938
rect 20466 23886 20478 23938
rect 23426 23886 23438 23938
rect 23490 23886 23502 23938
rect 18510 23874 18562 23886
rect 20078 23874 20130 23886
rect 27358 23874 27410 23886
rect 28030 23938 28082 23950
rect 29150 23938 29202 23950
rect 28466 23886 28478 23938
rect 28530 23886 28542 23938
rect 30258 23886 30270 23938
rect 30322 23886 30334 23938
rect 33170 23886 33182 23938
rect 33234 23886 33246 23938
rect 28030 23874 28082 23886
rect 29150 23874 29202 23886
rect 5854 23826 5906 23838
rect 10670 23826 10722 23838
rect 16158 23826 16210 23838
rect 19630 23826 19682 23838
rect 22878 23826 22930 23838
rect 27246 23826 27298 23838
rect 2482 23774 2494 23826
rect 2546 23774 2558 23826
rect 6962 23774 6974 23826
rect 7026 23774 7038 23826
rect 11554 23774 11566 23826
rect 11618 23774 11630 23826
rect 11890 23774 11902 23826
rect 11954 23774 11966 23826
rect 12562 23774 12574 23826
rect 12626 23774 12638 23826
rect 13906 23774 13918 23826
rect 13970 23774 13982 23826
rect 15026 23774 15038 23826
rect 15090 23774 15102 23826
rect 16594 23774 16606 23826
rect 16658 23774 16670 23826
rect 21298 23774 21310 23826
rect 21362 23774 21374 23826
rect 22418 23774 22430 23826
rect 22482 23774 22494 23826
rect 24210 23774 24222 23826
rect 24274 23774 24286 23826
rect 5854 23762 5906 23774
rect 10670 23762 10722 23774
rect 16158 23762 16210 23774
rect 19630 23762 19682 23774
rect 22878 23762 22930 23774
rect 27246 23762 27298 23774
rect 27582 23826 27634 23838
rect 32734 23826 32786 23838
rect 29474 23774 29486 23826
rect 29538 23774 29550 23826
rect 27582 23762 27634 23774
rect 32734 23762 32786 23774
rect 7646 23714 7698 23726
rect 7646 23650 7698 23662
rect 8430 23714 8482 23726
rect 8430 23650 8482 23662
rect 8654 23714 8706 23726
rect 8654 23650 8706 23662
rect 9886 23714 9938 23726
rect 9886 23650 9938 23662
rect 10222 23714 10274 23726
rect 10222 23650 10274 23662
rect 10782 23714 10834 23726
rect 10782 23650 10834 23662
rect 11230 23714 11282 23726
rect 11230 23650 11282 23662
rect 12238 23714 12290 23726
rect 12238 23650 12290 23662
rect 12910 23714 12962 23726
rect 12910 23650 12962 23662
rect 13582 23714 13634 23726
rect 13582 23650 13634 23662
rect 14254 23714 14306 23726
rect 14254 23650 14306 23662
rect 14702 23714 14754 23726
rect 14702 23650 14754 23662
rect 16046 23714 16098 23726
rect 16046 23650 16098 23662
rect 16942 23714 16994 23726
rect 16942 23650 16994 23662
rect 17614 23714 17666 23726
rect 17614 23650 17666 23662
rect 17838 23714 17890 23726
rect 17838 23650 17890 23662
rect 19294 23714 19346 23726
rect 21646 23714 21698 23726
rect 20066 23662 20078 23714
rect 20130 23662 20142 23714
rect 19294 23650 19346 23662
rect 21646 23650 21698 23662
rect 22094 23714 22146 23726
rect 22094 23650 22146 23662
rect 22990 23714 23042 23726
rect 22990 23650 23042 23662
rect 32622 23714 32674 23726
rect 32622 23650 32674 23662
rect 32958 23714 33010 23726
rect 32958 23650 33010 23662
rect 1344 23546 33760 23580
rect 1344 23494 9278 23546
rect 9330 23494 9382 23546
rect 9434 23494 9486 23546
rect 9538 23494 17342 23546
rect 17394 23494 17446 23546
rect 17498 23494 17550 23546
rect 17602 23494 25406 23546
rect 25458 23494 25510 23546
rect 25562 23494 25614 23546
rect 25666 23494 33470 23546
rect 33522 23494 33574 23546
rect 33626 23494 33678 23546
rect 33730 23494 33760 23546
rect 1344 23460 33760 23494
rect 5406 23378 5458 23390
rect 5406 23314 5458 23326
rect 6974 23378 7026 23390
rect 6974 23314 7026 23326
rect 8654 23378 8706 23390
rect 21310 23378 21362 23390
rect 29486 23378 29538 23390
rect 20402 23326 20414 23378
rect 20466 23326 20478 23378
rect 22306 23326 22318 23378
rect 22370 23326 22382 23378
rect 8654 23314 8706 23326
rect 21310 23314 21362 23326
rect 29486 23314 29538 23326
rect 30942 23378 30994 23390
rect 30942 23314 30994 23326
rect 4846 23266 4898 23278
rect 4846 23202 4898 23214
rect 5294 23266 5346 23278
rect 5294 23202 5346 23214
rect 5518 23266 5570 23278
rect 6750 23266 6802 23278
rect 5842 23214 5854 23266
rect 5906 23214 5918 23266
rect 5518 23202 5570 23214
rect 6750 23202 6802 23214
rect 7758 23266 7810 23278
rect 7758 23202 7810 23214
rect 8878 23266 8930 23278
rect 8878 23202 8930 23214
rect 8990 23266 9042 23278
rect 8990 23202 9042 23214
rect 9550 23266 9602 23278
rect 18734 23266 18786 23278
rect 12338 23214 12350 23266
rect 12402 23214 12414 23266
rect 18498 23214 18510 23266
rect 18562 23214 18574 23266
rect 9550 23202 9602 23214
rect 18734 23202 18786 23214
rect 21534 23266 21586 23278
rect 28478 23266 28530 23278
rect 22642 23214 22654 23266
rect 22706 23214 22718 23266
rect 22978 23214 22990 23266
rect 23042 23214 23054 23266
rect 21534 23202 21586 23214
rect 28478 23202 28530 23214
rect 29374 23266 29426 23278
rect 29374 23202 29426 23214
rect 33182 23266 33234 23278
rect 33182 23202 33234 23214
rect 6190 23154 6242 23166
rect 6190 23090 6242 23102
rect 6638 23154 6690 23166
rect 6638 23090 6690 23102
rect 7198 23154 7250 23166
rect 7198 23090 7250 23102
rect 7310 23154 7362 23166
rect 7310 23090 7362 23102
rect 7422 23154 7474 23166
rect 18286 23154 18338 23166
rect 9762 23102 9774 23154
rect 9826 23102 9838 23154
rect 11554 23102 11566 23154
rect 11618 23102 11630 23154
rect 7422 23090 7474 23102
rect 18286 23090 18338 23102
rect 18398 23154 18450 23166
rect 18398 23090 18450 23102
rect 19070 23154 19122 23166
rect 19070 23090 19122 23102
rect 19966 23154 20018 23166
rect 21646 23154 21698 23166
rect 23326 23154 23378 23166
rect 20626 23102 20638 23154
rect 20690 23102 20702 23154
rect 22530 23102 22542 23154
rect 22594 23102 22606 23154
rect 19966 23090 20018 23102
rect 21646 23090 21698 23102
rect 23326 23090 23378 23102
rect 23886 23154 23938 23166
rect 28254 23154 28306 23166
rect 25554 23102 25566 23154
rect 25618 23102 25630 23154
rect 23886 23090 23938 23102
rect 28254 23090 28306 23102
rect 28702 23154 28754 23166
rect 29922 23102 29934 23154
rect 29986 23102 29998 23154
rect 28702 23090 28754 23102
rect 16718 23042 16770 23054
rect 16718 22978 16770 22990
rect 17502 23042 17554 23054
rect 17502 22978 17554 22990
rect 24446 23042 24498 23054
rect 27458 22990 27470 23042
rect 27522 22990 27534 23042
rect 24446 22978 24498 22990
rect 15822 22930 15874 22942
rect 15822 22866 15874 22878
rect 16270 22930 16322 22942
rect 16270 22866 16322 22878
rect 16494 22930 16546 22942
rect 16494 22866 16546 22878
rect 19182 22930 19234 22942
rect 19182 22866 19234 22878
rect 19518 22930 19570 22942
rect 19518 22866 19570 22878
rect 19630 22930 19682 22942
rect 19630 22866 19682 22878
rect 19854 22930 19906 22942
rect 19854 22866 19906 22878
rect 28142 22930 28194 22942
rect 28142 22866 28194 22878
rect 28926 22930 28978 22942
rect 28926 22866 28978 22878
rect 29486 22930 29538 22942
rect 29486 22866 29538 22878
rect 33070 22930 33122 22942
rect 33070 22866 33122 22878
rect 1344 22762 33600 22796
rect 1344 22710 5246 22762
rect 5298 22710 5350 22762
rect 5402 22710 5454 22762
rect 5506 22710 13310 22762
rect 13362 22710 13414 22762
rect 13466 22710 13518 22762
rect 13570 22710 21374 22762
rect 21426 22710 21478 22762
rect 21530 22710 21582 22762
rect 21634 22710 29438 22762
rect 29490 22710 29542 22762
rect 29594 22710 29646 22762
rect 29698 22710 33600 22762
rect 1344 22676 33600 22710
rect 11342 22594 11394 22606
rect 11342 22530 11394 22542
rect 15038 22594 15090 22606
rect 15038 22530 15090 22542
rect 15374 22594 15426 22606
rect 20750 22594 20802 22606
rect 18050 22542 18062 22594
rect 18114 22591 18126 22594
rect 18610 22591 18622 22594
rect 18114 22545 18622 22591
rect 18114 22542 18126 22545
rect 18610 22542 18622 22545
rect 18674 22542 18686 22594
rect 15374 22530 15426 22542
rect 20750 22530 20802 22542
rect 32958 22594 33010 22606
rect 32958 22530 33010 22542
rect 5070 22482 5122 22494
rect 14814 22482 14866 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 5842 22430 5854 22482
rect 5906 22430 5918 22482
rect 5070 22418 5122 22430
rect 14814 22418 14866 22430
rect 18622 22482 18674 22494
rect 24882 22430 24894 22482
rect 24946 22430 24958 22482
rect 25554 22430 25566 22482
rect 25618 22430 25630 22482
rect 27570 22430 27582 22482
rect 27634 22430 27646 22482
rect 18622 22418 18674 22430
rect 12910 22370 12962 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 10882 22318 10894 22370
rect 10946 22318 10958 22370
rect 12910 22306 12962 22318
rect 16158 22370 16210 22382
rect 16158 22306 16210 22318
rect 16270 22370 16322 22382
rect 18846 22370 18898 22382
rect 25454 22370 25506 22382
rect 28142 22370 28194 22382
rect 16706 22318 16718 22370
rect 16770 22318 16782 22370
rect 19170 22318 19182 22370
rect 19234 22318 19246 22370
rect 21970 22318 21982 22370
rect 22034 22318 22046 22370
rect 25890 22318 25902 22370
rect 25954 22318 25966 22370
rect 16270 22306 16322 22318
rect 18846 22306 18898 22318
rect 25454 22306 25506 22318
rect 28142 22306 28194 22318
rect 29486 22370 29538 22382
rect 29486 22306 29538 22318
rect 30270 22370 30322 22382
rect 31042 22318 31054 22370
rect 31106 22318 31118 22370
rect 30270 22306 30322 22318
rect 11454 22258 11506 22270
rect 13470 22258 13522 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 11778 22206 11790 22258
rect 11842 22206 11854 22258
rect 12562 22206 12574 22258
rect 12626 22206 12638 22258
rect 11454 22194 11506 22206
rect 13470 22194 13522 22206
rect 13806 22258 13858 22270
rect 13806 22194 13858 22206
rect 14142 22258 14194 22270
rect 14142 22194 14194 22206
rect 14478 22258 14530 22270
rect 20638 22258 20690 22270
rect 17378 22206 17390 22258
rect 17442 22206 17454 22258
rect 14478 22194 14530 22206
rect 20638 22194 20690 22206
rect 21646 22258 21698 22270
rect 26798 22258 26850 22270
rect 22754 22206 22766 22258
rect 22818 22206 22830 22258
rect 21646 22194 21698 22206
rect 26798 22194 26850 22206
rect 27134 22258 27186 22270
rect 27918 22258 27970 22270
rect 27234 22206 27246 22258
rect 27298 22206 27310 22258
rect 27134 22194 27186 22206
rect 27918 22194 27970 22206
rect 28478 22258 28530 22270
rect 28478 22194 28530 22206
rect 29934 22258 29986 22270
rect 30146 22206 30158 22258
rect 30210 22206 30222 22258
rect 29934 22194 29986 22206
rect 11342 22146 11394 22158
rect 11342 22082 11394 22094
rect 12126 22146 12178 22158
rect 12126 22082 12178 22094
rect 15822 22146 15874 22158
rect 15822 22082 15874 22094
rect 16382 22146 16434 22158
rect 16382 22082 16434 22094
rect 17054 22146 17106 22158
rect 17054 22082 17106 22094
rect 18174 22146 18226 22158
rect 18174 22082 18226 22094
rect 19406 22146 19458 22158
rect 19406 22082 19458 22094
rect 19518 22146 19570 22158
rect 19518 22082 19570 22094
rect 19966 22146 20018 22158
rect 19966 22082 20018 22094
rect 20414 22146 20466 22158
rect 20414 22082 20466 22094
rect 21310 22146 21362 22158
rect 21310 22082 21362 22094
rect 21534 22146 21586 22158
rect 21534 22082 21586 22094
rect 25118 22146 25170 22158
rect 25118 22082 25170 22094
rect 27022 22146 27074 22158
rect 27022 22082 27074 22094
rect 28366 22146 28418 22158
rect 28366 22082 28418 22094
rect 29262 22146 29314 22158
rect 29262 22082 29314 22094
rect 1344 21978 33760 22012
rect 1344 21926 9278 21978
rect 9330 21926 9382 21978
rect 9434 21926 9486 21978
rect 9538 21926 17342 21978
rect 17394 21926 17446 21978
rect 17498 21926 17550 21978
rect 17602 21926 25406 21978
rect 25458 21926 25510 21978
rect 25562 21926 25614 21978
rect 25666 21926 33470 21978
rect 33522 21926 33574 21978
rect 33626 21926 33678 21978
rect 33730 21926 33760 21978
rect 1344 21892 33760 21926
rect 5294 21810 5346 21822
rect 5294 21746 5346 21758
rect 6190 21810 6242 21822
rect 6190 21746 6242 21758
rect 6750 21810 6802 21822
rect 13246 21810 13298 21822
rect 16046 21810 16098 21822
rect 11330 21758 11342 21810
rect 11394 21758 11406 21810
rect 14354 21758 14366 21810
rect 14418 21758 14430 21810
rect 6750 21746 6802 21758
rect 13246 21746 13298 21758
rect 16046 21746 16098 21758
rect 16494 21810 16546 21822
rect 16494 21746 16546 21758
rect 23774 21810 23826 21822
rect 23774 21746 23826 21758
rect 23886 21810 23938 21822
rect 23886 21746 23938 21758
rect 6078 21698 6130 21710
rect 6078 21634 6130 21646
rect 7534 21698 7586 21710
rect 7534 21634 7586 21646
rect 7646 21698 7698 21710
rect 7646 21634 7698 21646
rect 9550 21698 9602 21710
rect 9550 21634 9602 21646
rect 9662 21698 9714 21710
rect 9662 21634 9714 21646
rect 12910 21698 12962 21710
rect 12910 21634 12962 21646
rect 13022 21698 13074 21710
rect 13022 21634 13074 21646
rect 22878 21698 22930 21710
rect 22878 21634 22930 21646
rect 24222 21698 24274 21710
rect 24222 21634 24274 21646
rect 24446 21698 24498 21710
rect 24446 21634 24498 21646
rect 24670 21698 24722 21710
rect 24670 21634 24722 21646
rect 25342 21698 25394 21710
rect 27122 21646 27134 21698
rect 27186 21646 27198 21698
rect 28242 21646 28254 21698
rect 28306 21646 28318 21698
rect 32050 21646 32062 21698
rect 32114 21646 32126 21698
rect 25342 21634 25394 21646
rect 4958 21586 5010 21598
rect 1810 21534 1822 21586
rect 1874 21534 1886 21586
rect 4958 21522 5010 21534
rect 5294 21586 5346 21598
rect 5294 21522 5346 21534
rect 5630 21586 5682 21598
rect 5630 21522 5682 21534
rect 6638 21586 6690 21598
rect 6638 21522 6690 21534
rect 6974 21586 7026 21598
rect 6974 21522 7026 21534
rect 7310 21586 7362 21598
rect 7310 21522 7362 21534
rect 7870 21586 7922 21598
rect 7870 21522 7922 21534
rect 8318 21586 8370 21598
rect 8318 21522 8370 21534
rect 8430 21586 8482 21598
rect 8430 21522 8482 21534
rect 9886 21586 9938 21598
rect 12574 21586 12626 21598
rect 14814 21586 14866 21598
rect 23214 21586 23266 21598
rect 11106 21534 11118 21586
rect 11170 21534 11182 21586
rect 12114 21534 12126 21586
rect 12178 21534 12190 21586
rect 14130 21534 14142 21586
rect 14194 21534 14206 21586
rect 18722 21534 18734 21586
rect 18786 21534 18798 21586
rect 9886 21522 9938 21534
rect 12574 21522 12626 21534
rect 14814 21522 14866 21534
rect 23214 21522 23266 21534
rect 23662 21586 23714 21598
rect 23662 21522 23714 21534
rect 25230 21586 25282 21598
rect 30270 21586 30322 21598
rect 25778 21534 25790 21586
rect 25842 21534 25854 21586
rect 26898 21534 26910 21586
rect 26962 21534 26974 21586
rect 29810 21534 29822 21586
rect 29874 21534 29886 21586
rect 25230 21522 25282 21534
rect 30270 21522 30322 21534
rect 8094 21474 8146 21486
rect 2482 21422 2494 21474
rect 2546 21422 2558 21474
rect 4610 21422 4622 21474
rect 4674 21422 4686 21474
rect 8094 21410 8146 21422
rect 10334 21474 10386 21486
rect 10334 21410 10386 21422
rect 13694 21474 13746 21486
rect 13694 21410 13746 21422
rect 15486 21474 15538 21486
rect 15486 21410 15538 21422
rect 16942 21474 16994 21486
rect 16942 21410 16994 21422
rect 17614 21474 17666 21486
rect 17614 21410 17666 21422
rect 17950 21474 18002 21486
rect 17950 21410 18002 21422
rect 18398 21474 18450 21486
rect 21646 21474 21698 21486
rect 19506 21422 19518 21474
rect 19570 21422 19582 21474
rect 18398 21410 18450 21422
rect 21646 21410 21698 21422
rect 22318 21474 22370 21486
rect 30718 21474 30770 21486
rect 33182 21474 33234 21486
rect 26114 21422 26126 21474
rect 26178 21422 26190 21474
rect 27010 21422 27022 21474
rect 27074 21422 27086 21474
rect 31714 21422 31726 21474
rect 31778 21422 31790 21474
rect 22318 21410 22370 21422
rect 30718 21410 30770 21422
rect 33182 21410 33234 21422
rect 6190 21362 6242 21374
rect 6190 21298 6242 21310
rect 22654 21362 22706 21374
rect 22654 21298 22706 21310
rect 22990 21362 23042 21374
rect 22990 21298 23042 21310
rect 24782 21362 24834 21374
rect 31826 21310 31838 21362
rect 31890 21310 31902 21362
rect 24782 21298 24834 21310
rect 1344 21194 33600 21228
rect 1344 21142 5246 21194
rect 5298 21142 5350 21194
rect 5402 21142 5454 21194
rect 5506 21142 13310 21194
rect 13362 21142 13414 21194
rect 13466 21142 13518 21194
rect 13570 21142 21374 21194
rect 21426 21142 21478 21194
rect 21530 21142 21582 21194
rect 21634 21142 29438 21194
rect 29490 21142 29542 21194
rect 29594 21142 29646 21194
rect 29698 21142 33600 21194
rect 1344 21108 33600 21142
rect 5742 21026 5794 21038
rect 5742 20962 5794 20974
rect 4174 20914 4226 20926
rect 4174 20850 4226 20862
rect 5070 20914 5122 20926
rect 12014 20914 12066 20926
rect 17390 20914 17442 20926
rect 7970 20862 7982 20914
rect 8034 20862 8046 20914
rect 10098 20862 10110 20914
rect 10162 20862 10174 20914
rect 16370 20862 16382 20914
rect 16434 20862 16446 20914
rect 5070 20850 5122 20862
rect 12014 20850 12066 20862
rect 17390 20850 17442 20862
rect 19294 20914 19346 20926
rect 19294 20850 19346 20862
rect 20862 20914 20914 20926
rect 27246 20914 27298 20926
rect 24210 20862 24222 20914
rect 24274 20862 24286 20914
rect 26114 20862 26126 20914
rect 26178 20862 26190 20914
rect 20862 20850 20914 20862
rect 27246 20850 27298 20862
rect 27694 20914 27746 20926
rect 33294 20914 33346 20926
rect 30370 20862 30382 20914
rect 30434 20862 30446 20914
rect 27694 20850 27746 20862
rect 33294 20850 33346 20862
rect 4286 20802 4338 20814
rect 4286 20738 4338 20750
rect 4622 20802 4674 20814
rect 4622 20738 4674 20750
rect 5854 20802 5906 20814
rect 5854 20738 5906 20750
rect 6190 20802 6242 20814
rect 6190 20738 6242 20750
rect 6638 20802 6690 20814
rect 6638 20738 6690 20750
rect 6862 20802 6914 20814
rect 17838 20802 17890 20814
rect 7186 20750 7198 20802
rect 7250 20750 7262 20802
rect 13458 20750 13470 20802
rect 13522 20750 13534 20802
rect 6862 20738 6914 20750
rect 17838 20738 17890 20750
rect 18286 20802 18338 20814
rect 18286 20738 18338 20750
rect 19182 20802 19234 20814
rect 19182 20738 19234 20750
rect 19518 20802 19570 20814
rect 20302 20802 20354 20814
rect 27358 20802 27410 20814
rect 19954 20750 19966 20802
rect 20018 20750 20030 20802
rect 21410 20750 21422 20802
rect 21474 20750 21486 20802
rect 25330 20750 25342 20802
rect 25394 20750 25406 20802
rect 25666 20750 25678 20802
rect 25730 20750 25742 20802
rect 26898 20750 26910 20802
rect 26962 20750 26974 20802
rect 19518 20738 19570 20750
rect 20302 20738 20354 20750
rect 27358 20738 27410 20750
rect 27918 20802 27970 20814
rect 28354 20750 28366 20802
rect 28418 20750 28430 20802
rect 29138 20750 29150 20802
rect 29202 20750 29214 20802
rect 32050 20750 32062 20802
rect 32114 20750 32126 20802
rect 27918 20738 27970 20750
rect 4062 20690 4114 20702
rect 4062 20626 4114 20638
rect 11006 20690 11058 20702
rect 17614 20690 17666 20702
rect 14242 20638 14254 20690
rect 14306 20638 14318 20690
rect 11006 20626 11058 20638
rect 17614 20626 17666 20638
rect 18846 20690 18898 20702
rect 18846 20626 18898 20638
rect 19742 20690 19794 20702
rect 27134 20690 27186 20702
rect 22082 20638 22094 20690
rect 22146 20638 22158 20690
rect 26786 20638 26798 20690
rect 26850 20638 26862 20690
rect 28130 20638 28142 20690
rect 28194 20638 28206 20690
rect 32386 20638 32398 20690
rect 32450 20638 32462 20690
rect 32722 20638 32734 20690
rect 32786 20638 32798 20690
rect 19742 20626 19794 20638
rect 27134 20626 27186 20638
rect 5742 20578 5794 20590
rect 5742 20514 5794 20526
rect 6526 20578 6578 20590
rect 6526 20514 6578 20526
rect 10670 20578 10722 20590
rect 10670 20514 10722 20526
rect 10894 20578 10946 20590
rect 10894 20514 10946 20526
rect 11566 20578 11618 20590
rect 11566 20514 11618 20526
rect 16830 20578 16882 20590
rect 16830 20514 16882 20526
rect 18062 20578 18114 20590
rect 18062 20514 18114 20526
rect 19630 20578 19682 20590
rect 19630 20514 19682 20526
rect 24670 20578 24722 20590
rect 24670 20514 24722 20526
rect 24894 20578 24946 20590
rect 24894 20514 24946 20526
rect 28702 20578 28754 20590
rect 28702 20514 28754 20526
rect 1344 20410 33760 20444
rect 1344 20358 9278 20410
rect 9330 20358 9382 20410
rect 9434 20358 9486 20410
rect 9538 20358 17342 20410
rect 17394 20358 17446 20410
rect 17498 20358 17550 20410
rect 17602 20358 25406 20410
rect 25458 20358 25510 20410
rect 25562 20358 25614 20410
rect 25666 20358 33470 20410
rect 33522 20358 33574 20410
rect 33626 20358 33678 20410
rect 33730 20358 33760 20410
rect 1344 20324 33760 20358
rect 4286 20242 4338 20254
rect 4286 20178 4338 20190
rect 4510 20242 4562 20254
rect 14366 20242 14418 20254
rect 5394 20190 5406 20242
rect 5458 20190 5470 20242
rect 4510 20178 4562 20190
rect 14366 20178 14418 20190
rect 15262 20242 15314 20254
rect 15262 20178 15314 20190
rect 16158 20242 16210 20254
rect 16158 20178 16210 20190
rect 16942 20242 16994 20254
rect 16942 20178 16994 20190
rect 25342 20242 25394 20254
rect 25666 20190 25678 20242
rect 25730 20190 25742 20242
rect 25342 20178 25394 20190
rect 13022 20130 13074 20142
rect 6514 20078 6526 20130
rect 6578 20078 6590 20130
rect 13022 20066 13074 20078
rect 13694 20130 13746 20142
rect 20974 20130 21026 20142
rect 18162 20078 18174 20130
rect 18226 20078 18238 20130
rect 13694 20066 13746 20078
rect 20974 20066 21026 20078
rect 22430 20130 22482 20142
rect 22430 20066 22482 20078
rect 22542 20130 22594 20142
rect 22542 20066 22594 20078
rect 22878 20130 22930 20142
rect 30494 20130 30546 20142
rect 27234 20078 27246 20130
rect 27298 20078 27310 20130
rect 28354 20078 28366 20130
rect 28418 20078 28430 20130
rect 31826 20078 31838 20130
rect 31890 20078 31902 20130
rect 32162 20078 32174 20130
rect 32226 20078 32238 20130
rect 22878 20066 22930 20078
rect 30494 20066 30546 20078
rect 4622 20018 4674 20030
rect 13582 20018 13634 20030
rect 5170 19966 5182 20018
rect 5234 19966 5246 20018
rect 5730 19966 5742 20018
rect 5794 19966 5806 20018
rect 9762 19966 9774 20018
rect 9826 19966 9838 20018
rect 4622 19954 4674 19966
rect 13582 19954 13634 19966
rect 13918 20018 13970 20030
rect 13918 19954 13970 19966
rect 14142 20018 14194 20030
rect 14142 19954 14194 19966
rect 14366 20018 14418 20030
rect 14366 19954 14418 19966
rect 14590 20018 14642 20030
rect 14590 19954 14642 19966
rect 15038 20018 15090 20030
rect 15038 19954 15090 19966
rect 15374 20018 15426 20030
rect 15374 19954 15426 19966
rect 16046 20018 16098 20030
rect 16046 19954 16098 19966
rect 16382 20018 16434 20030
rect 23102 20018 23154 20030
rect 17490 19966 17502 20018
rect 17554 19966 17566 20018
rect 16382 19954 16434 19966
rect 23102 19954 23154 19966
rect 23550 20018 23602 20030
rect 23550 19954 23602 19966
rect 23774 20018 23826 20030
rect 33182 20018 33234 20030
rect 27346 19966 27358 20018
rect 27410 19966 27422 20018
rect 29810 19966 29822 20018
rect 29874 19966 29886 20018
rect 30258 19966 30270 20018
rect 30322 19966 30334 20018
rect 31042 19966 31054 20018
rect 31106 19966 31118 20018
rect 31490 19966 31502 20018
rect 31554 19966 31566 20018
rect 32498 19966 32510 20018
rect 32562 19966 32574 20018
rect 23774 19954 23826 19966
rect 33182 19954 33234 19966
rect 21534 19906 21586 19918
rect 8642 19854 8654 19906
rect 8706 19854 8718 19906
rect 10434 19854 10446 19906
rect 10498 19854 10510 19906
rect 12562 19854 12574 19906
rect 12626 19854 12638 19906
rect 20290 19854 20302 19906
rect 20354 19854 20366 19906
rect 21534 19842 21586 19854
rect 21982 19906 22034 19918
rect 21982 19842 22034 19854
rect 22990 19906 23042 19918
rect 26238 19906 26290 19918
rect 24210 19854 24222 19906
rect 24274 19854 24286 19906
rect 27010 19854 27022 19906
rect 27074 19854 27086 19906
rect 22990 19842 23042 19854
rect 26238 19842 26290 19854
rect 22430 19794 22482 19806
rect 22430 19730 22482 19742
rect 26014 19794 26066 19806
rect 26014 19730 26066 19742
rect 33070 19794 33122 19806
rect 33070 19730 33122 19742
rect 1344 19626 33600 19660
rect 1344 19574 5246 19626
rect 5298 19574 5350 19626
rect 5402 19574 5454 19626
rect 5506 19574 13310 19626
rect 13362 19574 13414 19626
rect 13466 19574 13518 19626
rect 13570 19574 21374 19626
rect 21426 19574 21478 19626
rect 21530 19574 21582 19626
rect 21634 19574 29438 19626
rect 29490 19574 29542 19626
rect 29594 19574 29646 19626
rect 29698 19574 33600 19626
rect 1344 19540 33600 19574
rect 5742 19458 5794 19470
rect 23774 19458 23826 19470
rect 18834 19406 18846 19458
rect 18898 19455 18910 19458
rect 19954 19455 19966 19458
rect 18898 19409 19966 19455
rect 18898 19406 18910 19409
rect 19954 19406 19966 19409
rect 20018 19406 20030 19458
rect 20290 19406 20302 19458
rect 20354 19455 20366 19458
rect 20514 19455 20526 19458
rect 20354 19409 20526 19455
rect 20354 19406 20366 19409
rect 20514 19406 20526 19409
rect 20578 19406 20590 19458
rect 22082 19406 22094 19458
rect 22146 19455 22158 19458
rect 22866 19455 22878 19458
rect 22146 19409 22878 19455
rect 22146 19406 22158 19409
rect 22866 19406 22878 19409
rect 22930 19406 22942 19458
rect 5742 19394 5794 19406
rect 23774 19394 23826 19406
rect 24334 19458 24386 19470
rect 24334 19394 24386 19406
rect 29150 19458 29202 19470
rect 29150 19394 29202 19406
rect 30830 19458 30882 19470
rect 30830 19394 30882 19406
rect 5070 19346 5122 19358
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 5070 19282 5122 19294
rect 9550 19346 9602 19358
rect 9550 19282 9602 19294
rect 10558 19346 10610 19358
rect 10558 19282 10610 19294
rect 12910 19346 12962 19358
rect 19070 19346 19122 19358
rect 17042 19294 17054 19346
rect 17106 19294 17118 19346
rect 12910 19282 12962 19294
rect 19070 19282 19122 19294
rect 19406 19346 19458 19358
rect 19406 19282 19458 19294
rect 19966 19346 20018 19358
rect 19966 19282 20018 19294
rect 20302 19346 20354 19358
rect 20302 19282 20354 19294
rect 21870 19346 21922 19358
rect 32846 19346 32898 19358
rect 25106 19294 25118 19346
rect 25170 19294 25182 19346
rect 27794 19294 27806 19346
rect 27858 19294 27870 19346
rect 21870 19282 21922 19294
rect 32846 19282 32898 19294
rect 5854 19234 5906 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 5854 19170 5906 19182
rect 7870 19234 7922 19246
rect 7870 19170 7922 19182
rect 8766 19234 8818 19246
rect 8766 19170 8818 19182
rect 10334 19234 10386 19246
rect 10334 19170 10386 19182
rect 10670 19234 10722 19246
rect 10670 19170 10722 19182
rect 10894 19234 10946 19246
rect 10894 19170 10946 19182
rect 13582 19234 13634 19246
rect 22990 19234 23042 19246
rect 14130 19182 14142 19234
rect 14194 19182 14206 19234
rect 17490 19182 17502 19234
rect 17554 19182 17566 19234
rect 13582 19170 13634 19182
rect 22990 19170 23042 19182
rect 23886 19234 23938 19246
rect 23886 19170 23938 19182
rect 24446 19234 24498 19246
rect 26014 19234 26066 19246
rect 29486 19234 29538 19246
rect 24994 19182 25006 19234
rect 25058 19182 25070 19234
rect 26786 19182 26798 19234
rect 26850 19182 26862 19234
rect 28018 19182 28030 19234
rect 28082 19182 28094 19234
rect 30034 19182 30046 19234
rect 30098 19182 30110 19234
rect 24446 19170 24498 19182
rect 26014 19170 26066 19182
rect 29486 19170 29538 19182
rect 8206 19122 8258 19134
rect 2482 19070 2494 19122
rect 2546 19070 2558 19122
rect 8206 19058 8258 19070
rect 8990 19122 9042 19134
rect 8990 19058 9042 19070
rect 9102 19122 9154 19134
rect 9102 19058 9154 19070
rect 11454 19122 11506 19134
rect 11454 19058 11506 19070
rect 11566 19122 11618 19134
rect 23326 19122 23378 19134
rect 14914 19070 14926 19122
rect 14978 19070 14990 19122
rect 17714 19070 17726 19122
rect 17778 19070 17790 19122
rect 11566 19058 11618 19070
rect 23326 19058 23378 19070
rect 24334 19122 24386 19134
rect 26238 19122 26290 19134
rect 25442 19070 25454 19122
rect 25506 19070 25518 19122
rect 24334 19058 24386 19070
rect 26238 19058 26290 19070
rect 26350 19122 26402 19134
rect 28366 19122 28418 19134
rect 27682 19070 27694 19122
rect 27746 19070 27758 19122
rect 26350 19058 26402 19070
rect 28366 19058 28418 19070
rect 5742 19010 5794 19022
rect 5742 18946 5794 18958
rect 8094 19010 8146 19022
rect 8094 18946 8146 18958
rect 11230 19010 11282 19022
rect 11230 18946 11282 18958
rect 13694 19010 13746 19022
rect 13694 18946 13746 18958
rect 13918 19010 13970 19022
rect 13918 18946 13970 18958
rect 18286 19010 18338 19022
rect 18286 18946 18338 18958
rect 20750 19010 20802 19022
rect 20750 18946 20802 18958
rect 21534 19010 21586 19022
rect 21534 18946 21586 18958
rect 22318 19010 22370 19022
rect 22318 18946 22370 18958
rect 22878 19010 22930 19022
rect 22878 18946 22930 18958
rect 23214 19010 23266 19022
rect 23214 18946 23266 18958
rect 23774 19010 23826 19022
rect 23774 18946 23826 18958
rect 26126 19010 26178 19022
rect 26126 18946 26178 18958
rect 28478 19010 28530 19022
rect 28478 18946 28530 18958
rect 28702 19010 28754 19022
rect 28702 18946 28754 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 1344 18842 33760 18876
rect 1344 18790 9278 18842
rect 9330 18790 9382 18842
rect 9434 18790 9486 18842
rect 9538 18790 17342 18842
rect 17394 18790 17446 18842
rect 17498 18790 17550 18842
rect 17602 18790 25406 18842
rect 25458 18790 25510 18842
rect 25562 18790 25614 18842
rect 25666 18790 33470 18842
rect 33522 18790 33574 18842
rect 33626 18790 33678 18842
rect 33730 18790 33760 18842
rect 1344 18756 33760 18790
rect 3054 18674 3106 18686
rect 3054 18610 3106 18622
rect 3614 18674 3666 18686
rect 11790 18674 11842 18686
rect 5954 18622 5966 18674
rect 6018 18622 6030 18674
rect 8194 18622 8206 18674
rect 8258 18622 8270 18674
rect 3614 18610 3666 18622
rect 11790 18610 11842 18622
rect 13134 18674 13186 18686
rect 13134 18610 13186 18622
rect 14926 18674 14978 18686
rect 14926 18610 14978 18622
rect 15486 18674 15538 18686
rect 15486 18610 15538 18622
rect 18622 18674 18674 18686
rect 27918 18674 27970 18686
rect 26674 18622 26686 18674
rect 26738 18622 26750 18674
rect 18622 18610 18674 18622
rect 27918 18610 27970 18622
rect 33070 18674 33122 18686
rect 33070 18610 33122 18622
rect 2942 18562 2994 18574
rect 2942 18498 2994 18510
rect 3726 18562 3778 18574
rect 3726 18498 3778 18510
rect 5070 18562 5122 18574
rect 5070 18498 5122 18510
rect 5182 18562 5234 18574
rect 5182 18498 5234 18510
rect 7422 18562 7474 18574
rect 7422 18498 7474 18510
rect 11342 18562 11394 18574
rect 11342 18498 11394 18510
rect 11678 18562 11730 18574
rect 11678 18498 11730 18510
rect 13022 18562 13074 18574
rect 13022 18498 13074 18510
rect 13358 18562 13410 18574
rect 13358 18498 13410 18510
rect 15038 18562 15090 18574
rect 15038 18498 15090 18510
rect 15598 18562 15650 18574
rect 15598 18498 15650 18510
rect 16046 18562 16098 18574
rect 16046 18498 16098 18510
rect 16158 18562 16210 18574
rect 16158 18498 16210 18510
rect 19966 18562 20018 18574
rect 24110 18562 24162 18574
rect 27694 18562 27746 18574
rect 22754 18510 22766 18562
rect 22818 18510 22830 18562
rect 26450 18510 26462 18562
rect 26514 18510 26526 18562
rect 27234 18510 27246 18562
rect 27298 18510 27310 18562
rect 19966 18498 20018 18510
rect 24110 18498 24162 18510
rect 27694 18498 27746 18510
rect 30494 18562 30546 18574
rect 31714 18510 31726 18562
rect 31778 18510 31790 18562
rect 32162 18510 32174 18562
rect 32226 18510 32238 18562
rect 30494 18498 30546 18510
rect 3278 18450 3330 18462
rect 3278 18386 3330 18398
rect 3950 18450 4002 18462
rect 3950 18386 4002 18398
rect 4398 18450 4450 18462
rect 4398 18386 4450 18398
rect 4510 18450 4562 18462
rect 4510 18386 4562 18398
rect 4846 18450 4898 18462
rect 4846 18386 4898 18398
rect 6302 18450 6354 18462
rect 6302 18386 6354 18398
rect 6750 18450 6802 18462
rect 6750 18386 6802 18398
rect 7758 18450 7810 18462
rect 7758 18386 7810 18398
rect 8542 18450 8594 18462
rect 8542 18386 8594 18398
rect 8990 18450 9042 18462
rect 8990 18386 9042 18398
rect 10894 18450 10946 18462
rect 10894 18386 10946 18398
rect 11118 18450 11170 18462
rect 11118 18386 11170 18398
rect 12014 18450 12066 18462
rect 12014 18386 12066 18398
rect 13470 18450 13522 18462
rect 13470 18386 13522 18398
rect 13918 18450 13970 18462
rect 13918 18386 13970 18398
rect 14030 18450 14082 18462
rect 14030 18386 14082 18398
rect 14478 18450 14530 18462
rect 14478 18386 14530 18398
rect 14814 18450 14866 18462
rect 14814 18386 14866 18398
rect 15262 18450 15314 18462
rect 15262 18386 15314 18398
rect 15822 18450 15874 18462
rect 15822 18386 15874 18398
rect 19854 18450 19906 18462
rect 19854 18386 19906 18398
rect 20526 18450 20578 18462
rect 21534 18450 21586 18462
rect 21298 18398 21310 18450
rect 21362 18398 21374 18450
rect 20526 18386 20578 18398
rect 21534 18386 21586 18398
rect 21646 18450 21698 18462
rect 23102 18450 23154 18462
rect 23774 18450 23826 18462
rect 22082 18398 22094 18450
rect 22146 18398 22158 18450
rect 23426 18398 23438 18450
rect 23490 18398 23502 18450
rect 21646 18386 21698 18398
rect 23102 18386 23154 18398
rect 23774 18386 23826 18398
rect 24670 18450 24722 18462
rect 25902 18450 25954 18462
rect 25442 18398 25454 18450
rect 25506 18398 25518 18450
rect 24670 18386 24722 18398
rect 25902 18386 25954 18398
rect 26350 18450 26402 18462
rect 26350 18386 26402 18398
rect 28254 18450 28306 18462
rect 29598 18450 29650 18462
rect 28690 18398 28702 18450
rect 28754 18398 28766 18450
rect 28254 18386 28306 18398
rect 29598 18386 29650 18398
rect 30270 18450 30322 18462
rect 30930 18398 30942 18450
rect 30994 18398 31006 18450
rect 31490 18398 31502 18450
rect 31554 18398 31566 18450
rect 32274 18398 32286 18450
rect 32338 18398 32350 18450
rect 30270 18386 30322 18398
rect 4174 18338 4226 18350
rect 4174 18274 4226 18286
rect 11230 18338 11282 18350
rect 11230 18274 11282 18286
rect 13694 18338 13746 18350
rect 13694 18274 13746 18286
rect 18958 18338 19010 18350
rect 18958 18274 19010 18286
rect 20974 18338 21026 18350
rect 29262 18338 29314 18350
rect 28578 18286 28590 18338
rect 28642 18286 28654 18338
rect 20974 18274 21026 18286
rect 29262 18274 29314 18286
rect 30046 18338 30098 18350
rect 33182 18338 33234 18350
rect 30370 18286 30382 18338
rect 30434 18286 30446 18338
rect 30046 18274 30098 18286
rect 33182 18274 33234 18286
rect 3614 18226 3666 18238
rect 3614 18162 3666 18174
rect 19182 18226 19234 18238
rect 19182 18162 19234 18174
rect 19518 18226 19570 18238
rect 19518 18162 19570 18174
rect 19966 18226 20018 18238
rect 19966 18162 20018 18174
rect 23438 18226 23490 18238
rect 23438 18162 23490 18174
rect 27582 18226 27634 18238
rect 27582 18162 27634 18174
rect 29822 18226 29874 18238
rect 29822 18162 29874 18174
rect 1344 18058 33600 18092
rect 1344 18006 5246 18058
rect 5298 18006 5350 18058
rect 5402 18006 5454 18058
rect 5506 18006 13310 18058
rect 13362 18006 13414 18058
rect 13466 18006 13518 18058
rect 13570 18006 21374 18058
rect 21426 18006 21478 18058
rect 21530 18006 21582 18058
rect 21634 18006 29438 18058
rect 29490 18006 29542 18058
rect 29594 18006 29646 18058
rect 29698 18006 33600 18058
rect 1344 17972 33600 18006
rect 20750 17890 20802 17902
rect 20750 17826 20802 17838
rect 27470 17890 27522 17902
rect 27470 17826 27522 17838
rect 27918 17890 27970 17902
rect 31714 17838 31726 17890
rect 31778 17838 31790 17890
rect 27918 17826 27970 17838
rect 5070 17778 5122 17790
rect 16830 17778 16882 17790
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 9874 17726 9886 17778
rect 9938 17726 9950 17778
rect 12002 17726 12014 17778
rect 12066 17726 12078 17778
rect 14242 17726 14254 17778
rect 14306 17726 14318 17778
rect 16370 17726 16382 17778
rect 16434 17726 16446 17778
rect 5070 17714 5122 17726
rect 16830 17714 16882 17726
rect 17614 17778 17666 17790
rect 21982 17778 22034 17790
rect 17826 17726 17838 17778
rect 17890 17726 17902 17778
rect 17614 17714 17666 17726
rect 21982 17714 22034 17726
rect 22206 17778 22258 17790
rect 22206 17714 22258 17726
rect 24782 17778 24834 17790
rect 24782 17714 24834 17726
rect 28590 17778 28642 17790
rect 30706 17726 30718 17778
rect 30770 17726 30782 17778
rect 28590 17714 28642 17726
rect 7086 17666 7138 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 5842 17614 5854 17666
rect 5906 17614 5918 17666
rect 7086 17602 7138 17614
rect 7310 17666 7362 17678
rect 18510 17666 18562 17678
rect 9202 17614 9214 17666
rect 9266 17614 9278 17666
rect 13570 17614 13582 17666
rect 13634 17614 13646 17666
rect 7310 17602 7362 17614
rect 18510 17602 18562 17614
rect 18958 17666 19010 17678
rect 27694 17666 27746 17678
rect 19842 17614 19854 17666
rect 19906 17614 19918 17666
rect 23202 17614 23214 17666
rect 23266 17614 23278 17666
rect 26786 17614 26798 17666
rect 26850 17614 26862 17666
rect 18958 17602 19010 17614
rect 27694 17602 27746 17614
rect 28142 17666 28194 17678
rect 31278 17666 31330 17678
rect 30594 17614 30606 17666
rect 30658 17614 30670 17666
rect 31490 17614 31502 17666
rect 31554 17614 31566 17666
rect 28142 17602 28194 17614
rect 31278 17602 31330 17614
rect 6750 17554 6802 17566
rect 2482 17502 2494 17554
rect 2546 17502 2558 17554
rect 5618 17502 5630 17554
rect 5682 17502 5694 17554
rect 6750 17490 6802 17502
rect 7646 17554 7698 17566
rect 18174 17554 18226 17566
rect 8530 17502 8542 17554
rect 8594 17502 8606 17554
rect 12338 17502 12350 17554
rect 12402 17502 12414 17554
rect 7646 17490 7698 17502
rect 18174 17490 18226 17502
rect 18846 17554 18898 17566
rect 18846 17490 18898 17502
rect 19630 17554 19682 17566
rect 20638 17554 20690 17566
rect 19954 17502 19966 17554
rect 20018 17502 20030 17554
rect 19630 17490 19682 17502
rect 20638 17490 20690 17502
rect 21310 17554 21362 17566
rect 21310 17490 21362 17502
rect 21646 17554 21698 17566
rect 23998 17554 24050 17566
rect 22530 17502 22542 17554
rect 22594 17502 22606 17554
rect 22978 17502 22990 17554
rect 23042 17502 23054 17554
rect 21646 17490 21698 17502
rect 23998 17490 24050 17502
rect 25342 17554 25394 17566
rect 33182 17554 33234 17566
rect 25890 17502 25902 17554
rect 25954 17502 25966 17554
rect 26450 17502 26462 17554
rect 26514 17502 26526 17554
rect 25342 17490 25394 17502
rect 33182 17490 33234 17502
rect 7534 17442 7586 17454
rect 7534 17378 7586 17390
rect 8206 17442 8258 17454
rect 8206 17378 8258 17390
rect 12686 17442 12738 17454
rect 12686 17378 12738 17390
rect 17950 17442 18002 17454
rect 17950 17378 18002 17390
rect 18622 17442 18674 17454
rect 18622 17378 18674 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 19518 17442 19570 17454
rect 24222 17442 24274 17454
rect 23426 17390 23438 17442
rect 23490 17390 23502 17442
rect 19518 17378 19570 17390
rect 24222 17378 24274 17390
rect 24446 17442 24498 17454
rect 24446 17378 24498 17390
rect 24558 17442 24610 17454
rect 27022 17442 27074 17454
rect 25778 17390 25790 17442
rect 25842 17390 25854 17442
rect 24558 17378 24610 17390
rect 27022 17378 27074 17390
rect 33070 17442 33122 17454
rect 33070 17378 33122 17390
rect 1344 17274 33760 17308
rect 1344 17222 9278 17274
rect 9330 17222 9382 17274
rect 9434 17222 9486 17274
rect 9538 17222 17342 17274
rect 17394 17222 17446 17274
rect 17498 17222 17550 17274
rect 17602 17222 25406 17274
rect 25458 17222 25510 17274
rect 25562 17222 25614 17274
rect 25666 17222 33470 17274
rect 33522 17222 33574 17274
rect 33626 17222 33678 17274
rect 33730 17222 33760 17274
rect 1344 17188 33760 17222
rect 4510 17106 4562 17118
rect 4510 17042 4562 17054
rect 5182 17106 5234 17118
rect 5182 17042 5234 17054
rect 5630 17106 5682 17118
rect 5630 17042 5682 17054
rect 6638 17106 6690 17118
rect 6638 17042 6690 17054
rect 8206 17106 8258 17118
rect 8206 17042 8258 17054
rect 8766 17106 8818 17118
rect 8766 17042 8818 17054
rect 9662 17106 9714 17118
rect 9662 17042 9714 17054
rect 10894 17106 10946 17118
rect 10894 17042 10946 17054
rect 12350 17106 12402 17118
rect 24558 17106 24610 17118
rect 14242 17054 14254 17106
rect 14306 17054 14318 17106
rect 12350 17042 12402 17054
rect 24558 17042 24610 17054
rect 26574 17106 26626 17118
rect 26574 17042 26626 17054
rect 28366 17106 28418 17118
rect 28802 17054 28814 17106
rect 28866 17054 28878 17106
rect 28366 17042 28418 17054
rect 4174 16994 4226 17006
rect 4174 16930 4226 16942
rect 4398 16994 4450 17006
rect 4398 16930 4450 16942
rect 4958 16994 5010 17006
rect 4958 16930 5010 16942
rect 5294 16994 5346 17006
rect 5294 16930 5346 16942
rect 5854 16994 5906 17006
rect 5854 16930 5906 16942
rect 5966 16994 6018 17006
rect 5966 16930 6018 16942
rect 6302 16994 6354 17006
rect 6302 16930 6354 16942
rect 6414 16994 6466 17006
rect 6414 16930 6466 16942
rect 6862 16994 6914 17006
rect 6862 16930 6914 16942
rect 7870 16994 7922 17006
rect 7870 16930 7922 16942
rect 7982 16994 8034 17006
rect 11230 16994 11282 17006
rect 23886 16994 23938 17006
rect 8418 16942 8430 16994
rect 8482 16942 8494 16994
rect 20066 16942 20078 16994
rect 20130 16942 20142 16994
rect 23650 16942 23662 16994
rect 23714 16942 23726 16994
rect 7982 16930 8034 16942
rect 11230 16930 11282 16942
rect 23886 16930 23938 16942
rect 26014 16994 26066 17006
rect 26014 16930 26066 16942
rect 26126 16994 26178 17006
rect 26126 16930 26178 16942
rect 26238 16994 26290 17006
rect 26238 16930 26290 16942
rect 29374 16994 29426 17006
rect 33182 16994 33234 17006
rect 30258 16942 30270 16994
rect 30322 16942 30334 16994
rect 31266 16942 31278 16994
rect 31330 16942 31342 16994
rect 29374 16930 29426 16942
rect 33182 16930 33234 16942
rect 4846 16882 4898 16894
rect 11566 16882 11618 16894
rect 7074 16830 7086 16882
rect 7138 16830 7150 16882
rect 10658 16830 10670 16882
rect 10722 16830 10734 16882
rect 4846 16818 4898 16830
rect 11566 16818 11618 16830
rect 13918 16882 13970 16894
rect 13918 16818 13970 16830
rect 16830 16882 16882 16894
rect 27470 16882 27522 16894
rect 22754 16830 22766 16882
rect 22818 16830 22830 16882
rect 24098 16830 24110 16882
rect 24162 16830 24174 16882
rect 27346 16830 27358 16882
rect 27410 16830 27422 16882
rect 30034 16830 30046 16882
rect 30098 16830 30110 16882
rect 31154 16830 31166 16882
rect 31218 16830 31230 16882
rect 31378 16830 31390 16882
rect 31442 16830 31454 16882
rect 32050 16830 32062 16882
rect 32114 16830 32126 16882
rect 16830 16818 16882 16830
rect 27470 16818 27522 16830
rect 23550 16770 23602 16782
rect 29150 16770 29202 16782
rect 27794 16718 27806 16770
rect 27858 16718 27870 16770
rect 30258 16718 30270 16770
rect 30322 16718 30334 16770
rect 23550 16706 23602 16718
rect 29150 16706 29202 16718
rect 25554 16606 25566 16658
rect 25618 16606 25630 16658
rect 1344 16490 33600 16524
rect 1344 16438 5246 16490
rect 5298 16438 5350 16490
rect 5402 16438 5454 16490
rect 5506 16438 13310 16490
rect 13362 16438 13414 16490
rect 13466 16438 13518 16490
rect 13570 16438 21374 16490
rect 21426 16438 21478 16490
rect 21530 16438 21582 16490
rect 21634 16438 29438 16490
rect 29490 16438 29542 16490
rect 29594 16438 29646 16490
rect 29698 16438 33600 16490
rect 1344 16404 33600 16438
rect 18510 16322 18562 16334
rect 18510 16258 18562 16270
rect 19294 16322 19346 16334
rect 23538 16270 23550 16322
rect 23602 16270 23614 16322
rect 19294 16258 19346 16270
rect 7534 16210 7586 16222
rect 7534 16146 7586 16158
rect 16942 16210 16994 16222
rect 26686 16210 26738 16222
rect 31502 16210 31554 16222
rect 18722 16158 18734 16210
rect 18786 16158 18798 16210
rect 22194 16158 22206 16210
rect 22258 16158 22270 16210
rect 26002 16158 26014 16210
rect 26066 16158 26078 16210
rect 27458 16158 27470 16210
rect 27522 16158 27534 16210
rect 32610 16158 32622 16210
rect 32674 16158 32686 16210
rect 16942 16146 16994 16158
rect 26686 16146 26738 16158
rect 31502 16146 31554 16158
rect 3838 16098 3890 16110
rect 3838 16034 3890 16046
rect 4958 16098 5010 16110
rect 4958 16034 5010 16046
rect 5630 16098 5682 16110
rect 5630 16034 5682 16046
rect 5966 16098 6018 16110
rect 5966 16034 6018 16046
rect 6414 16098 6466 16110
rect 6414 16034 6466 16046
rect 10894 16098 10946 16110
rect 10894 16034 10946 16046
rect 11678 16098 11730 16110
rect 11678 16034 11730 16046
rect 16382 16098 16434 16110
rect 16382 16034 16434 16046
rect 18622 16098 18674 16110
rect 18622 16034 18674 16046
rect 19070 16098 19122 16110
rect 23886 16098 23938 16110
rect 20178 16046 20190 16098
rect 20242 16046 20254 16098
rect 20514 16046 20526 16098
rect 20578 16046 20590 16098
rect 21298 16046 21310 16098
rect 21362 16046 21374 16098
rect 22642 16046 22654 16098
rect 22706 16046 22718 16098
rect 23202 16046 23214 16098
rect 23266 16046 23278 16098
rect 19070 16034 19122 16046
rect 23886 16034 23938 16046
rect 24110 16098 24162 16110
rect 24110 16034 24162 16046
rect 24782 16098 24834 16110
rect 24782 16034 24834 16046
rect 25006 16098 25058 16110
rect 28254 16098 28306 16110
rect 30270 16098 30322 16110
rect 27010 16046 27022 16098
rect 27074 16046 27086 16098
rect 28018 16046 28030 16098
rect 28082 16046 28094 16098
rect 29362 16046 29374 16098
rect 29426 16046 29438 16098
rect 31938 16046 31950 16098
rect 32002 16046 32014 16098
rect 32946 16046 32958 16098
rect 33010 16046 33022 16098
rect 25006 16034 25058 16046
rect 28254 16034 28306 16046
rect 30270 16034 30322 16046
rect 4174 15986 4226 15998
rect 4174 15922 4226 15934
rect 4398 15986 4450 15998
rect 4398 15922 4450 15934
rect 4734 15986 4786 15998
rect 4734 15922 4786 15934
rect 6190 15986 6242 15998
rect 6190 15922 6242 15934
rect 6750 15986 6802 15998
rect 16830 15986 16882 15998
rect 11330 15934 11342 15986
rect 11394 15934 11406 15986
rect 6750 15922 6802 15934
rect 16830 15922 16882 15934
rect 17054 15986 17106 15998
rect 17838 15986 17890 15998
rect 17602 15934 17614 15986
rect 17666 15934 17678 15986
rect 17054 15922 17106 15934
rect 17838 15922 17890 15934
rect 17950 15986 18002 15998
rect 17950 15922 18002 15934
rect 21534 15986 21586 15998
rect 21534 15922 21586 15934
rect 21646 15986 21698 15998
rect 22530 15934 22542 15986
rect 22594 15934 22606 15986
rect 27682 15934 27694 15986
rect 27746 15934 27758 15986
rect 21646 15922 21698 15934
rect 28590 15930 28642 15942
rect 29138 15934 29150 15986
rect 29202 15934 29214 15986
rect 30594 15934 30606 15986
rect 30658 15934 30670 15986
rect 30818 15934 30830 15986
rect 30882 15934 30894 15986
rect 3950 15874 4002 15886
rect 3950 15810 4002 15822
rect 4510 15874 4562 15886
rect 4510 15810 4562 15822
rect 5966 15874 6018 15886
rect 5966 15810 6018 15822
rect 6638 15874 6690 15886
rect 16606 15874 16658 15886
rect 10546 15822 10558 15874
rect 10610 15822 10622 15874
rect 6638 15810 6690 15822
rect 16606 15810 16658 15822
rect 18062 15874 18114 15886
rect 18062 15810 18114 15822
rect 18174 15874 18226 15886
rect 18174 15810 18226 15822
rect 19742 15874 19794 15886
rect 19742 15810 19794 15822
rect 19854 15874 19906 15886
rect 19854 15810 19906 15822
rect 19966 15874 20018 15886
rect 25566 15874 25618 15886
rect 24434 15822 24446 15874
rect 24498 15822 24510 15874
rect 19966 15810 20018 15822
rect 25566 15810 25618 15822
rect 28478 15874 28530 15886
rect 28590 15866 28642 15878
rect 29934 15874 29986 15886
rect 28478 15810 28530 15822
rect 29934 15810 29986 15822
rect 1344 15706 33760 15740
rect 1344 15654 9278 15706
rect 9330 15654 9382 15706
rect 9434 15654 9486 15706
rect 9538 15654 17342 15706
rect 17394 15654 17446 15706
rect 17498 15654 17550 15706
rect 17602 15654 25406 15706
rect 25458 15654 25510 15706
rect 25562 15654 25614 15706
rect 25666 15654 33470 15706
rect 33522 15654 33574 15706
rect 33626 15654 33678 15706
rect 33730 15654 33760 15706
rect 1344 15620 33760 15654
rect 5070 15538 5122 15550
rect 5070 15474 5122 15486
rect 5294 15538 5346 15550
rect 5294 15474 5346 15486
rect 6750 15538 6802 15550
rect 6750 15474 6802 15486
rect 7646 15538 7698 15550
rect 7646 15474 7698 15486
rect 8206 15538 8258 15550
rect 8206 15474 8258 15486
rect 10446 15538 10498 15550
rect 10446 15474 10498 15486
rect 12350 15538 12402 15550
rect 12350 15474 12402 15486
rect 17838 15538 17890 15550
rect 17838 15474 17890 15486
rect 18510 15538 18562 15550
rect 18510 15474 18562 15486
rect 19070 15538 19122 15550
rect 19070 15474 19122 15486
rect 19294 15538 19346 15550
rect 19294 15474 19346 15486
rect 21198 15538 21250 15550
rect 21198 15474 21250 15486
rect 22878 15538 22930 15550
rect 22878 15474 22930 15486
rect 23214 15538 23266 15550
rect 28142 15538 28194 15550
rect 24658 15486 24670 15538
rect 24722 15486 24734 15538
rect 23214 15474 23266 15486
rect 28142 15474 28194 15486
rect 28254 15538 28306 15550
rect 28254 15474 28306 15486
rect 29150 15538 29202 15550
rect 29150 15474 29202 15486
rect 6414 15426 6466 15438
rect 2482 15374 2494 15426
rect 2546 15374 2558 15426
rect 6414 15362 6466 15374
rect 6974 15426 7026 15438
rect 6974 15362 7026 15374
rect 8318 15426 8370 15438
rect 8318 15362 8370 15374
rect 10222 15426 10274 15438
rect 18398 15426 18450 15438
rect 13346 15374 13358 15426
rect 13410 15374 13422 15426
rect 10222 15362 10274 15374
rect 18398 15362 18450 15374
rect 18734 15426 18786 15438
rect 18734 15362 18786 15374
rect 19406 15426 19458 15438
rect 19406 15362 19458 15374
rect 20526 15426 20578 15438
rect 20526 15362 20578 15374
rect 20750 15426 20802 15438
rect 20750 15362 20802 15374
rect 21310 15426 21362 15438
rect 23550 15426 23602 15438
rect 21634 15374 21646 15426
rect 21698 15374 21710 15426
rect 21310 15362 21362 15374
rect 23550 15362 23602 15374
rect 24110 15426 24162 15438
rect 24110 15362 24162 15374
rect 25790 15426 25842 15438
rect 25790 15362 25842 15374
rect 26910 15426 26962 15438
rect 26910 15362 26962 15374
rect 27918 15426 27970 15438
rect 27918 15362 27970 15374
rect 28702 15426 28754 15438
rect 28702 15362 28754 15374
rect 33182 15426 33234 15438
rect 33182 15362 33234 15374
rect 5406 15314 5458 15326
rect 1810 15262 1822 15314
rect 1874 15262 1886 15314
rect 5406 15250 5458 15262
rect 5854 15314 5906 15326
rect 5854 15250 5906 15262
rect 6302 15314 6354 15326
rect 6302 15250 6354 15262
rect 6638 15314 6690 15326
rect 6638 15250 6690 15262
rect 7086 15314 7138 15326
rect 7086 15250 7138 15262
rect 7534 15314 7586 15326
rect 7534 15250 7586 15262
rect 7870 15314 7922 15326
rect 7870 15250 7922 15262
rect 7982 15314 8034 15326
rect 7982 15250 8034 15262
rect 10558 15314 10610 15326
rect 10558 15250 10610 15262
rect 10670 15314 10722 15326
rect 10670 15250 10722 15262
rect 11230 15314 11282 15326
rect 18174 15314 18226 15326
rect 13122 15262 13134 15314
rect 13186 15262 13198 15314
rect 13682 15262 13694 15314
rect 13746 15262 13758 15314
rect 11230 15250 11282 15262
rect 18174 15250 18226 15262
rect 18286 15314 18338 15326
rect 18286 15250 18338 15262
rect 20078 15314 20130 15326
rect 20078 15250 20130 15262
rect 20302 15314 20354 15326
rect 20302 15250 20354 15262
rect 20862 15314 20914 15326
rect 20862 15250 20914 15262
rect 21982 15314 22034 15326
rect 24222 15314 24274 15326
rect 23874 15262 23886 15314
rect 23938 15262 23950 15314
rect 21982 15250 22034 15262
rect 24222 15250 24274 15262
rect 25678 15314 25730 15326
rect 26574 15314 26626 15326
rect 26002 15262 26014 15314
rect 26066 15262 26078 15314
rect 25678 15250 25730 15262
rect 26574 15250 26626 15262
rect 27582 15314 27634 15326
rect 28466 15262 28478 15314
rect 28530 15262 28542 15314
rect 29586 15262 29598 15314
rect 29650 15262 29662 15314
rect 27582 15250 27634 15262
rect 12014 15202 12066 15214
rect 4610 15150 4622 15202
rect 4674 15150 4686 15202
rect 12014 15138 12066 15150
rect 12238 15202 12290 15214
rect 16606 15202 16658 15214
rect 14466 15150 14478 15202
rect 14530 15150 14542 15202
rect 22418 15150 22430 15202
rect 22482 15150 22494 15202
rect 30370 15150 30382 15202
rect 30434 15150 30446 15202
rect 32498 15150 32510 15202
rect 32562 15150 32574 15202
rect 12238 15138 12290 15150
rect 16606 15138 16658 15150
rect 19730 15038 19742 15090
rect 19794 15038 19806 15090
rect 25218 15038 25230 15090
rect 25282 15038 25294 15090
rect 1344 14922 33600 14956
rect 1344 14870 5246 14922
rect 5298 14870 5350 14922
rect 5402 14870 5454 14922
rect 5506 14870 13310 14922
rect 13362 14870 13414 14922
rect 13466 14870 13518 14922
rect 13570 14870 21374 14922
rect 21426 14870 21478 14922
rect 21530 14870 21582 14922
rect 21634 14870 29438 14922
rect 29490 14870 29542 14922
rect 29594 14870 29646 14922
rect 29698 14870 33600 14922
rect 1344 14836 33600 14870
rect 17166 14754 17218 14766
rect 17166 14690 17218 14702
rect 5182 14642 5234 14654
rect 18510 14642 18562 14654
rect 29150 14642 29202 14654
rect 2482 14590 2494 14642
rect 2546 14590 2558 14642
rect 4610 14590 4622 14642
rect 4674 14590 4686 14642
rect 8978 14590 8990 14642
rect 9042 14590 9054 14642
rect 11106 14590 11118 14642
rect 11170 14590 11182 14642
rect 16370 14590 16382 14642
rect 16434 14590 16446 14642
rect 24658 14590 24670 14642
rect 24722 14590 24734 14642
rect 25666 14590 25678 14642
rect 25730 14590 25742 14642
rect 30258 14590 30270 14642
rect 30322 14590 30334 14642
rect 5182 14578 5234 14590
rect 18510 14578 18562 14590
rect 29150 14578 29202 14590
rect 6526 14530 6578 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 6526 14466 6578 14478
rect 6862 14530 6914 14542
rect 6862 14466 6914 14478
rect 7198 14530 7250 14542
rect 7198 14466 7250 14478
rect 7646 14530 7698 14542
rect 7646 14466 7698 14478
rect 7870 14530 7922 14542
rect 7870 14466 7922 14478
rect 8654 14530 8706 14542
rect 12574 14530 12626 14542
rect 18286 14530 18338 14542
rect 11890 14478 11902 14530
rect 11954 14478 11966 14530
rect 13570 14478 13582 14530
rect 13634 14478 13646 14530
rect 17938 14478 17950 14530
rect 18002 14478 18014 14530
rect 8654 14466 8706 14478
rect 12574 14466 12626 14478
rect 18286 14466 18338 14478
rect 18622 14530 18674 14542
rect 18622 14466 18674 14478
rect 18958 14530 19010 14542
rect 20066 14478 20078 14530
rect 20130 14478 20142 14530
rect 20514 14478 20526 14530
rect 20578 14478 20590 14530
rect 23426 14478 23438 14530
rect 23490 14478 23502 14530
rect 23762 14478 23774 14530
rect 23826 14478 23838 14530
rect 28578 14478 28590 14530
rect 28642 14478 28654 14530
rect 33058 14478 33070 14530
rect 33122 14478 33134 14530
rect 18958 14466 19010 14478
rect 8094 14418 8146 14430
rect 8094 14354 8146 14366
rect 8318 14418 8370 14430
rect 19518 14418 19570 14430
rect 14242 14366 14254 14418
rect 14306 14366 14318 14418
rect 17826 14366 17838 14418
rect 17890 14366 17902 14418
rect 22642 14366 22654 14418
rect 22706 14366 22718 14418
rect 23650 14366 23662 14418
rect 23714 14366 23726 14418
rect 27794 14366 27806 14418
rect 27858 14366 27870 14418
rect 32386 14366 32398 14418
rect 32450 14366 32462 14418
rect 8318 14354 8370 14366
rect 19518 14354 19570 14366
rect 6750 14306 6802 14318
rect 6750 14242 6802 14254
rect 7870 14306 7922 14318
rect 7870 14242 7922 14254
rect 8542 14306 8594 14318
rect 16830 14306 16882 14318
rect 12226 14254 12238 14306
rect 12290 14254 12302 14306
rect 8542 14242 8594 14254
rect 16830 14242 16882 14254
rect 19182 14306 19234 14318
rect 19182 14242 19234 14254
rect 19406 14306 19458 14318
rect 19406 14242 19458 14254
rect 20638 14306 20690 14318
rect 20638 14242 20690 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 29710 14306 29762 14318
rect 29710 14242 29762 14254
rect 1344 14138 33760 14172
rect 1344 14086 9278 14138
rect 9330 14086 9382 14138
rect 9434 14086 9486 14138
rect 9538 14086 17342 14138
rect 17394 14086 17446 14138
rect 17498 14086 17550 14138
rect 17602 14086 25406 14138
rect 25458 14086 25510 14138
rect 25562 14086 25614 14138
rect 25666 14086 33470 14138
rect 33522 14086 33574 14138
rect 33626 14086 33678 14138
rect 33730 14086 33760 14138
rect 1344 14052 33760 14086
rect 10558 13970 10610 13982
rect 10558 13906 10610 13918
rect 10670 13970 10722 13982
rect 10670 13906 10722 13918
rect 10782 13970 10834 13982
rect 10782 13906 10834 13918
rect 12462 13970 12514 13982
rect 12462 13906 12514 13918
rect 14142 13970 14194 13982
rect 14142 13906 14194 13918
rect 15150 13970 15202 13982
rect 15150 13906 15202 13918
rect 17838 13970 17890 13982
rect 17838 13906 17890 13918
rect 18510 13970 18562 13982
rect 23886 13970 23938 13982
rect 19282 13918 19294 13970
rect 19346 13918 19358 13970
rect 18510 13906 18562 13918
rect 20190 13914 20242 13926
rect 22866 13918 22878 13970
rect 22930 13918 22942 13970
rect 11006 13858 11058 13870
rect 6850 13806 6862 13858
rect 6914 13806 6926 13858
rect 11006 13794 11058 13806
rect 11566 13858 11618 13870
rect 11566 13794 11618 13806
rect 14478 13858 14530 13870
rect 23886 13906 23938 13918
rect 25454 13970 25506 13982
rect 25454 13906 25506 13918
rect 30046 13970 30098 13982
rect 30046 13906 30098 13918
rect 31726 13970 31778 13982
rect 32162 13918 32174 13970
rect 32226 13918 32238 13970
rect 31726 13906 31778 13918
rect 16594 13806 16606 13858
rect 16658 13806 16670 13858
rect 20190 13850 20242 13862
rect 20302 13858 20354 13870
rect 22094 13858 22146 13870
rect 23774 13858 23826 13870
rect 21074 13806 21086 13858
rect 21138 13806 21150 13858
rect 21634 13806 21646 13858
rect 21698 13806 21710 13858
rect 23090 13806 23102 13858
rect 23154 13806 23166 13858
rect 14478 13794 14530 13806
rect 20302 13794 20354 13806
rect 22094 13794 22146 13806
rect 23774 13794 23826 13806
rect 25566 13858 25618 13870
rect 25566 13794 25618 13806
rect 27918 13858 27970 13870
rect 31614 13858 31666 13870
rect 28914 13806 28926 13858
rect 28978 13806 28990 13858
rect 30594 13806 30606 13858
rect 30658 13806 30670 13858
rect 31154 13806 31166 13858
rect 31218 13806 31230 13858
rect 27918 13794 27970 13806
rect 31614 13794 31666 13806
rect 14814 13746 14866 13758
rect 17614 13746 17666 13758
rect 6178 13694 6190 13746
rect 6242 13694 6254 13746
rect 11890 13694 11902 13746
rect 11954 13694 11966 13746
rect 16706 13694 16718 13746
rect 16770 13694 16782 13746
rect 14814 13682 14866 13694
rect 17614 13682 17666 13694
rect 17726 13746 17778 13758
rect 17726 13682 17778 13694
rect 18174 13746 18226 13758
rect 18174 13682 18226 13694
rect 18398 13746 18450 13758
rect 18398 13682 18450 13694
rect 18734 13746 18786 13758
rect 18734 13682 18786 13694
rect 18958 13746 19010 13758
rect 18958 13682 19010 13694
rect 20526 13746 20578 13758
rect 23998 13746 24050 13758
rect 26574 13746 26626 13758
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 23314 13694 23326 13746
rect 23378 13694 23390 13746
rect 24322 13694 24334 13746
rect 24386 13694 24398 13746
rect 25218 13694 25230 13746
rect 25282 13694 25294 13746
rect 20526 13682 20578 13694
rect 23998 13682 24050 13694
rect 26574 13682 26626 13694
rect 26910 13746 26962 13758
rect 26910 13682 26962 13694
rect 27470 13746 27522 13758
rect 27470 13682 27522 13694
rect 28254 13746 28306 13758
rect 30382 13746 30434 13758
rect 29026 13694 29038 13746
rect 29090 13694 29102 13746
rect 28254 13682 28306 13694
rect 30382 13682 30434 13694
rect 32510 13746 32562 13758
rect 32510 13682 32562 13694
rect 10222 13634 10274 13646
rect 8978 13582 8990 13634
rect 9042 13582 9054 13634
rect 10222 13570 10274 13582
rect 11678 13634 11730 13646
rect 11678 13570 11730 13582
rect 15934 13634 15986 13646
rect 15934 13570 15986 13582
rect 19854 13634 19906 13646
rect 29598 13634 29650 13646
rect 26114 13582 26126 13634
rect 26178 13582 26190 13634
rect 19854 13570 19906 13582
rect 29598 13570 29650 13582
rect 33182 13634 33234 13646
rect 33182 13570 33234 13582
rect 15598 13522 15650 13534
rect 15598 13458 15650 13470
rect 19630 13522 19682 13534
rect 19630 13458 19682 13470
rect 22206 13522 22258 13534
rect 22206 13458 22258 13470
rect 31726 13522 31778 13534
rect 31726 13458 31778 13470
rect 1344 13354 33600 13388
rect 1344 13302 5246 13354
rect 5298 13302 5350 13354
rect 5402 13302 5454 13354
rect 5506 13302 13310 13354
rect 13362 13302 13414 13354
rect 13466 13302 13518 13354
rect 13570 13302 21374 13354
rect 21426 13302 21478 13354
rect 21530 13302 21582 13354
rect 21634 13302 29438 13354
rect 29490 13302 29542 13354
rect 29594 13302 29646 13354
rect 29698 13302 33600 13354
rect 1344 13268 33600 13302
rect 17950 13186 18002 13198
rect 22430 13186 22482 13198
rect 19058 13183 19070 13186
rect 17950 13122 18002 13134
rect 18737 13137 19070 13183
rect 18737 13074 18783 13137
rect 19058 13134 19070 13137
rect 19122 13134 19134 13186
rect 22642 13134 22654 13186
rect 22706 13183 22718 13186
rect 22978 13183 22990 13186
rect 22706 13137 22990 13183
rect 22706 13134 22718 13137
rect 22978 13134 22990 13137
rect 23042 13134 23054 13186
rect 29026 13134 29038 13186
rect 29090 13183 29102 13186
rect 29474 13183 29486 13186
rect 29090 13137 29486 13183
rect 29090 13134 29102 13137
rect 29474 13134 29486 13137
rect 29538 13134 29550 13186
rect 22430 13122 22482 13134
rect 20862 13074 20914 13086
rect 5618 13022 5630 13074
rect 5682 13022 5694 13074
rect 10770 13022 10782 13074
rect 10834 13022 10846 13074
rect 12898 13022 12910 13074
rect 12962 13022 12974 13074
rect 16370 13022 16382 13074
rect 16434 13022 16446 13074
rect 18722 13022 18734 13074
rect 18786 13022 18798 13074
rect 20862 13010 20914 13022
rect 21422 13074 21474 13086
rect 21422 13010 21474 13022
rect 21982 13074 22034 13086
rect 21982 13010 22034 13022
rect 22318 13074 22370 13086
rect 22318 13010 22370 13022
rect 23550 13074 23602 13086
rect 23550 13010 23602 13022
rect 26462 13074 26514 13086
rect 26462 13010 26514 13022
rect 28030 13074 28082 13086
rect 28030 13010 28082 13022
rect 29710 13074 29762 13086
rect 29710 13010 29762 13022
rect 30718 13074 30770 13086
rect 32386 13022 32398 13074
rect 32450 13022 32462 13074
rect 30718 13010 30770 13022
rect 17166 12962 17218 12974
rect 18622 12962 18674 12974
rect 8530 12910 8542 12962
rect 8594 12910 8606 12962
rect 9986 12910 9998 12962
rect 10050 12910 10062 12962
rect 13570 12910 13582 12962
rect 13634 12910 13646 12962
rect 18274 12910 18286 12962
rect 18338 12910 18350 12962
rect 17166 12898 17218 12910
rect 18622 12898 18674 12910
rect 19070 12962 19122 12974
rect 19070 12898 19122 12910
rect 21310 12962 21362 12974
rect 21310 12898 21362 12910
rect 23102 12962 23154 12974
rect 23102 12898 23154 12910
rect 23326 12962 23378 12974
rect 23326 12898 23378 12910
rect 23774 12962 23826 12974
rect 23774 12898 23826 12910
rect 23998 12962 24050 12974
rect 23998 12898 24050 12910
rect 24558 12962 24610 12974
rect 24558 12898 24610 12910
rect 24894 12962 24946 12974
rect 31054 12962 31106 12974
rect 25666 12910 25678 12962
rect 25730 12910 25742 12962
rect 28466 12910 28478 12962
rect 28530 12910 28542 12962
rect 30146 12910 30158 12962
rect 30210 12910 30222 12962
rect 32722 12910 32734 12962
rect 32786 12910 32798 12962
rect 24894 12898 24946 12910
rect 31054 12898 31106 12910
rect 18062 12850 18114 12862
rect 7746 12798 7758 12850
rect 7810 12798 7822 12850
rect 14242 12798 14254 12850
rect 14306 12798 14318 12850
rect 18062 12786 18114 12798
rect 25230 12850 25282 12862
rect 25230 12786 25282 12798
rect 26574 12850 26626 12862
rect 29262 12850 29314 12862
rect 26898 12798 26910 12850
rect 26962 12798 26974 12850
rect 31266 12798 31278 12850
rect 31330 12798 31342 12850
rect 31714 12798 31726 12850
rect 31778 12798 31790 12850
rect 26574 12786 26626 12798
rect 29262 12786 29314 12798
rect 25902 12738 25954 12750
rect 25902 12674 25954 12686
rect 26350 12738 26402 12750
rect 26350 12674 26402 12686
rect 27246 12738 27298 12750
rect 27246 12674 27298 12686
rect 27694 12738 27746 12750
rect 27694 12674 27746 12686
rect 1344 12570 33760 12604
rect 1344 12518 9278 12570
rect 9330 12518 9382 12570
rect 9434 12518 9486 12570
rect 9538 12518 17342 12570
rect 17394 12518 17446 12570
rect 17498 12518 17550 12570
rect 17602 12518 25406 12570
rect 25458 12518 25510 12570
rect 25562 12518 25614 12570
rect 25666 12518 33470 12570
rect 33522 12518 33574 12570
rect 33626 12518 33678 12570
rect 33730 12518 33760 12570
rect 1344 12484 33760 12518
rect 12238 12402 12290 12414
rect 12238 12338 12290 12350
rect 14590 12402 14642 12414
rect 23214 12402 23266 12414
rect 22530 12350 22542 12402
rect 22594 12350 22606 12402
rect 14590 12338 14642 12350
rect 23214 12338 23266 12350
rect 23886 12402 23938 12414
rect 23886 12338 23938 12350
rect 33070 12402 33122 12414
rect 33070 12338 33122 12350
rect 7534 12290 7586 12302
rect 13358 12290 13410 12302
rect 12562 12238 12574 12290
rect 12626 12238 12638 12290
rect 7534 12226 7586 12238
rect 13358 12226 13410 12238
rect 13694 12290 13746 12302
rect 13694 12226 13746 12238
rect 14030 12290 14082 12302
rect 14030 12226 14082 12238
rect 14926 12290 14978 12302
rect 23538 12238 23550 12290
rect 23602 12238 23614 12290
rect 24210 12238 24222 12290
rect 24274 12238 24286 12290
rect 14926 12226 14978 12238
rect 7310 12178 7362 12190
rect 7310 12114 7362 12126
rect 7646 12178 7698 12190
rect 28926 12178 28978 12190
rect 12002 12126 12014 12178
rect 12066 12126 12078 12178
rect 12786 12126 12798 12178
rect 12850 12126 12862 12178
rect 19618 12126 19630 12178
rect 19682 12126 19694 12178
rect 20178 12126 20190 12178
rect 20242 12126 20254 12178
rect 25330 12126 25342 12178
rect 25394 12126 25406 12178
rect 28578 12126 28590 12178
rect 28642 12126 28654 12178
rect 7646 12114 7698 12126
rect 28926 12114 28978 12126
rect 29150 12178 29202 12190
rect 33182 12178 33234 12190
rect 32386 12126 32398 12178
rect 32450 12126 32462 12178
rect 29150 12114 29202 12126
rect 33182 12114 33234 12126
rect 8094 12066 8146 12078
rect 8094 12002 8146 12014
rect 8542 12066 8594 12078
rect 8542 12002 8594 12014
rect 24670 12066 24722 12078
rect 29038 12066 29090 12078
rect 26114 12014 26126 12066
rect 26178 12014 26190 12066
rect 28242 12014 28254 12066
rect 28306 12014 28318 12066
rect 29586 12014 29598 12066
rect 29650 12014 29662 12066
rect 31714 12014 31726 12066
rect 31778 12014 31790 12066
rect 24670 12002 24722 12014
rect 29038 12002 29090 12014
rect 1344 11786 33600 11820
rect 1344 11734 5246 11786
rect 5298 11734 5350 11786
rect 5402 11734 5454 11786
rect 5506 11734 13310 11786
rect 13362 11734 13414 11786
rect 13466 11734 13518 11786
rect 13570 11734 21374 11786
rect 21426 11734 21478 11786
rect 21530 11734 21582 11786
rect 21634 11734 29438 11786
rect 29490 11734 29542 11786
rect 29594 11734 29646 11786
rect 29698 11734 33600 11786
rect 1344 11700 33600 11734
rect 9438 11506 9490 11518
rect 8978 11454 8990 11506
rect 9042 11454 9054 11506
rect 9438 11442 9490 11454
rect 11454 11506 11506 11518
rect 11454 11442 11506 11454
rect 12574 11506 12626 11518
rect 33182 11506 33234 11518
rect 17826 11454 17838 11506
rect 17890 11454 17902 11506
rect 19954 11454 19966 11506
rect 20018 11454 20030 11506
rect 32050 11454 32062 11506
rect 32114 11454 32126 11506
rect 12574 11442 12626 11454
rect 33182 11442 33234 11454
rect 10446 11394 10498 11406
rect 6178 11342 6190 11394
rect 6242 11342 6254 11394
rect 10446 11330 10498 11342
rect 13470 11394 13522 11406
rect 21534 11394 21586 11406
rect 17042 11342 17054 11394
rect 17106 11342 17118 11394
rect 27122 11342 27134 11394
rect 27186 11342 27198 11394
rect 29250 11342 29262 11394
rect 29314 11342 29326 11394
rect 32610 11342 32622 11394
rect 32674 11342 32686 11394
rect 13470 11330 13522 11342
rect 21534 11330 21586 11342
rect 32398 11282 32450 11294
rect 6850 11230 6862 11282
rect 6914 11230 6926 11282
rect 24994 11230 25006 11282
rect 25058 11230 25070 11282
rect 28578 11230 28590 11282
rect 28642 11230 28654 11282
rect 29922 11230 29934 11282
rect 29986 11230 29998 11282
rect 32398 11218 32450 11230
rect 9886 11170 9938 11182
rect 9886 11106 9938 11118
rect 10894 11170 10946 11182
rect 14254 11170 14306 11182
rect 13794 11118 13806 11170
rect 13858 11118 13870 11170
rect 10894 11106 10946 11118
rect 14254 11106 14306 11118
rect 14814 11170 14866 11182
rect 14814 11106 14866 11118
rect 21870 11170 21922 11182
rect 21870 11106 21922 11118
rect 22318 11170 22370 11182
rect 22318 11106 22370 11118
rect 28254 11170 28306 11182
rect 28254 11106 28306 11118
rect 1344 11002 33760 11036
rect 1344 10950 9278 11002
rect 9330 10950 9382 11002
rect 9434 10950 9486 11002
rect 9538 10950 17342 11002
rect 17394 10950 17446 11002
rect 17498 10950 17550 11002
rect 17602 10950 25406 11002
rect 25458 10950 25510 11002
rect 25562 10950 25614 11002
rect 25666 10950 33470 11002
rect 33522 10950 33574 11002
rect 33626 10950 33678 11002
rect 33730 10950 33760 11002
rect 1344 10916 33760 10950
rect 4510 10834 4562 10846
rect 4510 10770 4562 10782
rect 5406 10834 5458 10846
rect 5406 10770 5458 10782
rect 5966 10834 6018 10846
rect 5966 10770 6018 10782
rect 6414 10834 6466 10846
rect 6414 10770 6466 10782
rect 6862 10834 6914 10846
rect 6862 10770 6914 10782
rect 7758 10834 7810 10846
rect 7758 10770 7810 10782
rect 7870 10834 7922 10846
rect 7870 10770 7922 10782
rect 8654 10834 8706 10846
rect 8654 10770 8706 10782
rect 11566 10834 11618 10846
rect 11566 10770 11618 10782
rect 19742 10834 19794 10846
rect 19742 10770 19794 10782
rect 20190 10834 20242 10846
rect 20190 10770 20242 10782
rect 21310 10834 21362 10846
rect 21310 10770 21362 10782
rect 26238 10834 26290 10846
rect 26238 10770 26290 10782
rect 33182 10834 33234 10846
rect 33182 10770 33234 10782
rect 3614 10722 3666 10734
rect 3614 10658 3666 10670
rect 6750 10722 6802 10734
rect 6750 10658 6802 10670
rect 7310 10722 7362 10734
rect 7310 10658 7362 10670
rect 9662 10722 9714 10734
rect 9662 10658 9714 10670
rect 11006 10722 11058 10734
rect 25678 10722 25730 10734
rect 11890 10670 11902 10722
rect 11954 10670 11966 10722
rect 19394 10670 19406 10722
rect 19458 10670 19470 10722
rect 20962 10670 20974 10722
rect 21026 10670 21038 10722
rect 11006 10658 11058 10670
rect 25678 10658 25730 10670
rect 26462 10722 26514 10734
rect 26462 10658 26514 10670
rect 3390 10610 3442 10622
rect 3390 10546 3442 10558
rect 3726 10610 3778 10622
rect 3726 10546 3778 10558
rect 5518 10610 5570 10622
rect 5518 10546 5570 10558
rect 6974 10610 7026 10622
rect 6974 10546 7026 10558
rect 7646 10610 7698 10622
rect 10558 10610 10610 10622
rect 8194 10558 8206 10610
rect 8258 10558 8270 10610
rect 7646 10546 7698 10558
rect 10558 10546 10610 10558
rect 11230 10610 11282 10622
rect 15598 10610 15650 10622
rect 12226 10558 12238 10610
rect 12290 10558 12302 10610
rect 11230 10546 11282 10558
rect 15598 10546 15650 10558
rect 15710 10610 15762 10622
rect 15710 10546 15762 10558
rect 16158 10610 16210 10622
rect 16158 10546 16210 10558
rect 17278 10610 17330 10622
rect 17278 10546 17330 10558
rect 17614 10610 17666 10622
rect 17614 10546 17666 10558
rect 17838 10610 17890 10622
rect 17838 10546 17890 10558
rect 19966 10610 20018 10622
rect 19966 10546 20018 10558
rect 20302 10610 20354 10622
rect 20302 10546 20354 10558
rect 20526 10610 20578 10622
rect 25230 10610 25282 10622
rect 21858 10558 21870 10610
rect 21922 10558 21934 10610
rect 20526 10546 20578 10558
rect 25230 10546 25282 10558
rect 25454 10610 25506 10622
rect 25454 10546 25506 10558
rect 26126 10610 26178 10622
rect 26126 10546 26178 10558
rect 26686 10610 26738 10622
rect 27122 10558 27134 10610
rect 27186 10558 27198 10610
rect 26686 10546 26738 10558
rect 4846 10498 4898 10510
rect 4846 10434 4898 10446
rect 10446 10498 10498 10510
rect 10446 10434 10498 10446
rect 10782 10498 10834 10510
rect 15934 10498 15986 10510
rect 13010 10446 13022 10498
rect 13074 10446 13086 10498
rect 15138 10446 15150 10498
rect 15202 10446 15214 10498
rect 10782 10434 10834 10446
rect 15934 10434 15986 10446
rect 17502 10498 17554 10510
rect 25342 10498 25394 10510
rect 22530 10446 22542 10498
rect 22594 10446 22606 10498
rect 24658 10446 24670 10498
rect 24722 10446 24734 10498
rect 31714 10446 31726 10498
rect 31778 10446 31790 10498
rect 17502 10434 17554 10446
rect 25342 10434 25394 10446
rect 5406 10386 5458 10398
rect 5730 10334 5742 10386
rect 5794 10383 5806 10386
rect 6514 10383 6526 10386
rect 5794 10337 6526 10383
rect 5794 10334 5806 10337
rect 6514 10334 6526 10337
rect 6578 10334 6590 10386
rect 5406 10322 5458 10334
rect 1344 10218 33600 10252
rect 1344 10166 5246 10218
rect 5298 10166 5350 10218
rect 5402 10166 5454 10218
rect 5506 10166 13310 10218
rect 13362 10166 13414 10218
rect 13466 10166 13518 10218
rect 13570 10166 21374 10218
rect 21426 10166 21478 10218
rect 21530 10166 21582 10218
rect 21634 10166 29438 10218
rect 29490 10166 29542 10218
rect 29594 10166 29646 10218
rect 29698 10166 33600 10218
rect 1344 10132 33600 10166
rect 8766 10050 8818 10062
rect 8766 9986 8818 9998
rect 5070 9938 5122 9950
rect 12574 9938 12626 9950
rect 9986 9886 9998 9938
rect 10050 9886 10062 9938
rect 12114 9886 12126 9938
rect 12178 9886 12190 9938
rect 5070 9874 5122 9886
rect 12574 9874 12626 9886
rect 13918 9938 13970 9950
rect 13918 9874 13970 9886
rect 15150 9938 15202 9950
rect 15150 9874 15202 9886
rect 15710 9938 15762 9950
rect 20078 9938 20130 9950
rect 17266 9886 17278 9938
rect 17330 9886 17342 9938
rect 19394 9886 19406 9938
rect 19458 9886 19470 9938
rect 15710 9874 15762 9886
rect 20078 9874 20130 9886
rect 22206 9938 22258 9950
rect 22206 9874 22258 9886
rect 23438 9938 23490 9950
rect 23438 9874 23490 9886
rect 26238 9938 26290 9950
rect 26238 9874 26290 9886
rect 27134 9938 27186 9950
rect 27134 9874 27186 9886
rect 28366 9938 28418 9950
rect 30258 9886 30270 9938
rect 30322 9886 30334 9938
rect 28366 9874 28418 9886
rect 2830 9826 2882 9838
rect 2830 9762 2882 9774
rect 3166 9826 3218 9838
rect 3166 9762 3218 9774
rect 3390 9826 3442 9838
rect 3390 9762 3442 9774
rect 3726 9826 3778 9838
rect 3726 9762 3778 9774
rect 4174 9826 4226 9838
rect 4174 9762 4226 9774
rect 4734 9826 4786 9838
rect 4734 9762 4786 9774
rect 5742 9826 5794 9838
rect 5742 9762 5794 9774
rect 6414 9826 6466 9838
rect 6414 9762 6466 9774
rect 7086 9826 7138 9838
rect 14142 9826 14194 9838
rect 9202 9774 9214 9826
rect 9266 9774 9278 9826
rect 7086 9762 7138 9774
rect 14142 9762 14194 9774
rect 14366 9826 14418 9838
rect 14366 9762 14418 9774
rect 16270 9826 16322 9838
rect 19966 9826 20018 9838
rect 16594 9774 16606 9826
rect 16658 9774 16670 9826
rect 16270 9762 16322 9774
rect 19966 9762 20018 9774
rect 20638 9826 20690 9838
rect 20638 9762 20690 9774
rect 22542 9826 22594 9838
rect 22542 9762 22594 9774
rect 23550 9826 23602 9838
rect 23550 9762 23602 9774
rect 23886 9826 23938 9838
rect 23886 9762 23938 9774
rect 24446 9826 24498 9838
rect 25454 9826 25506 9838
rect 24770 9774 24782 9826
rect 24834 9774 24846 9826
rect 24446 9762 24498 9774
rect 25454 9762 25506 9774
rect 26350 9826 26402 9838
rect 26350 9762 26402 9774
rect 26798 9826 26850 9838
rect 26798 9762 26850 9774
rect 27022 9826 27074 9838
rect 27022 9762 27074 9774
rect 27246 9826 27298 9838
rect 27246 9762 27298 9774
rect 28030 9826 28082 9838
rect 28030 9762 28082 9774
rect 28142 9826 28194 9838
rect 28142 9762 28194 9774
rect 28590 9826 28642 9838
rect 28590 9762 28642 9774
rect 29150 9826 29202 9838
rect 33058 9774 33070 9826
rect 33122 9774 33134 9826
rect 29150 9762 29202 9774
rect 7422 9714 7474 9726
rect 6738 9662 6750 9714
rect 6802 9662 6814 9714
rect 7422 9650 7474 9662
rect 7646 9714 7698 9726
rect 8654 9714 8706 9726
rect 8306 9662 8318 9714
rect 8370 9662 8382 9714
rect 7646 9650 7698 9662
rect 8654 9650 8706 9662
rect 13806 9714 13858 9726
rect 13806 9650 13858 9662
rect 20190 9714 20242 9726
rect 20190 9650 20242 9662
rect 23326 9714 23378 9726
rect 23326 9650 23378 9662
rect 24334 9714 24386 9726
rect 24334 9650 24386 9662
rect 25230 9714 25282 9726
rect 25230 9650 25282 9662
rect 25790 9714 25842 9726
rect 25790 9650 25842 9662
rect 29262 9714 29314 9726
rect 32386 9662 32398 9714
rect 32450 9662 32462 9714
rect 29262 9650 29314 9662
rect 2494 9602 2546 9614
rect 2494 9538 2546 9550
rect 2718 9602 2770 9614
rect 2718 9538 2770 9550
rect 3390 9602 3442 9614
rect 3390 9538 3442 9550
rect 4062 9602 4114 9614
rect 4062 9538 4114 9550
rect 4286 9602 4338 9614
rect 7310 9602 7362 9614
rect 6066 9550 6078 9602
rect 6130 9550 6142 9602
rect 4286 9538 4338 9550
rect 7310 9538 7362 9550
rect 7982 9602 8034 9614
rect 7982 9538 8034 9550
rect 8766 9602 8818 9614
rect 8766 9538 8818 9550
rect 14814 9602 14866 9614
rect 14814 9538 14866 9550
rect 15038 9602 15090 9614
rect 15038 9538 15090 9550
rect 15262 9602 15314 9614
rect 15262 9538 15314 9550
rect 15598 9602 15650 9614
rect 15598 9538 15650 9550
rect 15822 9602 15874 9614
rect 24222 9602 24274 9614
rect 22866 9550 22878 9602
rect 22930 9550 22942 9602
rect 15822 9538 15874 9550
rect 24222 9538 24274 9550
rect 25678 9602 25730 9614
rect 25678 9538 25730 9550
rect 26126 9602 26178 9614
rect 26126 9538 26178 9550
rect 27470 9602 27522 9614
rect 27470 9538 27522 9550
rect 29374 9602 29426 9614
rect 29374 9538 29426 9550
rect 29598 9602 29650 9614
rect 29598 9538 29650 9550
rect 1344 9434 33760 9468
rect 1344 9382 9278 9434
rect 9330 9382 9382 9434
rect 9434 9382 9486 9434
rect 9538 9382 17342 9434
rect 17394 9382 17446 9434
rect 17498 9382 17550 9434
rect 17602 9382 25406 9434
rect 25458 9382 25510 9434
rect 25562 9382 25614 9434
rect 25666 9382 33470 9434
rect 33522 9382 33574 9434
rect 33626 9382 33678 9434
rect 33730 9382 33760 9434
rect 1344 9348 33760 9382
rect 4958 9266 5010 9278
rect 4958 9202 5010 9214
rect 9662 9266 9714 9278
rect 11454 9266 11506 9278
rect 10658 9214 10670 9266
rect 10722 9214 10734 9266
rect 9662 9202 9714 9214
rect 11454 9202 11506 9214
rect 13134 9266 13186 9278
rect 13134 9202 13186 9214
rect 17502 9266 17554 9278
rect 17502 9202 17554 9214
rect 17838 9266 17890 9278
rect 17838 9202 17890 9214
rect 17950 9266 18002 9278
rect 17950 9202 18002 9214
rect 18174 9266 18226 9278
rect 18174 9202 18226 9214
rect 22318 9266 22370 9278
rect 22318 9202 22370 9214
rect 25566 9266 25618 9278
rect 25566 9202 25618 9214
rect 29262 9266 29314 9278
rect 29262 9202 29314 9214
rect 29374 9266 29426 9278
rect 31278 9266 31330 9278
rect 30258 9214 30270 9266
rect 30322 9214 30334 9266
rect 29374 9202 29426 9214
rect 31278 9202 31330 9214
rect 31390 9266 31442 9278
rect 31390 9202 31442 9214
rect 32286 9266 32338 9278
rect 32286 9202 32338 9214
rect 33294 9266 33346 9278
rect 33294 9202 33346 9214
rect 10222 9154 10274 9166
rect 3826 9102 3838 9154
rect 3890 9102 3902 9154
rect 8082 9102 8094 9154
rect 8146 9102 8158 9154
rect 10222 9090 10274 9102
rect 12350 9154 12402 9166
rect 18398 9154 18450 9166
rect 23550 9154 23602 9166
rect 29150 9154 29202 9166
rect 14466 9102 14478 9154
rect 14530 9102 14542 9154
rect 19730 9102 19742 9154
rect 19794 9102 19806 9154
rect 24546 9102 24558 9154
rect 24610 9102 24622 9154
rect 25218 9102 25230 9154
rect 25282 9102 25294 9154
rect 26674 9102 26686 9154
rect 26738 9102 26750 9154
rect 12350 9090 12402 9102
rect 18398 9090 18450 9102
rect 23550 9090 23602 9102
rect 29150 9090 29202 9102
rect 31838 9154 31890 9166
rect 31838 9090 31890 9102
rect 5182 9042 5234 9054
rect 9774 9042 9826 9054
rect 4610 8990 4622 9042
rect 4674 8990 4686 9042
rect 5506 8990 5518 9042
rect 5570 8990 5582 9042
rect 8866 8990 8878 9042
rect 8930 8990 8942 9042
rect 5182 8978 5234 8990
rect 9774 8978 9826 8990
rect 10110 9042 10162 9054
rect 10110 8978 10162 8990
rect 10446 9042 10498 9054
rect 11342 9042 11394 9054
rect 10882 8990 10894 9042
rect 10946 8990 10958 9042
rect 10446 8978 10498 8990
rect 11342 8978 11394 8990
rect 11566 9042 11618 9054
rect 12126 9042 12178 9054
rect 11890 8990 11902 9042
rect 11954 8990 11966 9042
rect 11566 8978 11618 8990
rect 12126 8978 12178 8990
rect 12462 9042 12514 9054
rect 17726 9042 17778 9054
rect 13682 8990 13694 9042
rect 13746 8990 13758 9042
rect 12462 8978 12514 8990
rect 17726 8978 17778 8990
rect 18510 9042 18562 9054
rect 29822 9042 29874 9054
rect 19058 8990 19070 9042
rect 19122 8990 19134 9042
rect 23762 8990 23774 9042
rect 23826 8990 23838 9042
rect 24322 8990 24334 9042
rect 24386 8990 24398 9042
rect 26002 8990 26014 9042
rect 26066 8990 26078 9042
rect 18510 8978 18562 8990
rect 29822 8978 29874 8990
rect 30606 9042 30658 9054
rect 31502 9042 31554 9054
rect 30930 8990 30942 9042
rect 30994 8990 31006 9042
rect 30606 8978 30658 8990
rect 31502 8978 31554 8990
rect 32062 9042 32114 9054
rect 32062 8978 32114 8990
rect 32398 9042 32450 9054
rect 32398 8978 32450 8990
rect 5070 8930 5122 8942
rect 22878 8930 22930 8942
rect 1698 8878 1710 8930
rect 1762 8878 1774 8930
rect 5954 8878 5966 8930
rect 6018 8878 6030 8930
rect 16594 8878 16606 8930
rect 16658 8878 16670 8930
rect 21858 8878 21870 8930
rect 21922 8878 21934 8930
rect 5070 8866 5122 8878
rect 22878 8866 22930 8878
rect 23214 8930 23266 8942
rect 28802 8878 28814 8930
rect 28866 8878 28878 8930
rect 23214 8866 23266 8878
rect 9662 8818 9714 8830
rect 9662 8754 9714 8766
rect 1344 8650 33600 8684
rect 1344 8598 5246 8650
rect 5298 8598 5350 8650
rect 5402 8598 5454 8650
rect 5506 8598 13310 8650
rect 13362 8598 13414 8650
rect 13466 8598 13518 8650
rect 13570 8598 21374 8650
rect 21426 8598 21478 8650
rect 21530 8598 21582 8650
rect 21634 8598 29438 8650
rect 29490 8598 29542 8650
rect 29594 8598 29646 8650
rect 29698 8598 33600 8650
rect 1344 8564 33600 8598
rect 24782 8482 24834 8494
rect 21970 8430 21982 8482
rect 22034 8479 22046 8482
rect 22754 8479 22766 8482
rect 22034 8433 22766 8479
rect 22034 8430 22046 8433
rect 22754 8430 22766 8433
rect 22818 8430 22830 8482
rect 24782 8418 24834 8430
rect 5854 8370 5906 8382
rect 22318 8370 22370 8382
rect 4610 8318 4622 8370
rect 4674 8318 4686 8370
rect 8866 8318 8878 8370
rect 8930 8318 8942 8370
rect 5854 8306 5906 8318
rect 22318 8306 22370 8318
rect 25342 8370 25394 8382
rect 25342 8306 25394 8318
rect 30046 8370 30098 8382
rect 30258 8318 30270 8370
rect 30322 8318 30334 8370
rect 30046 8306 30098 8318
rect 5966 8258 6018 8270
rect 12574 8258 12626 8270
rect 19630 8258 19682 8270
rect 1810 8206 1822 8258
rect 1874 8206 1886 8258
rect 11666 8206 11678 8258
rect 11730 8206 11742 8258
rect 14914 8206 14926 8258
rect 14978 8206 14990 8258
rect 5966 8194 6018 8206
rect 12574 8194 12626 8206
rect 19630 8194 19682 8206
rect 23214 8258 23266 8270
rect 23214 8194 23266 8206
rect 23774 8258 23826 8270
rect 23774 8194 23826 8206
rect 24334 8258 24386 8270
rect 24334 8194 24386 8206
rect 26238 8258 26290 8270
rect 26238 8194 26290 8206
rect 28030 8258 28082 8270
rect 28030 8194 28082 8206
rect 28142 8258 28194 8270
rect 28142 8194 28194 8206
rect 28254 8258 28306 8270
rect 28254 8194 28306 8206
rect 28702 8258 28754 8270
rect 33058 8206 33070 8258
rect 33122 8206 33134 8258
rect 28702 8194 28754 8206
rect 5742 8146 5794 8158
rect 2482 8094 2494 8146
rect 2546 8094 2558 8146
rect 5742 8082 5794 8094
rect 6302 8146 6354 8158
rect 21870 8146 21922 8158
rect 17826 8094 17838 8146
rect 17890 8094 17902 8146
rect 20290 8094 20302 8146
rect 20354 8094 20366 8146
rect 6302 8082 6354 8094
rect 21870 8082 21922 8094
rect 24670 8146 24722 8158
rect 24670 8082 24722 8094
rect 27246 8146 27298 8158
rect 27246 8082 27298 8094
rect 27694 8146 27746 8158
rect 29474 8094 29486 8146
rect 29538 8094 29550 8146
rect 32386 8094 32398 8146
rect 32450 8094 32462 8146
rect 27694 8082 27746 8094
rect 5182 8034 5234 8046
rect 19406 8034 19458 8046
rect 12898 7982 12910 8034
rect 12962 7982 12974 8034
rect 5182 7970 5234 7982
rect 19406 7970 19458 7982
rect 19518 8034 19570 8046
rect 19518 7970 19570 7982
rect 19854 8034 19906 8046
rect 19854 7970 19906 7982
rect 20638 8034 20690 8046
rect 20638 7970 20690 7982
rect 22766 8034 22818 8046
rect 22766 7970 22818 7982
rect 22878 8034 22930 8046
rect 22878 7970 22930 7982
rect 23102 8034 23154 8046
rect 23102 7970 23154 7982
rect 23438 8034 23490 8046
rect 23438 7970 23490 7982
rect 23662 8034 23714 8046
rect 23662 7970 23714 7982
rect 23998 8034 24050 8046
rect 23998 7970 24050 7982
rect 24222 8034 24274 8046
rect 24222 7970 24274 7982
rect 24782 8034 24834 8046
rect 24782 7970 24834 7982
rect 25902 8034 25954 8046
rect 25902 7970 25954 7982
rect 26798 8034 26850 8046
rect 26798 7970 26850 7982
rect 27358 8034 27410 8046
rect 27358 7970 27410 7982
rect 27582 8034 27634 8046
rect 27582 7970 27634 7982
rect 29150 8034 29202 8046
rect 29150 7970 29202 7982
rect 1344 7866 33760 7900
rect 1344 7814 9278 7866
rect 9330 7814 9382 7866
rect 9434 7814 9486 7866
rect 9538 7814 17342 7866
rect 17394 7814 17446 7866
rect 17498 7814 17550 7866
rect 17602 7814 25406 7866
rect 25458 7814 25510 7866
rect 25562 7814 25614 7866
rect 25666 7814 33470 7866
rect 33522 7814 33574 7866
rect 33626 7814 33678 7866
rect 33730 7814 33760 7866
rect 1344 7780 33760 7814
rect 3054 7698 3106 7710
rect 3054 7634 3106 7646
rect 4174 7698 4226 7710
rect 4174 7634 4226 7646
rect 4398 7698 4450 7710
rect 4398 7634 4450 7646
rect 5854 7698 5906 7710
rect 5854 7634 5906 7646
rect 7758 7698 7810 7710
rect 7758 7634 7810 7646
rect 7870 7698 7922 7710
rect 7870 7634 7922 7646
rect 13246 7698 13298 7710
rect 13246 7634 13298 7646
rect 17502 7698 17554 7710
rect 17502 7634 17554 7646
rect 17614 7698 17666 7710
rect 17614 7634 17666 7646
rect 19854 7698 19906 7710
rect 19854 7634 19906 7646
rect 20302 7698 20354 7710
rect 20302 7634 20354 7646
rect 21646 7698 21698 7710
rect 21646 7634 21698 7646
rect 23326 7698 23378 7710
rect 23326 7634 23378 7646
rect 24670 7698 24722 7710
rect 24670 7634 24722 7646
rect 27470 7698 27522 7710
rect 27470 7634 27522 7646
rect 28366 7698 28418 7710
rect 28366 7634 28418 7646
rect 29598 7698 29650 7710
rect 29598 7634 29650 7646
rect 30046 7698 30098 7710
rect 30046 7634 30098 7646
rect 31054 7698 31106 7710
rect 31054 7634 31106 7646
rect 32062 7698 32114 7710
rect 32062 7634 32114 7646
rect 33182 7698 33234 7710
rect 33182 7634 33234 7646
rect 2494 7586 2546 7598
rect 2494 7522 2546 7534
rect 3278 7586 3330 7598
rect 3278 7522 3330 7534
rect 3502 7586 3554 7598
rect 3502 7522 3554 7534
rect 4958 7586 5010 7598
rect 4958 7522 5010 7534
rect 5966 7586 6018 7598
rect 16718 7586 16770 7598
rect 8530 7534 8542 7586
rect 8594 7534 8606 7586
rect 5966 7522 6018 7534
rect 16718 7522 16770 7534
rect 19294 7586 19346 7598
rect 19294 7522 19346 7534
rect 21758 7586 21810 7598
rect 21758 7522 21810 7534
rect 22094 7586 22146 7598
rect 28590 7586 28642 7598
rect 29374 7586 29426 7598
rect 25554 7534 25566 7586
rect 25618 7534 25630 7586
rect 26674 7534 26686 7586
rect 26738 7534 26750 7586
rect 27794 7534 27806 7586
rect 27858 7534 27870 7586
rect 28914 7534 28926 7586
rect 28978 7534 28990 7586
rect 22094 7522 22146 7534
rect 28590 7522 28642 7534
rect 29374 7522 29426 7534
rect 30382 7586 30434 7598
rect 30382 7522 30434 7534
rect 2382 7474 2434 7486
rect 2034 7422 2046 7474
rect 2098 7422 2110 7474
rect 2382 7410 2434 7422
rect 2606 7474 2658 7486
rect 2606 7410 2658 7422
rect 2830 7474 2882 7486
rect 4286 7474 4338 7486
rect 3826 7422 3838 7474
rect 3890 7422 3902 7474
rect 2830 7410 2882 7422
rect 4286 7410 4338 7422
rect 4846 7474 4898 7486
rect 4846 7410 4898 7422
rect 5406 7474 5458 7486
rect 5406 7410 5458 7422
rect 5630 7474 5682 7486
rect 5630 7410 5682 7422
rect 6078 7474 6130 7486
rect 6078 7410 6130 7422
rect 6750 7474 6802 7486
rect 6750 7410 6802 7422
rect 6974 7474 7026 7486
rect 6974 7410 7026 7422
rect 7422 7474 7474 7486
rect 7422 7410 7474 7422
rect 7646 7474 7698 7486
rect 13134 7474 13186 7486
rect 16606 7474 16658 7486
rect 8194 7422 8206 7474
rect 8258 7422 8270 7474
rect 8754 7422 8766 7474
rect 8818 7422 8830 7474
rect 12338 7422 12350 7474
rect 12402 7422 12414 7474
rect 13682 7422 13694 7474
rect 13746 7422 13758 7474
rect 7646 7410 7698 7422
rect 13134 7410 13186 7422
rect 16606 7410 16658 7422
rect 16942 7474 16994 7486
rect 16942 7410 16994 7422
rect 17390 7474 17442 7486
rect 17390 7410 17442 7422
rect 18062 7474 18114 7486
rect 18062 7410 18114 7422
rect 18286 7474 18338 7486
rect 18286 7410 18338 7422
rect 18622 7474 18674 7486
rect 18622 7410 18674 7422
rect 18846 7474 18898 7486
rect 18846 7410 18898 7422
rect 19406 7474 19458 7486
rect 19406 7410 19458 7422
rect 22318 7474 22370 7486
rect 22318 7410 22370 7422
rect 22766 7474 22818 7486
rect 22766 7410 22818 7422
rect 23102 7474 23154 7486
rect 23102 7410 23154 7422
rect 23438 7474 23490 7486
rect 23438 7410 23490 7422
rect 25230 7474 25282 7486
rect 25230 7410 25282 7422
rect 27022 7474 27074 7486
rect 27022 7410 27074 7422
rect 29262 7474 29314 7486
rect 29262 7410 29314 7422
rect 30606 7474 30658 7486
rect 30606 7410 30658 7422
rect 31278 7474 31330 7486
rect 31278 7410 31330 7422
rect 31614 7474 31666 7486
rect 31614 7410 31666 7422
rect 31950 7474 32002 7486
rect 31950 7410 32002 7422
rect 32174 7474 32226 7486
rect 32174 7410 32226 7422
rect 5182 7362 5234 7374
rect 5182 7298 5234 7310
rect 6862 7362 6914 7374
rect 18734 7362 18786 7374
rect 9538 7310 9550 7362
rect 9602 7310 9614 7362
rect 11666 7310 11678 7362
rect 11730 7310 11742 7362
rect 14914 7310 14926 7362
rect 14978 7310 14990 7362
rect 6862 7298 6914 7310
rect 18734 7298 18786 7310
rect 21310 7362 21362 7374
rect 21310 7298 21362 7310
rect 22206 7362 22258 7374
rect 22206 7298 22258 7310
rect 24334 7362 24386 7374
rect 24334 7298 24386 7310
rect 26462 7362 26514 7374
rect 26462 7298 26514 7310
rect 31166 7362 31218 7374
rect 31166 7298 31218 7310
rect 13246 7250 13298 7262
rect 13246 7186 13298 7198
rect 19294 7250 19346 7262
rect 19294 7186 19346 7198
rect 21646 7250 21698 7262
rect 21646 7186 21698 7198
rect 1344 7082 33600 7116
rect 1344 7030 5246 7082
rect 5298 7030 5350 7082
rect 5402 7030 5454 7082
rect 5506 7030 13310 7082
rect 13362 7030 13414 7082
rect 13466 7030 13518 7082
rect 13570 7030 21374 7082
rect 21426 7030 21478 7082
rect 21530 7030 21582 7082
rect 21634 7030 29438 7082
rect 29490 7030 29542 7082
rect 29594 7030 29646 7082
rect 29698 7030 33600 7082
rect 1344 6996 33600 7030
rect 10894 6802 10946 6814
rect 16942 6802 16994 6814
rect 23550 6802 23602 6814
rect 16482 6750 16494 6802
rect 16546 6750 16558 6802
rect 20738 6750 20750 6802
rect 20802 6750 20814 6802
rect 10894 6738 10946 6750
rect 16942 6738 16994 6750
rect 23550 6738 23602 6750
rect 31502 6802 31554 6814
rect 31502 6738 31554 6750
rect 10670 6690 10722 6702
rect 4050 6638 4062 6690
rect 4114 6638 4126 6690
rect 4834 6638 4846 6690
rect 4898 6638 4910 6690
rect 5842 6638 5854 6690
rect 5906 6638 5918 6690
rect 9650 6638 9662 6690
rect 9714 6638 9726 6690
rect 10670 6626 10722 6638
rect 11342 6690 11394 6702
rect 11342 6626 11394 6638
rect 11902 6690 11954 6702
rect 11902 6626 11954 6638
rect 12462 6690 12514 6702
rect 12462 6626 12514 6638
rect 12910 6690 12962 6702
rect 17054 6690 17106 6702
rect 21646 6690 21698 6702
rect 13570 6638 13582 6690
rect 13634 6638 13646 6690
rect 17826 6638 17838 6690
rect 17890 6638 17902 6690
rect 12910 6626 12962 6638
rect 17054 6626 17106 6638
rect 21646 6626 21698 6638
rect 22430 6690 22482 6702
rect 22430 6626 22482 6638
rect 22766 6690 22818 6702
rect 22766 6626 22818 6638
rect 23102 6690 23154 6702
rect 23102 6626 23154 6638
rect 24110 6690 24162 6702
rect 24110 6626 24162 6638
rect 24558 6690 24610 6702
rect 24558 6626 24610 6638
rect 25678 6690 25730 6702
rect 25678 6626 25730 6638
rect 26350 6690 26402 6702
rect 26350 6626 26402 6638
rect 27134 6690 27186 6702
rect 27134 6626 27186 6638
rect 28366 6690 28418 6702
rect 28366 6626 28418 6638
rect 28702 6690 28754 6702
rect 28702 6626 28754 6638
rect 30046 6690 30098 6702
rect 30046 6626 30098 6638
rect 30606 6690 30658 6702
rect 30606 6626 30658 6638
rect 30718 6690 30770 6702
rect 30718 6626 30770 6638
rect 31390 6690 31442 6702
rect 31390 6626 31442 6638
rect 32510 6690 32562 6702
rect 32510 6626 32562 6638
rect 33182 6690 33234 6702
rect 33182 6626 33234 6638
rect 10222 6578 10274 6590
rect 9426 6526 9438 6578
rect 9490 6526 9502 6578
rect 10222 6514 10274 6526
rect 10334 6578 10386 6590
rect 10334 6514 10386 6526
rect 11118 6578 11170 6590
rect 11118 6514 11170 6526
rect 11790 6578 11842 6590
rect 11790 6514 11842 6526
rect 12798 6578 12850 6590
rect 21982 6578 22034 6590
rect 14354 6526 14366 6578
rect 14418 6526 14430 6578
rect 18610 6526 18622 6578
rect 18674 6526 18686 6578
rect 12798 6514 12850 6526
rect 21982 6514 22034 6526
rect 22206 6578 22258 6590
rect 22206 6514 22258 6526
rect 24446 6578 24498 6590
rect 27470 6578 27522 6590
rect 26786 6526 26798 6578
rect 26850 6526 26862 6578
rect 24446 6514 24498 6526
rect 27470 6514 27522 6526
rect 27806 6578 27858 6590
rect 27806 6514 27858 6526
rect 29486 6578 29538 6590
rect 29486 6514 29538 6526
rect 29822 6578 29874 6590
rect 29822 6514 29874 6526
rect 31614 6578 31666 6590
rect 31614 6514 31666 6526
rect 32174 6578 32226 6590
rect 32174 6514 32226 6526
rect 32846 6578 32898 6590
rect 32846 6514 32898 6526
rect 3278 6466 3330 6478
rect 6862 6466 6914 6478
rect 9102 6466 9154 6478
rect 5058 6414 5070 6466
rect 5122 6414 5134 6466
rect 8754 6414 8766 6466
rect 8818 6414 8830 6466
rect 3278 6402 3330 6414
rect 6862 6402 6914 6414
rect 9102 6402 9154 6414
rect 10558 6466 10610 6478
rect 10558 6402 10610 6414
rect 11566 6466 11618 6478
rect 11566 6402 11618 6414
rect 12574 6466 12626 6478
rect 12574 6402 12626 6414
rect 16830 6466 16882 6478
rect 16830 6402 16882 6414
rect 17278 6466 17330 6478
rect 17278 6402 17330 6414
rect 21758 6466 21810 6478
rect 21758 6402 21810 6414
rect 22654 6466 22706 6478
rect 22654 6402 22706 6414
rect 23438 6466 23490 6478
rect 23438 6402 23490 6414
rect 23662 6466 23714 6478
rect 23662 6402 23714 6414
rect 24222 6466 24274 6478
rect 24222 6402 24274 6414
rect 25118 6466 25170 6478
rect 28478 6466 28530 6478
rect 25330 6414 25342 6466
rect 25394 6414 25406 6466
rect 26002 6414 26014 6466
rect 26066 6414 26078 6466
rect 25118 6402 25170 6414
rect 28478 6402 28530 6414
rect 30494 6466 30546 6478
rect 30494 6402 30546 6414
rect 31166 6466 31218 6478
rect 31166 6402 31218 6414
rect 1344 6298 33760 6332
rect 1344 6246 9278 6298
rect 9330 6246 9382 6298
rect 9434 6246 9486 6298
rect 9538 6246 17342 6298
rect 17394 6246 17446 6298
rect 17498 6246 17550 6298
rect 17602 6246 25406 6298
rect 25458 6246 25510 6298
rect 25562 6246 25614 6298
rect 25666 6246 33470 6298
rect 33522 6246 33574 6298
rect 33626 6246 33678 6298
rect 33730 6246 33760 6298
rect 1344 6212 33760 6246
rect 5294 6130 5346 6142
rect 5294 6066 5346 6078
rect 22206 6130 22258 6142
rect 22206 6066 22258 6078
rect 22318 6130 22370 6142
rect 22318 6066 22370 6078
rect 22430 6130 22482 6142
rect 22430 6066 22482 6078
rect 23550 6130 23602 6142
rect 23550 6066 23602 6078
rect 24110 6130 24162 6142
rect 24110 6066 24162 6078
rect 26126 6130 26178 6142
rect 26126 6066 26178 6078
rect 27358 6130 27410 6142
rect 27358 6066 27410 6078
rect 28254 6130 28306 6142
rect 28254 6066 28306 6078
rect 29150 6130 29202 6142
rect 29150 6066 29202 6078
rect 29374 6130 29426 6142
rect 29374 6066 29426 6078
rect 29598 6130 29650 6142
rect 29598 6066 29650 6078
rect 31726 6130 31778 6142
rect 31726 6066 31778 6078
rect 31950 6130 32002 6142
rect 31950 6066 32002 6078
rect 33070 6130 33122 6142
rect 33070 6066 33122 6078
rect 5070 6018 5122 6030
rect 9662 6018 9714 6030
rect 3826 5966 3838 6018
rect 3890 5966 3902 6018
rect 8082 5966 8094 6018
rect 8146 5966 8158 6018
rect 5070 5954 5122 5966
rect 9662 5954 9714 5966
rect 9774 6018 9826 6030
rect 9774 5954 9826 5966
rect 10446 6018 10498 6030
rect 10446 5954 10498 5966
rect 10782 6018 10834 6030
rect 10782 5954 10834 5966
rect 11006 6018 11058 6030
rect 11006 5954 11058 5966
rect 17726 6018 17778 6030
rect 17726 5954 17778 5966
rect 17950 6018 18002 6030
rect 24558 6018 24610 6030
rect 19730 5966 19742 6018
rect 19794 5966 19806 6018
rect 17950 5954 18002 5966
rect 24558 5954 24610 5966
rect 25566 6018 25618 6030
rect 25566 5954 25618 5966
rect 27246 6018 27298 6030
rect 27246 5954 27298 5966
rect 27918 6018 27970 6030
rect 27918 5954 27970 5966
rect 28030 6018 28082 6030
rect 28030 5954 28082 5966
rect 28478 6018 28530 6030
rect 28478 5954 28530 5966
rect 28590 6018 28642 6030
rect 28590 5954 28642 5966
rect 29038 6018 29090 6030
rect 29038 5954 29090 5966
rect 29822 6018 29874 6030
rect 29822 5954 29874 5966
rect 31054 6018 31106 6030
rect 31054 5954 31106 5966
rect 5406 5906 5458 5918
rect 4498 5854 4510 5906
rect 4562 5854 4574 5906
rect 5406 5842 5458 5854
rect 5518 5906 5570 5918
rect 17278 5906 17330 5918
rect 8866 5854 8878 5906
rect 8930 5854 8942 5906
rect 11778 5854 11790 5906
rect 11842 5854 11854 5906
rect 14242 5854 14254 5906
rect 14306 5854 14318 5906
rect 5518 5842 5570 5854
rect 17278 5842 17330 5854
rect 17502 5906 17554 5918
rect 23102 5906 23154 5918
rect 19058 5854 19070 5906
rect 19122 5854 19134 5906
rect 22754 5854 22766 5906
rect 22818 5854 22830 5906
rect 17502 5842 17554 5854
rect 23102 5842 23154 5854
rect 23326 5906 23378 5918
rect 23326 5842 23378 5854
rect 24334 5906 24386 5918
rect 24334 5842 24386 5854
rect 25230 5906 25282 5918
rect 25230 5842 25282 5854
rect 25342 5906 25394 5918
rect 25342 5842 25394 5854
rect 25790 5906 25842 5918
rect 25790 5842 25842 5854
rect 26238 5906 26290 5918
rect 26238 5842 26290 5854
rect 26350 5906 26402 5918
rect 27582 5906 27634 5918
rect 26674 5854 26686 5906
rect 26738 5854 26750 5906
rect 26350 5842 26402 5854
rect 27582 5842 27634 5854
rect 28814 5906 28866 5918
rect 30382 5906 30434 5918
rect 30146 5854 30158 5906
rect 30210 5854 30222 5906
rect 28814 5842 28866 5854
rect 30382 5842 30434 5854
rect 30830 5906 30882 5918
rect 30830 5842 30882 5854
rect 31278 5906 31330 5918
rect 31278 5842 31330 5854
rect 10558 5794 10610 5806
rect 1698 5742 1710 5794
rect 1762 5742 1774 5794
rect 5954 5742 5966 5794
rect 6018 5742 6030 5794
rect 10558 5730 10610 5742
rect 18398 5794 18450 5806
rect 23214 5794 23266 5806
rect 21858 5742 21870 5794
rect 21922 5742 21934 5794
rect 18398 5730 18450 5742
rect 23214 5730 23266 5742
rect 24446 5794 24498 5806
rect 24446 5730 24498 5742
rect 29710 5794 29762 5806
rect 29710 5730 29762 5742
rect 30942 5794 30994 5806
rect 30942 5730 30994 5742
rect 31838 5794 31890 5806
rect 31838 5730 31890 5742
rect 32398 5794 32450 5806
rect 32398 5730 32450 5742
rect 33182 5794 33234 5806
rect 33182 5730 33234 5742
rect 9774 5682 9826 5694
rect 9774 5618 9826 5630
rect 12350 5682 12402 5694
rect 12350 5618 12402 5630
rect 15262 5682 15314 5694
rect 15262 5618 15314 5630
rect 32286 5682 32338 5694
rect 32286 5618 32338 5630
rect 1344 5514 33600 5548
rect 1344 5462 5246 5514
rect 5298 5462 5350 5514
rect 5402 5462 5454 5514
rect 5506 5462 13310 5514
rect 13362 5462 13414 5514
rect 13466 5462 13518 5514
rect 13570 5462 21374 5514
rect 21426 5462 21478 5514
rect 21530 5462 21582 5514
rect 21634 5462 29438 5514
rect 29490 5462 29542 5514
rect 29594 5462 29646 5514
rect 29698 5462 33600 5514
rect 1344 5428 33600 5462
rect 26798 5346 26850 5358
rect 26798 5282 26850 5294
rect 2718 5234 2770 5246
rect 20302 5234 20354 5246
rect 9762 5182 9774 5234
rect 9826 5182 9838 5234
rect 11890 5182 11902 5234
rect 11954 5182 11966 5234
rect 18722 5182 18734 5234
rect 18786 5182 18798 5234
rect 2718 5170 2770 5182
rect 20302 5170 20354 5182
rect 20750 5234 20802 5246
rect 20750 5170 20802 5182
rect 22542 5234 22594 5246
rect 22542 5170 22594 5182
rect 24558 5234 24610 5246
rect 24558 5170 24610 5182
rect 25454 5234 25506 5246
rect 25454 5170 25506 5182
rect 28478 5234 28530 5246
rect 30258 5182 30270 5234
rect 30322 5182 30334 5234
rect 28478 5170 28530 5182
rect 2270 5122 2322 5134
rect 5854 5122 5906 5134
rect 12126 5122 12178 5134
rect 4610 5070 4622 5122
rect 4674 5070 4686 5122
rect 8418 5070 8430 5122
rect 8482 5070 8494 5122
rect 8978 5070 8990 5122
rect 9042 5070 9054 5122
rect 2270 5058 2322 5070
rect 5854 5058 5906 5070
rect 12126 5058 12178 5070
rect 12350 5122 12402 5134
rect 12350 5058 12402 5070
rect 12574 5122 12626 5134
rect 12574 5058 12626 5070
rect 12798 5122 12850 5134
rect 12798 5058 12850 5070
rect 13918 5122 13970 5134
rect 13918 5058 13970 5070
rect 14142 5122 14194 5134
rect 14142 5058 14194 5070
rect 14478 5122 14530 5134
rect 14478 5058 14530 5070
rect 14814 5122 14866 5134
rect 18958 5122 19010 5134
rect 15362 5070 15374 5122
rect 15426 5070 15438 5122
rect 15810 5070 15822 5122
rect 15874 5070 15886 5122
rect 14814 5058 14866 5070
rect 18958 5058 19010 5070
rect 19966 5122 20018 5134
rect 24334 5122 24386 5134
rect 21522 5070 21534 5122
rect 21586 5070 21598 5122
rect 19966 5058 20018 5070
rect 24334 5058 24386 5070
rect 24782 5122 24834 5134
rect 24782 5058 24834 5070
rect 24894 5122 24946 5134
rect 24894 5058 24946 5070
rect 25342 5122 25394 5134
rect 25342 5058 25394 5070
rect 26014 5122 26066 5134
rect 26014 5058 26066 5070
rect 26126 5122 26178 5134
rect 26126 5058 26178 5070
rect 26462 5122 26514 5134
rect 28030 5122 28082 5134
rect 27570 5070 27582 5122
rect 27634 5070 27646 5122
rect 26462 5058 26514 5070
rect 28030 5058 28082 5070
rect 28142 5122 28194 5134
rect 28142 5058 28194 5070
rect 29038 5122 29090 5134
rect 29038 5058 29090 5070
rect 29374 5122 29426 5134
rect 29374 5058 29426 5070
rect 29710 5122 29762 5134
rect 32386 5070 32398 5122
rect 32450 5070 32462 5122
rect 33058 5070 33070 5122
rect 33122 5070 33134 5122
rect 29710 5058 29762 5070
rect 1934 5010 1986 5022
rect 1934 4946 1986 4958
rect 2046 5010 2098 5022
rect 15150 5010 15202 5022
rect 19294 5010 19346 5022
rect 7074 4958 7086 5010
rect 7138 4958 7150 5010
rect 13570 4958 13582 5010
rect 13634 4958 13646 5010
rect 16594 4958 16606 5010
rect 16658 4958 16670 5010
rect 2046 4946 2098 4958
rect 15150 4946 15202 4958
rect 19294 4946 19346 4958
rect 19630 5010 19682 5022
rect 19630 4946 19682 4958
rect 26350 5010 26402 5022
rect 26350 4946 26402 4958
rect 26910 5010 26962 5022
rect 26910 4946 26962 4958
rect 27918 5010 27970 5022
rect 27918 4946 27970 4958
rect 28590 5010 28642 5022
rect 28590 4946 28642 4958
rect 14478 4898 14530 4910
rect 14478 4834 14530 4846
rect 19182 4898 19234 4910
rect 19182 4834 19234 4846
rect 19742 4898 19794 4910
rect 19742 4834 19794 4846
rect 25566 4898 25618 4910
rect 25566 4834 25618 4846
rect 29262 4898 29314 4910
rect 29262 4834 29314 4846
rect 1344 4730 33760 4764
rect 1344 4678 9278 4730
rect 9330 4678 9382 4730
rect 9434 4678 9486 4730
rect 9538 4678 17342 4730
rect 17394 4678 17446 4730
rect 17498 4678 17550 4730
rect 17602 4678 25406 4730
rect 25458 4678 25510 4730
rect 25562 4678 25614 4730
rect 25666 4678 33470 4730
rect 33522 4678 33574 4730
rect 33626 4678 33678 4730
rect 33730 4678 33760 4730
rect 1344 4644 33760 4678
rect 8206 4562 8258 4574
rect 8206 4498 8258 4510
rect 8318 4562 8370 4574
rect 8318 4498 8370 4510
rect 16606 4562 16658 4574
rect 16606 4498 16658 4510
rect 24110 4562 24162 4574
rect 24110 4498 24162 4510
rect 31838 4562 31890 4574
rect 31838 4498 31890 4510
rect 33070 4562 33122 4574
rect 33070 4498 33122 4510
rect 24558 4450 24610 4462
rect 32062 4450 32114 4462
rect 3826 4398 3838 4450
rect 3890 4398 3902 4450
rect 5730 4398 5742 4450
rect 5794 4398 5806 4450
rect 14802 4398 14814 4450
rect 14866 4398 14878 4450
rect 18162 4398 18174 4450
rect 18226 4398 18238 4450
rect 21634 4398 21646 4450
rect 21698 4398 21710 4450
rect 26002 4398 26014 4450
rect 26066 4398 26078 4450
rect 29250 4398 29262 4450
rect 29314 4398 29326 4450
rect 24558 4386 24610 4398
rect 32062 4386 32114 4398
rect 8430 4338 8482 4350
rect 16382 4338 16434 4350
rect 4498 4286 4510 4338
rect 4562 4286 4574 4338
rect 4946 4286 4958 4338
rect 5010 4286 5022 4338
rect 8754 4286 8766 4338
rect 8818 4286 8830 4338
rect 12002 4286 12014 4338
rect 12066 4286 12078 4338
rect 15586 4286 15598 4338
rect 15650 4286 15662 4338
rect 8430 4274 8482 4286
rect 16382 4274 16434 4286
rect 16606 4338 16658 4350
rect 16606 4274 16658 4286
rect 16942 4338 16994 4350
rect 31614 4338 31666 4350
rect 17378 4286 17390 4338
rect 17442 4286 17454 4338
rect 20850 4286 20862 4338
rect 20914 4286 20926 4338
rect 25330 4286 25342 4338
rect 25394 4286 25406 4338
rect 28578 4286 28590 4338
rect 28642 4286 28654 4338
rect 16942 4274 16994 4286
rect 31614 4274 31666 4286
rect 32174 4338 32226 4350
rect 32174 4274 32226 4286
rect 24222 4226 24274 4238
rect 1698 4174 1710 4226
rect 1762 4174 1774 4226
rect 7858 4174 7870 4226
rect 7922 4174 7934 4226
rect 10322 4174 10334 4226
rect 10386 4174 10398 4226
rect 12674 4174 12686 4226
rect 12738 4174 12750 4226
rect 20290 4174 20302 4226
rect 20354 4174 20366 4226
rect 23762 4174 23774 4226
rect 23826 4174 23838 4226
rect 24222 4162 24274 4174
rect 24670 4226 24722 4238
rect 33182 4226 33234 4238
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 31378 4174 31390 4226
rect 31442 4174 31454 4226
rect 24670 4162 24722 4174
rect 33182 4162 33234 4174
rect 1344 3946 33600 3980
rect 1344 3894 5246 3946
rect 5298 3894 5350 3946
rect 5402 3894 5454 3946
rect 5506 3894 13310 3946
rect 13362 3894 13414 3946
rect 13466 3894 13518 3946
rect 13570 3894 21374 3946
rect 21426 3894 21478 3946
rect 21530 3894 21582 3946
rect 21634 3894 29438 3946
rect 29490 3894 29542 3946
rect 29594 3894 29646 3946
rect 29698 3894 33600 3946
rect 1344 3860 33600 3894
rect 26898 3726 26910 3778
rect 26962 3775 26974 3778
rect 27906 3775 27918 3778
rect 26962 3729 27918 3775
rect 26962 3726 26974 3729
rect 27906 3726 27918 3729
rect 27970 3726 27982 3778
rect 8542 3666 8594 3678
rect 16158 3666 16210 3678
rect 25566 3666 25618 3678
rect 9538 3614 9550 3666
rect 9602 3614 9614 3666
rect 11666 3614 11678 3666
rect 11730 3614 11742 3666
rect 18162 3614 18174 3666
rect 18226 3614 18238 3666
rect 21858 3614 21870 3666
rect 21922 3614 21934 3666
rect 8542 3602 8594 3614
rect 16158 3602 16210 3614
rect 25566 3602 25618 3614
rect 13246 3554 13298 3566
rect 2370 3502 2382 3554
rect 2434 3502 2446 3554
rect 6178 3502 6190 3554
rect 6242 3502 6254 3554
rect 12450 3502 12462 3554
rect 12514 3502 12526 3554
rect 13246 3490 13298 3502
rect 13582 3554 13634 3566
rect 16942 3554 16994 3566
rect 13794 3502 13806 3554
rect 13858 3502 13870 3554
rect 13582 3490 13634 3502
rect 16942 3490 16994 3502
rect 17278 3554 17330 3566
rect 27022 3554 27074 3566
rect 30270 3554 30322 3566
rect 33182 3554 33234 3566
rect 20066 3502 20078 3554
rect 20130 3502 20142 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 24882 3502 24894 3554
rect 24946 3502 24958 3554
rect 26450 3502 26462 3554
rect 26514 3502 26526 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 29586 3502 29598 3554
rect 29650 3502 29662 3554
rect 32274 3502 32286 3554
rect 32338 3502 32350 3554
rect 17278 3490 17330 3502
rect 27022 3490 27074 3502
rect 30270 3490 30322 3502
rect 33182 3490 33234 3502
rect 1822 3442 1874 3454
rect 5742 3442 5794 3454
rect 4050 3390 4062 3442
rect 4114 3390 4126 3442
rect 13358 3442 13410 3454
rect 1822 3378 1874 3390
rect 5742 3378 5794 3390
rect 5854 3386 5906 3398
rect 1934 3330 1986 3342
rect 1934 3266 1986 3278
rect 2158 3330 2210 3342
rect 2158 3266 2210 3278
rect 5518 3330 5570 3342
rect 13358 3378 13410 3390
rect 17166 3442 17218 3454
rect 17166 3378 17218 3390
rect 23662 3442 23714 3454
rect 23662 3378 23714 3390
rect 23998 3442 24050 3454
rect 23998 3378 24050 3390
rect 24670 3442 24722 3454
rect 24670 3378 24722 3390
rect 25902 3442 25954 3454
rect 25902 3378 25954 3390
rect 26238 3442 26290 3454
rect 26238 3378 26290 3390
rect 27470 3442 27522 3454
rect 27470 3378 27522 3390
rect 28366 3442 28418 3454
rect 28366 3378 28418 3390
rect 29374 3442 29426 3454
rect 29374 3378 29426 3390
rect 30606 3442 30658 3454
rect 30606 3378 30658 3390
rect 30942 3442 30994 3454
rect 30942 3378 30994 3390
rect 31278 3442 31330 3454
rect 31278 3378 31330 3390
rect 32510 3442 32562 3454
rect 32510 3378 32562 3390
rect 32846 3442 32898 3454
rect 32846 3378 32898 3390
rect 5854 3322 5906 3334
rect 5518 3266 5570 3278
rect 1344 3162 33760 3196
rect 1344 3110 9278 3162
rect 9330 3110 9382 3162
rect 9434 3110 9486 3162
rect 9538 3110 17342 3162
rect 17394 3110 17446 3162
rect 17498 3110 17550 3162
rect 17602 3110 25406 3162
rect 25458 3110 25510 3162
rect 25562 3110 25614 3162
rect 25666 3110 33470 3162
rect 33522 3110 33574 3162
rect 33626 3110 33678 3162
rect 33730 3110 33760 3162
rect 1344 3076 33760 3110
<< via1 >>
rect 478 31502 530 31554
rect 2270 31502 2322 31554
rect 9278 31334 9330 31386
rect 9382 31334 9434 31386
rect 9486 31334 9538 31386
rect 17342 31334 17394 31386
rect 17446 31334 17498 31386
rect 17550 31334 17602 31386
rect 25406 31334 25458 31386
rect 25510 31334 25562 31386
rect 25614 31334 25666 31386
rect 33470 31334 33522 31386
rect 33574 31334 33626 31386
rect 33678 31334 33730 31386
rect 1822 31166 1874 31218
rect 2270 31166 2322 31218
rect 2942 31166 2994 31218
rect 3950 31166 4002 31218
rect 4510 31166 4562 31218
rect 4958 31166 5010 31218
rect 5854 31166 5906 31218
rect 18622 31166 18674 31218
rect 21758 31166 21810 31218
rect 24558 31166 24610 31218
rect 26238 31166 26290 31218
rect 3726 31054 3778 31106
rect 7982 31054 8034 31106
rect 16942 31054 16994 31106
rect 23662 31054 23714 31106
rect 24894 31054 24946 31106
rect 29150 31054 29202 31106
rect 6638 30942 6690 30994
rect 9438 30942 9490 30994
rect 13806 30942 13858 30994
rect 17278 30942 17330 30994
rect 17950 30942 18002 30994
rect 20750 30942 20802 30994
rect 23886 30942 23938 30994
rect 25342 30942 25394 30994
rect 28366 30942 28418 30994
rect 32286 30942 32338 30994
rect 32734 30942 32786 30994
rect 10110 30830 10162 30882
rect 12238 30830 12290 30882
rect 13358 30830 13410 30882
rect 16158 30830 16210 30882
rect 31278 30830 31330 30882
rect 32174 30830 32226 30882
rect 13470 30718 13522 30770
rect 32286 30718 32338 30770
rect 32958 30718 33010 30770
rect 5246 30550 5298 30602
rect 5350 30550 5402 30602
rect 5454 30550 5506 30602
rect 13310 30550 13362 30602
rect 13414 30550 13466 30602
rect 13518 30550 13570 30602
rect 21374 30550 21426 30602
rect 21478 30550 21530 30602
rect 21582 30550 21634 30602
rect 29438 30550 29490 30602
rect 29542 30550 29594 30602
rect 29646 30550 29698 30602
rect 5070 30270 5122 30322
rect 8542 30270 8594 30322
rect 18622 30270 18674 30322
rect 20638 30270 20690 30322
rect 27694 30270 27746 30322
rect 32510 30270 32562 30322
rect 2270 30158 2322 30210
rect 5630 30158 5682 30210
rect 9774 30158 9826 30210
rect 13806 30158 13858 30210
rect 14814 30158 14866 30210
rect 14926 30158 14978 30210
rect 15710 30158 15762 30210
rect 16494 30158 16546 30210
rect 19070 30158 19122 30210
rect 19630 30158 19682 30210
rect 21310 30158 21362 30210
rect 24894 30158 24946 30210
rect 29262 30158 29314 30210
rect 29598 30158 29650 30210
rect 33070 30158 33122 30210
rect 2942 30046 2994 30098
rect 6414 30046 6466 30098
rect 9326 30046 9378 30098
rect 10558 30046 10610 30098
rect 15038 30046 15090 30098
rect 20302 30046 20354 30098
rect 20414 30046 20466 30098
rect 22094 30046 22146 30098
rect 25566 30046 25618 30098
rect 30382 30046 30434 30098
rect 32846 30046 32898 30098
rect 8878 29934 8930 29986
rect 9438 29934 9490 29986
rect 12798 29934 12850 29986
rect 14030 29934 14082 29986
rect 14366 29934 14418 29986
rect 20526 29934 20578 29986
rect 20750 29934 20802 29986
rect 24334 29934 24386 29986
rect 28030 29934 28082 29986
rect 28366 29934 28418 29986
rect 9278 29766 9330 29818
rect 9382 29766 9434 29818
rect 9486 29766 9538 29818
rect 17342 29766 17394 29818
rect 17446 29766 17498 29818
rect 17550 29766 17602 29818
rect 25406 29766 25458 29818
rect 25510 29766 25562 29818
rect 25614 29766 25666 29818
rect 33470 29766 33522 29818
rect 33574 29766 33626 29818
rect 33678 29766 33730 29818
rect 3950 29598 4002 29650
rect 5070 29598 5122 29650
rect 5518 29598 5570 29650
rect 7198 29598 7250 29650
rect 9102 29598 9154 29650
rect 10110 29598 10162 29650
rect 11678 29598 11730 29650
rect 18398 29598 18450 29650
rect 22318 29598 22370 29650
rect 22542 29598 22594 29650
rect 6078 29486 6130 29538
rect 7422 29486 7474 29538
rect 8206 29486 8258 29538
rect 8542 29486 8594 29538
rect 10222 29486 10274 29538
rect 11342 29486 11394 29538
rect 12798 29486 12850 29538
rect 15934 29486 15986 29538
rect 22990 29486 23042 29538
rect 23102 29486 23154 29538
rect 30606 29486 30658 29538
rect 5854 29374 5906 29426
rect 7758 29374 7810 29426
rect 8654 29374 8706 29426
rect 12126 29374 12178 29426
rect 15710 29374 15762 29426
rect 15822 29374 15874 29426
rect 16158 29374 16210 29426
rect 17726 29374 17778 29426
rect 18174 29374 18226 29426
rect 18846 29374 18898 29426
rect 22206 29374 22258 29426
rect 22766 29374 22818 29426
rect 22878 29374 22930 29426
rect 23438 29374 23490 29426
rect 24110 29374 24162 29426
rect 24446 29374 24498 29426
rect 25454 29374 25506 29426
rect 26126 29374 26178 29426
rect 26574 29374 26626 29426
rect 31950 29374 32002 29426
rect 4062 29262 4114 29314
rect 4510 29262 4562 29314
rect 6750 29262 6802 29314
rect 8094 29262 8146 29314
rect 9662 29262 9714 29314
rect 10894 29262 10946 29314
rect 14926 29262 14978 29314
rect 17390 29262 17442 29314
rect 18286 29262 18338 29314
rect 19518 29262 19570 29314
rect 21758 29262 21810 29314
rect 23886 29262 23938 29314
rect 27358 29262 27410 29314
rect 29486 29262 29538 29314
rect 33182 29262 33234 29314
rect 9998 29150 10050 29202
rect 11006 29150 11058 29202
rect 16606 29150 16658 29202
rect 17502 29150 17554 29202
rect 25678 29150 25730 29202
rect 26126 29150 26178 29202
rect 26238 29150 26290 29202
rect 5246 28982 5298 29034
rect 5350 28982 5402 29034
rect 5454 28982 5506 29034
rect 13310 28982 13362 29034
rect 13414 28982 13466 29034
rect 13518 28982 13570 29034
rect 21374 28982 21426 29034
rect 21478 28982 21530 29034
rect 21582 28982 21634 29034
rect 29438 28982 29490 29034
rect 29542 28982 29594 29034
rect 29646 28982 29698 29034
rect 8430 28814 8482 28866
rect 9326 28814 9378 28866
rect 9662 28814 9714 28866
rect 11342 28814 11394 28866
rect 18734 28814 18786 28866
rect 26910 28814 26962 28866
rect 4622 28702 4674 28754
rect 6078 28702 6130 28754
rect 7646 28702 7698 28754
rect 8430 28702 8482 28754
rect 9326 28702 9378 28754
rect 13470 28702 13522 28754
rect 18286 28702 18338 28754
rect 21870 28702 21922 28754
rect 23438 28702 23490 28754
rect 25566 28702 25618 28754
rect 29934 28702 29986 28754
rect 31054 28702 31106 28754
rect 33182 28702 33234 28754
rect 1710 28590 1762 28642
rect 5182 28590 5234 28642
rect 6414 28590 6466 28642
rect 7870 28590 7922 28642
rect 10334 28590 10386 28642
rect 14142 28590 14194 28642
rect 14478 28590 14530 28642
rect 15038 28590 15090 28642
rect 15486 28590 15538 28642
rect 19294 28590 19346 28642
rect 19966 28590 20018 28642
rect 20302 28590 20354 28642
rect 22206 28590 22258 28642
rect 22654 28590 22706 28642
rect 25902 28590 25954 28642
rect 30270 28590 30322 28642
rect 2494 28478 2546 28530
rect 6302 28478 6354 28530
rect 6638 28478 6690 28530
rect 7534 28478 7586 28530
rect 9998 28478 10050 28530
rect 13694 28478 13746 28530
rect 13806 28478 13858 28530
rect 14702 28478 14754 28530
rect 16158 28478 16210 28530
rect 18734 28478 18786 28530
rect 18846 28478 18898 28530
rect 20638 28478 20690 28530
rect 21534 28478 21586 28530
rect 21870 28478 21922 28530
rect 29374 28478 29426 28530
rect 29486 28478 29538 28530
rect 29598 28478 29650 28530
rect 5742 28366 5794 28418
rect 6862 28366 6914 28418
rect 8990 28366 9042 28418
rect 9774 28366 9826 28418
rect 19182 28366 19234 28418
rect 19406 28366 19458 28418
rect 19630 28366 19682 28418
rect 20190 28366 20242 28418
rect 21758 28366 21810 28418
rect 29150 28366 29202 28418
rect 9278 28198 9330 28250
rect 9382 28198 9434 28250
rect 9486 28198 9538 28250
rect 17342 28198 17394 28250
rect 17446 28198 17498 28250
rect 17550 28198 17602 28250
rect 25406 28198 25458 28250
rect 25510 28198 25562 28250
rect 25614 28198 25666 28250
rect 33470 28198 33522 28250
rect 33574 28198 33626 28250
rect 33678 28198 33730 28250
rect 5070 28030 5122 28082
rect 5518 28030 5570 28082
rect 8094 28030 8146 28082
rect 12238 28030 12290 28082
rect 15150 28030 15202 28082
rect 18510 28030 18562 28082
rect 20526 28030 20578 28082
rect 24334 28030 24386 28082
rect 24558 28030 24610 28082
rect 25790 28030 25842 28082
rect 26126 28030 26178 28082
rect 26238 28030 26290 28082
rect 26350 28030 26402 28082
rect 7758 27918 7810 27970
rect 9662 27918 9714 27970
rect 9886 27918 9938 27970
rect 10782 27918 10834 27970
rect 24670 27918 24722 27970
rect 26462 27918 26514 27970
rect 30270 27918 30322 27970
rect 1710 27806 1762 27858
rect 6302 27806 6354 27858
rect 7198 27806 7250 27858
rect 9774 27806 9826 27858
rect 10670 27806 10722 27858
rect 11230 27806 11282 27858
rect 14142 27806 14194 27858
rect 17726 27806 17778 27858
rect 20414 27806 20466 27858
rect 20974 27806 21026 27858
rect 25454 27806 25506 27858
rect 26910 27806 26962 27858
rect 27246 27806 27298 27858
rect 2494 27694 2546 27746
rect 4622 27694 4674 27746
rect 6750 27694 6802 27746
rect 8542 27694 8594 27746
rect 9102 27694 9154 27746
rect 21758 27694 21810 27746
rect 23998 27694 24050 27746
rect 25230 27694 25282 27746
rect 33182 27694 33234 27746
rect 7310 27582 7362 27634
rect 7534 27582 7586 27634
rect 10334 27582 10386 27634
rect 10782 27582 10834 27634
rect 20526 27582 20578 27634
rect 5246 27414 5298 27466
rect 5350 27414 5402 27466
rect 5454 27414 5506 27466
rect 13310 27414 13362 27466
rect 13414 27414 13466 27466
rect 13518 27414 13570 27466
rect 21374 27414 21426 27466
rect 21478 27414 21530 27466
rect 21582 27414 21634 27466
rect 29438 27414 29490 27466
rect 29542 27414 29594 27466
rect 29646 27414 29698 27466
rect 2830 27246 2882 27298
rect 3278 27246 3330 27298
rect 12574 27246 12626 27298
rect 12910 27246 12962 27298
rect 14142 27246 14194 27298
rect 18734 27246 18786 27298
rect 28478 27246 28530 27298
rect 2942 27134 2994 27186
rect 6302 27134 6354 27186
rect 6750 27134 6802 27186
rect 7982 27134 8034 27186
rect 9214 27134 9266 27186
rect 9998 27134 10050 27186
rect 10670 27134 10722 27186
rect 12350 27134 12402 27186
rect 16830 27134 16882 27186
rect 22318 27134 22370 27186
rect 26014 27134 26066 27186
rect 28142 27134 28194 27186
rect 28590 27134 28642 27186
rect 31054 27134 31106 27186
rect 33182 27134 33234 27186
rect 4846 27022 4898 27074
rect 7534 27022 7586 27074
rect 8542 27022 8594 27074
rect 9550 27022 9602 27074
rect 10222 27022 10274 27074
rect 10782 27022 10834 27074
rect 11790 27022 11842 27074
rect 14478 27022 14530 27074
rect 14590 27022 14642 27074
rect 15710 27022 15762 27074
rect 18734 27022 18786 27074
rect 19294 27022 19346 27074
rect 19966 27022 20018 27074
rect 20526 27022 20578 27074
rect 24110 27022 24162 27074
rect 25342 27022 25394 27074
rect 29598 27022 29650 27074
rect 29934 27022 29986 27074
rect 30270 27022 30322 27074
rect 3390 26910 3442 26962
rect 5182 26910 5234 26962
rect 5966 26910 6018 26962
rect 6078 26910 6130 26962
rect 6190 26910 6242 26962
rect 6974 26910 7026 26962
rect 7198 26910 7250 26962
rect 8094 26910 8146 26962
rect 8206 26910 8258 26962
rect 10670 26910 10722 26962
rect 11006 26910 11058 26962
rect 11230 26910 11282 26962
rect 11902 26910 11954 26962
rect 13470 26910 13522 26962
rect 14814 26910 14866 26962
rect 18174 26910 18226 26962
rect 18398 26910 18450 26962
rect 20638 26910 20690 26962
rect 21310 26910 21362 26962
rect 29262 26910 29314 26962
rect 29374 26910 29426 26962
rect 4958 26798 5010 26850
rect 6414 26798 6466 26850
rect 7310 26798 7362 26850
rect 7870 26798 7922 26850
rect 9774 26798 9826 26850
rect 9998 26798 10050 26850
rect 12126 26798 12178 26850
rect 13806 26798 13858 26850
rect 14702 26798 14754 26850
rect 18958 26798 19010 26850
rect 19406 26798 19458 26850
rect 21646 26798 21698 26850
rect 29150 26798 29202 26850
rect 9278 26630 9330 26682
rect 9382 26630 9434 26682
rect 9486 26630 9538 26682
rect 17342 26630 17394 26682
rect 17446 26630 17498 26682
rect 17550 26630 17602 26682
rect 25406 26630 25458 26682
rect 25510 26630 25562 26682
rect 25614 26630 25666 26682
rect 33470 26630 33522 26682
rect 33574 26630 33626 26682
rect 33678 26630 33730 26682
rect 7758 26462 7810 26514
rect 12462 26462 12514 26514
rect 12574 26462 12626 26514
rect 14030 26462 14082 26514
rect 16270 26462 16322 26514
rect 17726 26462 17778 26514
rect 18398 26462 18450 26514
rect 18622 26462 18674 26514
rect 19966 26462 20018 26514
rect 6526 26350 6578 26402
rect 7422 26350 7474 26402
rect 8542 26350 8594 26402
rect 9774 26350 9826 26402
rect 11118 26350 11170 26402
rect 15934 26350 15986 26402
rect 26910 26350 26962 26402
rect 29598 26350 29650 26402
rect 30718 26350 30770 26402
rect 5070 26238 5122 26290
rect 6302 26238 6354 26290
rect 6750 26238 6802 26290
rect 6974 26238 7026 26290
rect 8430 26238 8482 26290
rect 8990 26238 9042 26290
rect 9998 26238 10050 26290
rect 10558 26238 10610 26290
rect 11902 26238 11954 26290
rect 12238 26238 12290 26290
rect 12686 26238 12738 26290
rect 13022 26238 13074 26290
rect 16158 26238 16210 26290
rect 16830 26238 16882 26290
rect 18174 26238 18226 26290
rect 18846 26238 18898 26290
rect 19182 26238 19234 26290
rect 19518 26238 19570 26290
rect 19742 26238 19794 26290
rect 20190 26238 20242 26290
rect 20638 26238 20690 26290
rect 20750 26238 20802 26290
rect 21646 26238 21698 26290
rect 25342 26238 25394 26290
rect 28814 26238 28866 26290
rect 29038 26238 29090 26290
rect 29486 26238 29538 26290
rect 32174 26238 32226 26290
rect 5182 26126 5234 26178
rect 5518 26126 5570 26178
rect 7086 26126 7138 26178
rect 8766 26126 8818 26178
rect 16606 26126 16658 26178
rect 17838 26126 17890 26178
rect 18734 26126 18786 26178
rect 19630 26126 19682 26178
rect 20414 26126 20466 26178
rect 22318 26126 22370 26178
rect 24446 26126 24498 26178
rect 28478 26126 28530 26178
rect 33182 26126 33234 26178
rect 10782 26014 10834 26066
rect 11230 26014 11282 26066
rect 11342 26014 11394 26066
rect 16382 26014 16434 26066
rect 17502 26014 17554 26066
rect 29486 26014 29538 26066
rect 5246 25846 5298 25898
rect 5350 25846 5402 25898
rect 5454 25846 5506 25898
rect 13310 25846 13362 25898
rect 13414 25846 13466 25898
rect 13518 25846 13570 25898
rect 21374 25846 21426 25898
rect 21478 25846 21530 25898
rect 21582 25846 21634 25898
rect 29438 25846 29490 25898
rect 29542 25846 29594 25898
rect 29646 25846 29698 25898
rect 9550 25678 9602 25730
rect 9886 25678 9938 25730
rect 16830 25678 16882 25730
rect 27806 25678 27858 25730
rect 4174 25566 4226 25618
rect 4622 25566 4674 25618
rect 5742 25566 5794 25618
rect 6526 25566 6578 25618
rect 9214 25566 9266 25618
rect 12126 25566 12178 25618
rect 15486 25566 15538 25618
rect 16942 25566 16994 25618
rect 17726 25566 17778 25618
rect 18958 25566 19010 25618
rect 27470 25566 27522 25618
rect 28254 25566 28306 25618
rect 31054 25566 31106 25618
rect 33182 25566 33234 25618
rect 4734 25454 4786 25506
rect 5182 25454 5234 25506
rect 7422 25454 7474 25506
rect 7758 25454 7810 25506
rect 10222 25454 10274 25506
rect 10558 25454 10610 25506
rect 6526 25398 6578 25450
rect 11006 25454 11058 25506
rect 11342 25454 11394 25506
rect 6302 25342 6354 25394
rect 6638 25342 6690 25394
rect 7198 25342 7250 25394
rect 9662 25342 9714 25394
rect 3950 25230 4002 25282
rect 4062 25230 4114 25282
rect 4510 25230 4562 25282
rect 6862 25230 6914 25282
rect 7086 25230 7138 25282
rect 9550 25230 9602 25282
rect 9998 25230 10050 25282
rect 10670 25230 10722 25282
rect 10894 25230 10946 25282
rect 11454 25286 11506 25338
rect 11678 25342 11730 25394
rect 12350 25342 12402 25394
rect 12574 25342 12626 25394
rect 12686 25398 12738 25450
rect 13918 25454 13970 25506
rect 14254 25454 14306 25506
rect 14478 25454 14530 25506
rect 15374 25454 15426 25506
rect 15822 25454 15874 25506
rect 16270 25454 16322 25506
rect 17502 25454 17554 25506
rect 17838 25454 17890 25506
rect 18510 25454 18562 25506
rect 18846 25454 18898 25506
rect 19182 25454 19234 25506
rect 26574 25454 26626 25506
rect 27022 25454 27074 25506
rect 27246 25454 27298 25506
rect 28142 25454 28194 25506
rect 29374 25454 29426 25506
rect 29710 25454 29762 25506
rect 30270 25454 30322 25506
rect 12910 25342 12962 25394
rect 13694 25342 13746 25394
rect 14926 25342 14978 25394
rect 15150 25342 15202 25394
rect 16494 25342 16546 25394
rect 17278 25342 17330 25394
rect 20526 25342 20578 25394
rect 20638 25342 20690 25394
rect 21982 25342 22034 25394
rect 27582 25342 27634 25394
rect 28590 25342 28642 25394
rect 14590 25230 14642 25282
rect 15486 25230 15538 25282
rect 16046 25230 16098 25282
rect 18062 25230 18114 25282
rect 19406 25230 19458 25282
rect 19518 25230 19570 25282
rect 19630 25230 19682 25282
rect 19854 25230 19906 25282
rect 20302 25230 20354 25282
rect 28366 25230 28418 25282
rect 29822 25230 29874 25282
rect 9278 25062 9330 25114
rect 9382 25062 9434 25114
rect 9486 25062 9538 25114
rect 17342 25062 17394 25114
rect 17446 25062 17498 25114
rect 17550 25062 17602 25114
rect 25406 25062 25458 25114
rect 25510 25062 25562 25114
rect 25614 25062 25666 25114
rect 33470 25062 33522 25114
rect 33574 25062 33626 25114
rect 33678 25062 33730 25114
rect 6862 24894 6914 24946
rect 7646 24894 7698 24946
rect 7758 24894 7810 24946
rect 8318 24894 8370 24946
rect 8542 24894 8594 24946
rect 10558 24894 10610 24946
rect 11678 24894 11730 24946
rect 12574 24894 12626 24946
rect 12686 24894 12738 24946
rect 13246 24894 13298 24946
rect 13358 24894 13410 24946
rect 15486 24894 15538 24946
rect 16494 24894 16546 24946
rect 18398 24894 18450 24946
rect 18846 24894 18898 24946
rect 24670 24894 24722 24946
rect 25566 24894 25618 24946
rect 2494 24782 2546 24834
rect 5294 24782 5346 24834
rect 12798 24782 12850 24834
rect 13470 24782 13522 24834
rect 14366 24782 14418 24834
rect 16270 24782 16322 24834
rect 16718 24782 16770 24834
rect 16830 24782 16882 24834
rect 17390 24782 17442 24834
rect 17502 24782 17554 24834
rect 18286 24782 18338 24834
rect 18734 24782 18786 24834
rect 20190 24782 20242 24834
rect 30718 24782 30770 24834
rect 33182 24782 33234 24834
rect 1822 24670 1874 24722
rect 5518 24670 5570 24722
rect 5966 24670 6018 24722
rect 6414 24670 6466 24722
rect 6750 24670 6802 24722
rect 6974 24670 7026 24722
rect 7310 24670 7362 24722
rect 7534 24670 7586 24722
rect 7982 24670 8034 24722
rect 8878 24670 8930 24722
rect 9550 24670 9602 24722
rect 9774 24670 9826 24722
rect 10894 24670 10946 24722
rect 13134 24670 13186 24722
rect 13918 24670 13970 24722
rect 14590 24670 14642 24722
rect 14926 24670 14978 24722
rect 15374 24670 15426 24722
rect 15598 24670 15650 24722
rect 15934 24670 15986 24722
rect 19294 24670 19346 24722
rect 19518 24670 19570 24722
rect 19854 24670 19906 24722
rect 20414 24670 20466 24722
rect 20638 24670 20690 24722
rect 21198 24670 21250 24722
rect 24334 24670 24386 24722
rect 25230 24670 25282 24722
rect 28142 24670 28194 24722
rect 28926 24670 28978 24722
rect 32510 24670 32562 24722
rect 4622 24558 4674 24610
rect 5406 24558 5458 24610
rect 8430 24558 8482 24610
rect 12238 24558 12290 24610
rect 19406 24558 19458 24610
rect 20302 24558 20354 24610
rect 21870 24558 21922 24610
rect 23998 24558 24050 24610
rect 27358 24558 27410 24610
rect 31950 24558 32002 24610
rect 9998 24446 10050 24498
rect 10110 24446 10162 24498
rect 17502 24446 17554 24498
rect 18846 24446 18898 24498
rect 33070 24446 33122 24498
rect 5246 24278 5298 24330
rect 5350 24278 5402 24330
rect 5454 24278 5506 24330
rect 13310 24278 13362 24330
rect 13414 24278 13466 24330
rect 13518 24278 13570 24330
rect 21374 24278 21426 24330
rect 21478 24278 21530 24330
rect 21582 24278 21634 24330
rect 29438 24278 29490 24330
rect 29542 24278 29594 24330
rect 29646 24278 29698 24330
rect 6414 24110 6466 24162
rect 19070 24110 19122 24162
rect 23102 24110 23154 24162
rect 26798 24110 26850 24162
rect 30830 24110 30882 24162
rect 4734 23998 4786 24050
rect 5966 23998 6018 24050
rect 7758 23998 7810 24050
rect 26350 23998 26402 24050
rect 27022 23998 27074 24050
rect 1822 23886 1874 23938
rect 6190 23886 6242 23938
rect 6638 23886 6690 23938
rect 7198 23886 7250 23938
rect 7870 23886 7922 23938
rect 8206 23886 8258 23938
rect 8766 23886 8818 23938
rect 10110 23886 10162 23938
rect 10446 23886 10498 23938
rect 11006 23886 11058 23938
rect 15262 23886 15314 23938
rect 15598 23886 15650 23938
rect 16270 23886 16322 23938
rect 18174 23886 18226 23938
rect 18510 23886 18562 23938
rect 18734 23886 18786 23938
rect 19182 23886 19234 23938
rect 19854 23886 19906 23938
rect 20078 23886 20130 23938
rect 20414 23886 20466 23938
rect 23438 23886 23490 23938
rect 27358 23886 27410 23938
rect 28030 23886 28082 23938
rect 28478 23886 28530 23938
rect 29150 23886 29202 23938
rect 30270 23886 30322 23938
rect 33182 23886 33234 23938
rect 2494 23774 2546 23826
rect 5854 23774 5906 23826
rect 6974 23774 7026 23826
rect 10670 23774 10722 23826
rect 11566 23774 11618 23826
rect 11902 23774 11954 23826
rect 12574 23774 12626 23826
rect 13918 23774 13970 23826
rect 15038 23774 15090 23826
rect 16158 23774 16210 23826
rect 16606 23774 16658 23826
rect 19630 23774 19682 23826
rect 21310 23774 21362 23826
rect 22430 23774 22482 23826
rect 22878 23774 22930 23826
rect 24222 23774 24274 23826
rect 27246 23774 27298 23826
rect 27582 23774 27634 23826
rect 29486 23774 29538 23826
rect 32734 23774 32786 23826
rect 7646 23662 7698 23714
rect 8430 23662 8482 23714
rect 8654 23662 8706 23714
rect 9886 23662 9938 23714
rect 10222 23662 10274 23714
rect 10782 23662 10834 23714
rect 11230 23662 11282 23714
rect 12238 23662 12290 23714
rect 12910 23662 12962 23714
rect 13582 23662 13634 23714
rect 14254 23662 14306 23714
rect 14702 23662 14754 23714
rect 16046 23662 16098 23714
rect 16942 23662 16994 23714
rect 17614 23662 17666 23714
rect 17838 23662 17890 23714
rect 19294 23662 19346 23714
rect 20078 23662 20130 23714
rect 21646 23662 21698 23714
rect 22094 23662 22146 23714
rect 22990 23662 23042 23714
rect 32622 23662 32674 23714
rect 32958 23662 33010 23714
rect 9278 23494 9330 23546
rect 9382 23494 9434 23546
rect 9486 23494 9538 23546
rect 17342 23494 17394 23546
rect 17446 23494 17498 23546
rect 17550 23494 17602 23546
rect 25406 23494 25458 23546
rect 25510 23494 25562 23546
rect 25614 23494 25666 23546
rect 33470 23494 33522 23546
rect 33574 23494 33626 23546
rect 33678 23494 33730 23546
rect 5406 23326 5458 23378
rect 6974 23326 7026 23378
rect 8654 23326 8706 23378
rect 20414 23326 20466 23378
rect 21310 23326 21362 23378
rect 22318 23326 22370 23378
rect 29486 23326 29538 23378
rect 30942 23326 30994 23378
rect 4846 23214 4898 23266
rect 5294 23214 5346 23266
rect 5518 23214 5570 23266
rect 5854 23214 5906 23266
rect 6750 23214 6802 23266
rect 7758 23214 7810 23266
rect 8878 23214 8930 23266
rect 8990 23214 9042 23266
rect 9550 23214 9602 23266
rect 12350 23214 12402 23266
rect 18510 23214 18562 23266
rect 18734 23214 18786 23266
rect 21534 23214 21586 23266
rect 22654 23214 22706 23266
rect 22990 23214 23042 23266
rect 28478 23214 28530 23266
rect 29374 23214 29426 23266
rect 33182 23214 33234 23266
rect 6190 23102 6242 23154
rect 6638 23102 6690 23154
rect 7198 23102 7250 23154
rect 7310 23102 7362 23154
rect 7422 23102 7474 23154
rect 9774 23102 9826 23154
rect 11566 23102 11618 23154
rect 18286 23102 18338 23154
rect 18398 23102 18450 23154
rect 19070 23102 19122 23154
rect 19966 23102 20018 23154
rect 20638 23102 20690 23154
rect 21646 23102 21698 23154
rect 22542 23102 22594 23154
rect 23326 23102 23378 23154
rect 23886 23102 23938 23154
rect 25566 23102 25618 23154
rect 28254 23102 28306 23154
rect 28702 23102 28754 23154
rect 29934 23102 29986 23154
rect 16718 22990 16770 23042
rect 17502 22990 17554 23042
rect 24446 22990 24498 23042
rect 27470 22990 27522 23042
rect 15822 22878 15874 22930
rect 16270 22878 16322 22930
rect 16494 22878 16546 22930
rect 19182 22878 19234 22930
rect 19518 22878 19570 22930
rect 19630 22878 19682 22930
rect 19854 22878 19906 22930
rect 28142 22878 28194 22930
rect 28926 22878 28978 22930
rect 29486 22878 29538 22930
rect 33070 22878 33122 22930
rect 5246 22710 5298 22762
rect 5350 22710 5402 22762
rect 5454 22710 5506 22762
rect 13310 22710 13362 22762
rect 13414 22710 13466 22762
rect 13518 22710 13570 22762
rect 21374 22710 21426 22762
rect 21478 22710 21530 22762
rect 21582 22710 21634 22762
rect 29438 22710 29490 22762
rect 29542 22710 29594 22762
rect 29646 22710 29698 22762
rect 11342 22542 11394 22594
rect 15038 22542 15090 22594
rect 15374 22542 15426 22594
rect 18062 22542 18114 22594
rect 18622 22542 18674 22594
rect 20750 22542 20802 22594
rect 32958 22542 33010 22594
rect 4622 22430 4674 22482
rect 5070 22430 5122 22482
rect 5854 22430 5906 22482
rect 14814 22430 14866 22482
rect 18622 22430 18674 22482
rect 24894 22430 24946 22482
rect 25566 22430 25618 22482
rect 27582 22430 27634 22482
rect 1822 22318 1874 22370
rect 10894 22318 10946 22370
rect 12910 22318 12962 22370
rect 16158 22318 16210 22370
rect 16270 22318 16322 22370
rect 16718 22318 16770 22370
rect 18846 22318 18898 22370
rect 19182 22318 19234 22370
rect 21982 22318 22034 22370
rect 25454 22318 25506 22370
rect 25902 22318 25954 22370
rect 28142 22318 28194 22370
rect 29486 22318 29538 22370
rect 30270 22318 30322 22370
rect 31054 22318 31106 22370
rect 2494 22206 2546 22258
rect 11454 22206 11506 22258
rect 11790 22206 11842 22258
rect 12574 22206 12626 22258
rect 13470 22206 13522 22258
rect 13806 22206 13858 22258
rect 14142 22206 14194 22258
rect 14478 22206 14530 22258
rect 17390 22206 17442 22258
rect 20638 22206 20690 22258
rect 21646 22206 21698 22258
rect 22766 22206 22818 22258
rect 26798 22206 26850 22258
rect 27134 22206 27186 22258
rect 27246 22206 27298 22258
rect 27918 22206 27970 22258
rect 28478 22206 28530 22258
rect 29934 22206 29986 22258
rect 30158 22206 30210 22258
rect 11342 22094 11394 22146
rect 12126 22094 12178 22146
rect 15822 22094 15874 22146
rect 16382 22094 16434 22146
rect 17054 22094 17106 22146
rect 18174 22094 18226 22146
rect 19406 22094 19458 22146
rect 19518 22094 19570 22146
rect 19966 22094 20018 22146
rect 20414 22094 20466 22146
rect 21310 22094 21362 22146
rect 21534 22094 21586 22146
rect 25118 22094 25170 22146
rect 27022 22094 27074 22146
rect 28366 22094 28418 22146
rect 29262 22094 29314 22146
rect 9278 21926 9330 21978
rect 9382 21926 9434 21978
rect 9486 21926 9538 21978
rect 17342 21926 17394 21978
rect 17446 21926 17498 21978
rect 17550 21926 17602 21978
rect 25406 21926 25458 21978
rect 25510 21926 25562 21978
rect 25614 21926 25666 21978
rect 33470 21926 33522 21978
rect 33574 21926 33626 21978
rect 33678 21926 33730 21978
rect 5294 21758 5346 21810
rect 6190 21758 6242 21810
rect 6750 21758 6802 21810
rect 11342 21758 11394 21810
rect 13246 21758 13298 21810
rect 14366 21758 14418 21810
rect 16046 21758 16098 21810
rect 16494 21758 16546 21810
rect 23774 21758 23826 21810
rect 23886 21758 23938 21810
rect 6078 21646 6130 21698
rect 7534 21646 7586 21698
rect 7646 21646 7698 21698
rect 9550 21646 9602 21698
rect 9662 21646 9714 21698
rect 12910 21646 12962 21698
rect 13022 21646 13074 21698
rect 22878 21646 22930 21698
rect 24222 21646 24274 21698
rect 24446 21646 24498 21698
rect 24670 21646 24722 21698
rect 25342 21646 25394 21698
rect 27134 21646 27186 21698
rect 28254 21646 28306 21698
rect 32062 21646 32114 21698
rect 1822 21534 1874 21586
rect 4958 21534 5010 21586
rect 5294 21534 5346 21586
rect 5630 21534 5682 21586
rect 6638 21534 6690 21586
rect 6974 21534 7026 21586
rect 7310 21534 7362 21586
rect 7870 21534 7922 21586
rect 8318 21534 8370 21586
rect 8430 21534 8482 21586
rect 9886 21534 9938 21586
rect 11118 21534 11170 21586
rect 12126 21534 12178 21586
rect 12574 21534 12626 21586
rect 14142 21534 14194 21586
rect 14814 21534 14866 21586
rect 18734 21534 18786 21586
rect 23214 21534 23266 21586
rect 23662 21534 23714 21586
rect 25230 21534 25282 21586
rect 25790 21534 25842 21586
rect 26910 21534 26962 21586
rect 29822 21534 29874 21586
rect 30270 21534 30322 21586
rect 2494 21422 2546 21474
rect 4622 21422 4674 21474
rect 8094 21422 8146 21474
rect 10334 21422 10386 21474
rect 13694 21422 13746 21474
rect 15486 21422 15538 21474
rect 16942 21422 16994 21474
rect 17614 21422 17666 21474
rect 17950 21422 18002 21474
rect 18398 21422 18450 21474
rect 19518 21422 19570 21474
rect 21646 21422 21698 21474
rect 22318 21422 22370 21474
rect 26126 21422 26178 21474
rect 27022 21422 27074 21474
rect 30718 21422 30770 21474
rect 31726 21422 31778 21474
rect 33182 21422 33234 21474
rect 6190 21310 6242 21362
rect 22654 21310 22706 21362
rect 22990 21310 23042 21362
rect 24782 21310 24834 21362
rect 31838 21310 31890 21362
rect 5246 21142 5298 21194
rect 5350 21142 5402 21194
rect 5454 21142 5506 21194
rect 13310 21142 13362 21194
rect 13414 21142 13466 21194
rect 13518 21142 13570 21194
rect 21374 21142 21426 21194
rect 21478 21142 21530 21194
rect 21582 21142 21634 21194
rect 29438 21142 29490 21194
rect 29542 21142 29594 21194
rect 29646 21142 29698 21194
rect 5742 20974 5794 21026
rect 4174 20862 4226 20914
rect 5070 20862 5122 20914
rect 7982 20862 8034 20914
rect 10110 20862 10162 20914
rect 12014 20862 12066 20914
rect 16382 20862 16434 20914
rect 17390 20862 17442 20914
rect 19294 20862 19346 20914
rect 20862 20862 20914 20914
rect 24222 20862 24274 20914
rect 26126 20862 26178 20914
rect 27246 20862 27298 20914
rect 27694 20862 27746 20914
rect 30382 20862 30434 20914
rect 33294 20862 33346 20914
rect 4286 20750 4338 20802
rect 4622 20750 4674 20802
rect 5854 20750 5906 20802
rect 6190 20750 6242 20802
rect 6638 20750 6690 20802
rect 6862 20750 6914 20802
rect 7198 20750 7250 20802
rect 13470 20750 13522 20802
rect 17838 20750 17890 20802
rect 18286 20750 18338 20802
rect 19182 20750 19234 20802
rect 19518 20750 19570 20802
rect 19966 20750 20018 20802
rect 20302 20750 20354 20802
rect 21422 20750 21474 20802
rect 25342 20750 25394 20802
rect 25678 20750 25730 20802
rect 26910 20750 26962 20802
rect 27358 20750 27410 20802
rect 27918 20750 27970 20802
rect 28366 20750 28418 20802
rect 29150 20750 29202 20802
rect 32062 20750 32114 20802
rect 4062 20638 4114 20690
rect 11006 20638 11058 20690
rect 14254 20638 14306 20690
rect 17614 20638 17666 20690
rect 18846 20638 18898 20690
rect 19742 20638 19794 20690
rect 22094 20638 22146 20690
rect 26798 20638 26850 20690
rect 27134 20638 27186 20690
rect 28142 20638 28194 20690
rect 32398 20638 32450 20690
rect 32734 20638 32786 20690
rect 5742 20526 5794 20578
rect 6526 20526 6578 20578
rect 10670 20526 10722 20578
rect 10894 20526 10946 20578
rect 11566 20526 11618 20578
rect 16830 20526 16882 20578
rect 18062 20526 18114 20578
rect 19630 20526 19682 20578
rect 24670 20526 24722 20578
rect 24894 20526 24946 20578
rect 28702 20526 28754 20578
rect 9278 20358 9330 20410
rect 9382 20358 9434 20410
rect 9486 20358 9538 20410
rect 17342 20358 17394 20410
rect 17446 20358 17498 20410
rect 17550 20358 17602 20410
rect 25406 20358 25458 20410
rect 25510 20358 25562 20410
rect 25614 20358 25666 20410
rect 33470 20358 33522 20410
rect 33574 20358 33626 20410
rect 33678 20358 33730 20410
rect 4286 20190 4338 20242
rect 4510 20190 4562 20242
rect 5406 20190 5458 20242
rect 14366 20190 14418 20242
rect 15262 20190 15314 20242
rect 16158 20190 16210 20242
rect 16942 20190 16994 20242
rect 25342 20190 25394 20242
rect 25678 20190 25730 20242
rect 6526 20078 6578 20130
rect 13022 20078 13074 20130
rect 13694 20078 13746 20130
rect 18174 20078 18226 20130
rect 20974 20078 21026 20130
rect 22430 20078 22482 20130
rect 22542 20078 22594 20130
rect 22878 20078 22930 20130
rect 27246 20078 27298 20130
rect 28366 20078 28418 20130
rect 30494 20078 30546 20130
rect 31838 20078 31890 20130
rect 32174 20078 32226 20130
rect 4622 19966 4674 20018
rect 5182 19966 5234 20018
rect 5742 19966 5794 20018
rect 9774 19966 9826 20018
rect 13582 19966 13634 20018
rect 13918 19966 13970 20018
rect 14142 19966 14194 20018
rect 14366 19966 14418 20018
rect 14590 19966 14642 20018
rect 15038 19966 15090 20018
rect 15374 19966 15426 20018
rect 16046 19966 16098 20018
rect 16382 19966 16434 20018
rect 17502 19966 17554 20018
rect 23102 19966 23154 20018
rect 23550 19966 23602 20018
rect 23774 19966 23826 20018
rect 27358 19966 27410 20018
rect 29822 19966 29874 20018
rect 30270 19966 30322 20018
rect 31054 19966 31106 20018
rect 31502 19966 31554 20018
rect 32510 19966 32562 20018
rect 33182 19966 33234 20018
rect 8654 19854 8706 19906
rect 10446 19854 10498 19906
rect 12574 19854 12626 19906
rect 20302 19854 20354 19906
rect 21534 19854 21586 19906
rect 21982 19854 22034 19906
rect 22990 19854 23042 19906
rect 24222 19854 24274 19906
rect 26238 19854 26290 19906
rect 27022 19854 27074 19906
rect 22430 19742 22482 19794
rect 26014 19742 26066 19794
rect 33070 19742 33122 19794
rect 5246 19574 5298 19626
rect 5350 19574 5402 19626
rect 5454 19574 5506 19626
rect 13310 19574 13362 19626
rect 13414 19574 13466 19626
rect 13518 19574 13570 19626
rect 21374 19574 21426 19626
rect 21478 19574 21530 19626
rect 21582 19574 21634 19626
rect 29438 19574 29490 19626
rect 29542 19574 29594 19626
rect 29646 19574 29698 19626
rect 5742 19406 5794 19458
rect 18846 19406 18898 19458
rect 19966 19406 20018 19458
rect 20302 19406 20354 19458
rect 20526 19406 20578 19458
rect 22094 19406 22146 19458
rect 22878 19406 22930 19458
rect 23774 19406 23826 19458
rect 24334 19406 24386 19458
rect 29150 19406 29202 19458
rect 30830 19406 30882 19458
rect 4622 19294 4674 19346
rect 5070 19294 5122 19346
rect 9550 19294 9602 19346
rect 10558 19294 10610 19346
rect 12910 19294 12962 19346
rect 17054 19294 17106 19346
rect 19070 19294 19122 19346
rect 19406 19294 19458 19346
rect 19966 19294 20018 19346
rect 20302 19294 20354 19346
rect 21870 19294 21922 19346
rect 25118 19294 25170 19346
rect 27806 19294 27858 19346
rect 32846 19294 32898 19346
rect 1822 19182 1874 19234
rect 5854 19182 5906 19234
rect 7870 19182 7922 19234
rect 8766 19182 8818 19234
rect 10334 19182 10386 19234
rect 10670 19182 10722 19234
rect 10894 19182 10946 19234
rect 13582 19182 13634 19234
rect 14142 19182 14194 19234
rect 17502 19182 17554 19234
rect 22990 19182 23042 19234
rect 23886 19182 23938 19234
rect 24446 19182 24498 19234
rect 25006 19182 25058 19234
rect 26014 19182 26066 19234
rect 26798 19182 26850 19234
rect 28030 19182 28082 19234
rect 29486 19182 29538 19234
rect 30046 19182 30098 19234
rect 2494 19070 2546 19122
rect 8206 19070 8258 19122
rect 8990 19070 9042 19122
rect 9102 19070 9154 19122
rect 11454 19070 11506 19122
rect 11566 19070 11618 19122
rect 14926 19070 14978 19122
rect 17726 19070 17778 19122
rect 23326 19070 23378 19122
rect 24334 19070 24386 19122
rect 25454 19070 25506 19122
rect 26238 19070 26290 19122
rect 26350 19070 26402 19122
rect 27694 19070 27746 19122
rect 28366 19070 28418 19122
rect 5742 18958 5794 19010
rect 8094 18958 8146 19010
rect 11230 18958 11282 19010
rect 13694 18958 13746 19010
rect 13918 18958 13970 19010
rect 18286 18958 18338 19010
rect 20750 18958 20802 19010
rect 21534 18958 21586 19010
rect 22318 18958 22370 19010
rect 22878 18958 22930 19010
rect 23214 18958 23266 19010
rect 23774 18958 23826 19010
rect 26126 18958 26178 19010
rect 28478 18958 28530 19010
rect 28702 18958 28754 19010
rect 29262 18958 29314 19010
rect 9278 18790 9330 18842
rect 9382 18790 9434 18842
rect 9486 18790 9538 18842
rect 17342 18790 17394 18842
rect 17446 18790 17498 18842
rect 17550 18790 17602 18842
rect 25406 18790 25458 18842
rect 25510 18790 25562 18842
rect 25614 18790 25666 18842
rect 33470 18790 33522 18842
rect 33574 18790 33626 18842
rect 33678 18790 33730 18842
rect 3054 18622 3106 18674
rect 3614 18622 3666 18674
rect 5966 18622 6018 18674
rect 8206 18622 8258 18674
rect 11790 18622 11842 18674
rect 13134 18622 13186 18674
rect 14926 18622 14978 18674
rect 15486 18622 15538 18674
rect 18622 18622 18674 18674
rect 26686 18622 26738 18674
rect 27918 18622 27970 18674
rect 33070 18622 33122 18674
rect 2942 18510 2994 18562
rect 3726 18510 3778 18562
rect 5070 18510 5122 18562
rect 5182 18510 5234 18562
rect 7422 18510 7474 18562
rect 11342 18510 11394 18562
rect 11678 18510 11730 18562
rect 13022 18510 13074 18562
rect 13358 18510 13410 18562
rect 15038 18510 15090 18562
rect 15598 18510 15650 18562
rect 16046 18510 16098 18562
rect 16158 18510 16210 18562
rect 19966 18510 20018 18562
rect 22766 18510 22818 18562
rect 24110 18510 24162 18562
rect 26462 18510 26514 18562
rect 27246 18510 27298 18562
rect 27694 18510 27746 18562
rect 30494 18510 30546 18562
rect 31726 18510 31778 18562
rect 32174 18510 32226 18562
rect 3278 18398 3330 18450
rect 3950 18398 4002 18450
rect 4398 18398 4450 18450
rect 4510 18398 4562 18450
rect 4846 18398 4898 18450
rect 6302 18398 6354 18450
rect 6750 18398 6802 18450
rect 7758 18398 7810 18450
rect 8542 18398 8594 18450
rect 8990 18398 9042 18450
rect 10894 18398 10946 18450
rect 11118 18398 11170 18450
rect 12014 18398 12066 18450
rect 13470 18398 13522 18450
rect 13918 18398 13970 18450
rect 14030 18398 14082 18450
rect 14478 18398 14530 18450
rect 14814 18398 14866 18450
rect 15262 18398 15314 18450
rect 15822 18398 15874 18450
rect 19854 18398 19906 18450
rect 20526 18398 20578 18450
rect 21310 18398 21362 18450
rect 21534 18398 21586 18450
rect 21646 18398 21698 18450
rect 22094 18398 22146 18450
rect 23102 18398 23154 18450
rect 23438 18398 23490 18450
rect 23774 18398 23826 18450
rect 24670 18398 24722 18450
rect 25454 18398 25506 18450
rect 25902 18398 25954 18450
rect 26350 18398 26402 18450
rect 28254 18398 28306 18450
rect 28702 18398 28754 18450
rect 29598 18398 29650 18450
rect 30270 18398 30322 18450
rect 30942 18398 30994 18450
rect 31502 18398 31554 18450
rect 32286 18398 32338 18450
rect 4174 18286 4226 18338
rect 11230 18286 11282 18338
rect 13694 18286 13746 18338
rect 18958 18286 19010 18338
rect 20974 18286 21026 18338
rect 28590 18286 28642 18338
rect 29262 18286 29314 18338
rect 30046 18286 30098 18338
rect 30382 18286 30434 18338
rect 33182 18286 33234 18338
rect 3614 18174 3666 18226
rect 19182 18174 19234 18226
rect 19518 18174 19570 18226
rect 19966 18174 20018 18226
rect 23438 18174 23490 18226
rect 27582 18174 27634 18226
rect 29822 18174 29874 18226
rect 5246 18006 5298 18058
rect 5350 18006 5402 18058
rect 5454 18006 5506 18058
rect 13310 18006 13362 18058
rect 13414 18006 13466 18058
rect 13518 18006 13570 18058
rect 21374 18006 21426 18058
rect 21478 18006 21530 18058
rect 21582 18006 21634 18058
rect 29438 18006 29490 18058
rect 29542 18006 29594 18058
rect 29646 18006 29698 18058
rect 20750 17838 20802 17890
rect 27470 17838 27522 17890
rect 27918 17838 27970 17890
rect 31726 17838 31778 17890
rect 4622 17726 4674 17778
rect 5070 17726 5122 17778
rect 9886 17726 9938 17778
rect 12014 17726 12066 17778
rect 14254 17726 14306 17778
rect 16382 17726 16434 17778
rect 16830 17726 16882 17778
rect 17614 17726 17666 17778
rect 17838 17726 17890 17778
rect 21982 17726 22034 17778
rect 22206 17726 22258 17778
rect 24782 17726 24834 17778
rect 28590 17726 28642 17778
rect 30718 17726 30770 17778
rect 1822 17614 1874 17666
rect 5854 17614 5906 17666
rect 7086 17614 7138 17666
rect 7310 17614 7362 17666
rect 9214 17614 9266 17666
rect 13582 17614 13634 17666
rect 18510 17614 18562 17666
rect 18958 17614 19010 17666
rect 19854 17614 19906 17666
rect 23214 17614 23266 17666
rect 26798 17614 26850 17666
rect 27694 17614 27746 17666
rect 28142 17614 28194 17666
rect 30606 17614 30658 17666
rect 31278 17614 31330 17666
rect 31502 17614 31554 17666
rect 2494 17502 2546 17554
rect 5630 17502 5682 17554
rect 6750 17502 6802 17554
rect 7646 17502 7698 17554
rect 8542 17502 8594 17554
rect 12350 17502 12402 17554
rect 18174 17502 18226 17554
rect 18846 17502 18898 17554
rect 19630 17502 19682 17554
rect 19966 17502 20018 17554
rect 20638 17502 20690 17554
rect 21310 17502 21362 17554
rect 21646 17502 21698 17554
rect 22542 17502 22594 17554
rect 22990 17502 23042 17554
rect 23998 17502 24050 17554
rect 25342 17502 25394 17554
rect 25902 17502 25954 17554
rect 26462 17502 26514 17554
rect 33182 17502 33234 17554
rect 7534 17390 7586 17442
rect 8206 17390 8258 17442
rect 12686 17390 12738 17442
rect 17950 17390 18002 17442
rect 18622 17390 18674 17442
rect 19406 17390 19458 17442
rect 19518 17390 19570 17442
rect 23438 17390 23490 17442
rect 24222 17390 24274 17442
rect 24446 17390 24498 17442
rect 24558 17390 24610 17442
rect 25790 17390 25842 17442
rect 27022 17390 27074 17442
rect 33070 17390 33122 17442
rect 9278 17222 9330 17274
rect 9382 17222 9434 17274
rect 9486 17222 9538 17274
rect 17342 17222 17394 17274
rect 17446 17222 17498 17274
rect 17550 17222 17602 17274
rect 25406 17222 25458 17274
rect 25510 17222 25562 17274
rect 25614 17222 25666 17274
rect 33470 17222 33522 17274
rect 33574 17222 33626 17274
rect 33678 17222 33730 17274
rect 4510 17054 4562 17106
rect 5182 17054 5234 17106
rect 5630 17054 5682 17106
rect 6638 17054 6690 17106
rect 8206 17054 8258 17106
rect 8766 17054 8818 17106
rect 9662 17054 9714 17106
rect 10894 17054 10946 17106
rect 12350 17054 12402 17106
rect 14254 17054 14306 17106
rect 24558 17054 24610 17106
rect 26574 17054 26626 17106
rect 28366 17054 28418 17106
rect 28814 17054 28866 17106
rect 4174 16942 4226 16994
rect 4398 16942 4450 16994
rect 4958 16942 5010 16994
rect 5294 16942 5346 16994
rect 5854 16942 5906 16994
rect 5966 16942 6018 16994
rect 6302 16942 6354 16994
rect 6414 16942 6466 16994
rect 6862 16942 6914 16994
rect 7870 16942 7922 16994
rect 7982 16942 8034 16994
rect 8430 16942 8482 16994
rect 11230 16942 11282 16994
rect 20078 16942 20130 16994
rect 23662 16942 23714 16994
rect 23886 16942 23938 16994
rect 26014 16942 26066 16994
rect 26126 16942 26178 16994
rect 26238 16942 26290 16994
rect 29374 16942 29426 16994
rect 30270 16942 30322 16994
rect 31278 16942 31330 16994
rect 33182 16942 33234 16994
rect 4846 16830 4898 16882
rect 7086 16830 7138 16882
rect 10670 16830 10722 16882
rect 11566 16830 11618 16882
rect 13918 16830 13970 16882
rect 16830 16830 16882 16882
rect 22766 16830 22818 16882
rect 24110 16830 24162 16882
rect 27358 16830 27410 16882
rect 27470 16830 27522 16882
rect 30046 16830 30098 16882
rect 31166 16830 31218 16882
rect 31390 16830 31442 16882
rect 32062 16830 32114 16882
rect 23550 16718 23602 16770
rect 27806 16718 27858 16770
rect 29150 16718 29202 16770
rect 30270 16718 30322 16770
rect 25566 16606 25618 16658
rect 5246 16438 5298 16490
rect 5350 16438 5402 16490
rect 5454 16438 5506 16490
rect 13310 16438 13362 16490
rect 13414 16438 13466 16490
rect 13518 16438 13570 16490
rect 21374 16438 21426 16490
rect 21478 16438 21530 16490
rect 21582 16438 21634 16490
rect 29438 16438 29490 16490
rect 29542 16438 29594 16490
rect 29646 16438 29698 16490
rect 18510 16270 18562 16322
rect 19294 16270 19346 16322
rect 23550 16270 23602 16322
rect 7534 16158 7586 16210
rect 16942 16158 16994 16210
rect 18734 16158 18786 16210
rect 22206 16158 22258 16210
rect 26014 16158 26066 16210
rect 26686 16158 26738 16210
rect 27470 16158 27522 16210
rect 31502 16158 31554 16210
rect 32622 16158 32674 16210
rect 3838 16046 3890 16098
rect 4958 16046 5010 16098
rect 5630 16046 5682 16098
rect 5966 16046 6018 16098
rect 6414 16046 6466 16098
rect 10894 16046 10946 16098
rect 11678 16046 11730 16098
rect 16382 16046 16434 16098
rect 18622 16046 18674 16098
rect 19070 16046 19122 16098
rect 20190 16046 20242 16098
rect 20526 16046 20578 16098
rect 21310 16046 21362 16098
rect 22654 16046 22706 16098
rect 23214 16046 23266 16098
rect 23886 16046 23938 16098
rect 24110 16046 24162 16098
rect 24782 16046 24834 16098
rect 25006 16046 25058 16098
rect 27022 16046 27074 16098
rect 28030 16046 28082 16098
rect 28254 16046 28306 16098
rect 29374 16046 29426 16098
rect 30270 16046 30322 16098
rect 31950 16046 32002 16098
rect 32958 16046 33010 16098
rect 4174 15934 4226 15986
rect 4398 15934 4450 15986
rect 4734 15934 4786 15986
rect 6190 15934 6242 15986
rect 6750 15934 6802 15986
rect 11342 15934 11394 15986
rect 16830 15934 16882 15986
rect 17054 15934 17106 15986
rect 17614 15934 17666 15986
rect 17838 15934 17890 15986
rect 17950 15934 18002 15986
rect 21534 15934 21586 15986
rect 21646 15934 21698 15986
rect 22542 15934 22594 15986
rect 27694 15934 27746 15986
rect 29150 15934 29202 15986
rect 30606 15934 30658 15986
rect 30830 15934 30882 15986
rect 3950 15822 4002 15874
rect 4510 15822 4562 15874
rect 5966 15822 6018 15874
rect 6638 15822 6690 15874
rect 10558 15822 10610 15874
rect 16606 15822 16658 15874
rect 18062 15822 18114 15874
rect 18174 15822 18226 15874
rect 19742 15822 19794 15874
rect 19854 15822 19906 15874
rect 19966 15822 20018 15874
rect 24446 15822 24498 15874
rect 25566 15822 25618 15874
rect 28478 15822 28530 15874
rect 28590 15878 28642 15930
rect 29934 15822 29986 15874
rect 9278 15654 9330 15706
rect 9382 15654 9434 15706
rect 9486 15654 9538 15706
rect 17342 15654 17394 15706
rect 17446 15654 17498 15706
rect 17550 15654 17602 15706
rect 25406 15654 25458 15706
rect 25510 15654 25562 15706
rect 25614 15654 25666 15706
rect 33470 15654 33522 15706
rect 33574 15654 33626 15706
rect 33678 15654 33730 15706
rect 5070 15486 5122 15538
rect 5294 15486 5346 15538
rect 6750 15486 6802 15538
rect 7646 15486 7698 15538
rect 8206 15486 8258 15538
rect 10446 15486 10498 15538
rect 12350 15486 12402 15538
rect 17838 15486 17890 15538
rect 18510 15486 18562 15538
rect 19070 15486 19122 15538
rect 19294 15486 19346 15538
rect 21198 15486 21250 15538
rect 22878 15486 22930 15538
rect 23214 15486 23266 15538
rect 24670 15486 24722 15538
rect 28142 15486 28194 15538
rect 28254 15486 28306 15538
rect 29150 15486 29202 15538
rect 2494 15374 2546 15426
rect 6414 15374 6466 15426
rect 6974 15374 7026 15426
rect 8318 15374 8370 15426
rect 10222 15374 10274 15426
rect 13358 15374 13410 15426
rect 18398 15374 18450 15426
rect 18734 15374 18786 15426
rect 19406 15374 19458 15426
rect 20526 15374 20578 15426
rect 20750 15374 20802 15426
rect 21310 15374 21362 15426
rect 21646 15374 21698 15426
rect 23550 15374 23602 15426
rect 24110 15374 24162 15426
rect 25790 15374 25842 15426
rect 26910 15374 26962 15426
rect 27918 15374 27970 15426
rect 28702 15374 28754 15426
rect 33182 15374 33234 15426
rect 1822 15262 1874 15314
rect 5406 15262 5458 15314
rect 5854 15262 5906 15314
rect 6302 15262 6354 15314
rect 6638 15262 6690 15314
rect 7086 15262 7138 15314
rect 7534 15262 7586 15314
rect 7870 15262 7922 15314
rect 7982 15262 8034 15314
rect 10558 15262 10610 15314
rect 10670 15262 10722 15314
rect 11230 15262 11282 15314
rect 13134 15262 13186 15314
rect 13694 15262 13746 15314
rect 18174 15262 18226 15314
rect 18286 15262 18338 15314
rect 20078 15262 20130 15314
rect 20302 15262 20354 15314
rect 20862 15262 20914 15314
rect 21982 15262 22034 15314
rect 23886 15262 23938 15314
rect 24222 15262 24274 15314
rect 25678 15262 25730 15314
rect 26014 15262 26066 15314
rect 26574 15262 26626 15314
rect 27582 15262 27634 15314
rect 28478 15262 28530 15314
rect 29598 15262 29650 15314
rect 4622 15150 4674 15202
rect 12014 15150 12066 15202
rect 12238 15150 12290 15202
rect 14478 15150 14530 15202
rect 16606 15150 16658 15202
rect 22430 15150 22482 15202
rect 30382 15150 30434 15202
rect 32510 15150 32562 15202
rect 19742 15038 19794 15090
rect 25230 15038 25282 15090
rect 5246 14870 5298 14922
rect 5350 14870 5402 14922
rect 5454 14870 5506 14922
rect 13310 14870 13362 14922
rect 13414 14870 13466 14922
rect 13518 14870 13570 14922
rect 21374 14870 21426 14922
rect 21478 14870 21530 14922
rect 21582 14870 21634 14922
rect 29438 14870 29490 14922
rect 29542 14870 29594 14922
rect 29646 14870 29698 14922
rect 17166 14702 17218 14754
rect 2494 14590 2546 14642
rect 4622 14590 4674 14642
rect 5182 14590 5234 14642
rect 8990 14590 9042 14642
rect 11118 14590 11170 14642
rect 16382 14590 16434 14642
rect 18510 14590 18562 14642
rect 24670 14590 24722 14642
rect 25678 14590 25730 14642
rect 29150 14590 29202 14642
rect 30270 14590 30322 14642
rect 1822 14478 1874 14530
rect 6526 14478 6578 14530
rect 6862 14478 6914 14530
rect 7198 14478 7250 14530
rect 7646 14478 7698 14530
rect 7870 14478 7922 14530
rect 8654 14478 8706 14530
rect 11902 14478 11954 14530
rect 12574 14478 12626 14530
rect 13582 14478 13634 14530
rect 17950 14478 18002 14530
rect 18286 14478 18338 14530
rect 18622 14478 18674 14530
rect 18958 14478 19010 14530
rect 20078 14478 20130 14530
rect 20526 14478 20578 14530
rect 23438 14478 23490 14530
rect 23774 14478 23826 14530
rect 28590 14478 28642 14530
rect 33070 14478 33122 14530
rect 8094 14366 8146 14418
rect 8318 14366 8370 14418
rect 14254 14366 14306 14418
rect 17838 14366 17890 14418
rect 19518 14366 19570 14418
rect 22654 14366 22706 14418
rect 23662 14366 23714 14418
rect 27806 14366 27858 14418
rect 32398 14366 32450 14418
rect 6750 14254 6802 14306
rect 7870 14254 7922 14306
rect 8542 14254 8594 14306
rect 12238 14254 12290 14306
rect 16830 14254 16882 14306
rect 19182 14254 19234 14306
rect 19406 14254 19458 14306
rect 20638 14254 20690 14306
rect 21422 14254 21474 14306
rect 29710 14254 29762 14306
rect 9278 14086 9330 14138
rect 9382 14086 9434 14138
rect 9486 14086 9538 14138
rect 17342 14086 17394 14138
rect 17446 14086 17498 14138
rect 17550 14086 17602 14138
rect 25406 14086 25458 14138
rect 25510 14086 25562 14138
rect 25614 14086 25666 14138
rect 33470 14086 33522 14138
rect 33574 14086 33626 14138
rect 33678 14086 33730 14138
rect 10558 13918 10610 13970
rect 10670 13918 10722 13970
rect 10782 13918 10834 13970
rect 12462 13918 12514 13970
rect 14142 13918 14194 13970
rect 15150 13918 15202 13970
rect 17838 13918 17890 13970
rect 18510 13918 18562 13970
rect 19294 13918 19346 13970
rect 22878 13918 22930 13970
rect 23886 13918 23938 13970
rect 6862 13806 6914 13858
rect 11006 13806 11058 13858
rect 11566 13806 11618 13858
rect 20190 13862 20242 13914
rect 25454 13918 25506 13970
rect 30046 13918 30098 13970
rect 31726 13918 31778 13970
rect 32174 13918 32226 13970
rect 14478 13806 14530 13858
rect 16606 13806 16658 13858
rect 20302 13806 20354 13858
rect 21086 13806 21138 13858
rect 21646 13806 21698 13858
rect 22094 13806 22146 13858
rect 23102 13806 23154 13858
rect 23774 13806 23826 13858
rect 25566 13806 25618 13858
rect 27918 13806 27970 13858
rect 28926 13806 28978 13858
rect 30606 13806 30658 13858
rect 31166 13806 31218 13858
rect 31614 13806 31666 13858
rect 6190 13694 6242 13746
rect 11902 13694 11954 13746
rect 14814 13694 14866 13746
rect 16718 13694 16770 13746
rect 17614 13694 17666 13746
rect 17726 13694 17778 13746
rect 18174 13694 18226 13746
rect 18398 13694 18450 13746
rect 18734 13694 18786 13746
rect 18958 13694 19010 13746
rect 20526 13694 20578 13746
rect 21758 13694 21810 13746
rect 23326 13694 23378 13746
rect 23998 13694 24050 13746
rect 24334 13694 24386 13746
rect 25230 13694 25282 13746
rect 26574 13694 26626 13746
rect 26910 13694 26962 13746
rect 27470 13694 27522 13746
rect 28254 13694 28306 13746
rect 29038 13694 29090 13746
rect 30382 13694 30434 13746
rect 32510 13694 32562 13746
rect 8990 13582 9042 13634
rect 10222 13582 10274 13634
rect 11678 13582 11730 13634
rect 15934 13582 15986 13634
rect 19854 13582 19906 13634
rect 26126 13582 26178 13634
rect 29598 13582 29650 13634
rect 33182 13582 33234 13634
rect 15598 13470 15650 13522
rect 19630 13470 19682 13522
rect 22206 13470 22258 13522
rect 31726 13470 31778 13522
rect 5246 13302 5298 13354
rect 5350 13302 5402 13354
rect 5454 13302 5506 13354
rect 13310 13302 13362 13354
rect 13414 13302 13466 13354
rect 13518 13302 13570 13354
rect 21374 13302 21426 13354
rect 21478 13302 21530 13354
rect 21582 13302 21634 13354
rect 29438 13302 29490 13354
rect 29542 13302 29594 13354
rect 29646 13302 29698 13354
rect 17950 13134 18002 13186
rect 19070 13134 19122 13186
rect 22430 13134 22482 13186
rect 22654 13134 22706 13186
rect 22990 13134 23042 13186
rect 29038 13134 29090 13186
rect 29486 13134 29538 13186
rect 5630 13022 5682 13074
rect 10782 13022 10834 13074
rect 12910 13022 12962 13074
rect 16382 13022 16434 13074
rect 18734 13022 18786 13074
rect 20862 13022 20914 13074
rect 21422 13022 21474 13074
rect 21982 13022 22034 13074
rect 22318 13022 22370 13074
rect 23550 13022 23602 13074
rect 26462 13022 26514 13074
rect 28030 13022 28082 13074
rect 29710 13022 29762 13074
rect 30718 13022 30770 13074
rect 32398 13022 32450 13074
rect 8542 12910 8594 12962
rect 9998 12910 10050 12962
rect 13582 12910 13634 12962
rect 17166 12910 17218 12962
rect 18286 12910 18338 12962
rect 18622 12910 18674 12962
rect 19070 12910 19122 12962
rect 21310 12910 21362 12962
rect 23102 12910 23154 12962
rect 23326 12910 23378 12962
rect 23774 12910 23826 12962
rect 23998 12910 24050 12962
rect 24558 12910 24610 12962
rect 24894 12910 24946 12962
rect 25678 12910 25730 12962
rect 28478 12910 28530 12962
rect 30158 12910 30210 12962
rect 31054 12910 31106 12962
rect 32734 12910 32786 12962
rect 7758 12798 7810 12850
rect 14254 12798 14306 12850
rect 18062 12798 18114 12850
rect 25230 12798 25282 12850
rect 26574 12798 26626 12850
rect 26910 12798 26962 12850
rect 29262 12798 29314 12850
rect 31278 12798 31330 12850
rect 31726 12798 31778 12850
rect 25902 12686 25954 12738
rect 26350 12686 26402 12738
rect 27246 12686 27298 12738
rect 27694 12686 27746 12738
rect 9278 12518 9330 12570
rect 9382 12518 9434 12570
rect 9486 12518 9538 12570
rect 17342 12518 17394 12570
rect 17446 12518 17498 12570
rect 17550 12518 17602 12570
rect 25406 12518 25458 12570
rect 25510 12518 25562 12570
rect 25614 12518 25666 12570
rect 33470 12518 33522 12570
rect 33574 12518 33626 12570
rect 33678 12518 33730 12570
rect 12238 12350 12290 12402
rect 14590 12350 14642 12402
rect 22542 12350 22594 12402
rect 23214 12350 23266 12402
rect 23886 12350 23938 12402
rect 33070 12350 33122 12402
rect 7534 12238 7586 12290
rect 12574 12238 12626 12290
rect 13358 12238 13410 12290
rect 13694 12238 13746 12290
rect 14030 12238 14082 12290
rect 14926 12238 14978 12290
rect 23550 12238 23602 12290
rect 24222 12238 24274 12290
rect 7310 12126 7362 12178
rect 7646 12126 7698 12178
rect 12014 12126 12066 12178
rect 12798 12126 12850 12178
rect 19630 12126 19682 12178
rect 20190 12126 20242 12178
rect 25342 12126 25394 12178
rect 28590 12126 28642 12178
rect 28926 12126 28978 12178
rect 29150 12126 29202 12178
rect 32398 12126 32450 12178
rect 33182 12126 33234 12178
rect 8094 12014 8146 12066
rect 8542 12014 8594 12066
rect 24670 12014 24722 12066
rect 26126 12014 26178 12066
rect 28254 12014 28306 12066
rect 29038 12014 29090 12066
rect 29598 12014 29650 12066
rect 31726 12014 31778 12066
rect 5246 11734 5298 11786
rect 5350 11734 5402 11786
rect 5454 11734 5506 11786
rect 13310 11734 13362 11786
rect 13414 11734 13466 11786
rect 13518 11734 13570 11786
rect 21374 11734 21426 11786
rect 21478 11734 21530 11786
rect 21582 11734 21634 11786
rect 29438 11734 29490 11786
rect 29542 11734 29594 11786
rect 29646 11734 29698 11786
rect 8990 11454 9042 11506
rect 9438 11454 9490 11506
rect 11454 11454 11506 11506
rect 12574 11454 12626 11506
rect 17838 11454 17890 11506
rect 19966 11454 20018 11506
rect 32062 11454 32114 11506
rect 33182 11454 33234 11506
rect 6190 11342 6242 11394
rect 10446 11342 10498 11394
rect 13470 11342 13522 11394
rect 17054 11342 17106 11394
rect 21534 11342 21586 11394
rect 27134 11342 27186 11394
rect 29262 11342 29314 11394
rect 32622 11342 32674 11394
rect 6862 11230 6914 11282
rect 25006 11230 25058 11282
rect 28590 11230 28642 11282
rect 29934 11230 29986 11282
rect 32398 11230 32450 11282
rect 9886 11118 9938 11170
rect 10894 11118 10946 11170
rect 13806 11118 13858 11170
rect 14254 11118 14306 11170
rect 14814 11118 14866 11170
rect 21870 11118 21922 11170
rect 22318 11118 22370 11170
rect 28254 11118 28306 11170
rect 9278 10950 9330 11002
rect 9382 10950 9434 11002
rect 9486 10950 9538 11002
rect 17342 10950 17394 11002
rect 17446 10950 17498 11002
rect 17550 10950 17602 11002
rect 25406 10950 25458 11002
rect 25510 10950 25562 11002
rect 25614 10950 25666 11002
rect 33470 10950 33522 11002
rect 33574 10950 33626 11002
rect 33678 10950 33730 11002
rect 4510 10782 4562 10834
rect 5406 10782 5458 10834
rect 5966 10782 6018 10834
rect 6414 10782 6466 10834
rect 6862 10782 6914 10834
rect 7758 10782 7810 10834
rect 7870 10782 7922 10834
rect 8654 10782 8706 10834
rect 11566 10782 11618 10834
rect 19742 10782 19794 10834
rect 20190 10782 20242 10834
rect 21310 10782 21362 10834
rect 26238 10782 26290 10834
rect 33182 10782 33234 10834
rect 3614 10670 3666 10722
rect 6750 10670 6802 10722
rect 7310 10670 7362 10722
rect 9662 10670 9714 10722
rect 11006 10670 11058 10722
rect 11902 10670 11954 10722
rect 19406 10670 19458 10722
rect 20974 10670 21026 10722
rect 25678 10670 25730 10722
rect 26462 10670 26514 10722
rect 3390 10558 3442 10610
rect 3726 10558 3778 10610
rect 5518 10558 5570 10610
rect 6974 10558 7026 10610
rect 7646 10558 7698 10610
rect 8206 10558 8258 10610
rect 10558 10558 10610 10610
rect 11230 10558 11282 10610
rect 12238 10558 12290 10610
rect 15598 10558 15650 10610
rect 15710 10558 15762 10610
rect 16158 10558 16210 10610
rect 17278 10558 17330 10610
rect 17614 10558 17666 10610
rect 17838 10558 17890 10610
rect 19966 10558 20018 10610
rect 20302 10558 20354 10610
rect 20526 10558 20578 10610
rect 21870 10558 21922 10610
rect 25230 10558 25282 10610
rect 25454 10558 25506 10610
rect 26126 10558 26178 10610
rect 26686 10558 26738 10610
rect 27134 10558 27186 10610
rect 4846 10446 4898 10498
rect 10446 10446 10498 10498
rect 10782 10446 10834 10498
rect 13022 10446 13074 10498
rect 15150 10446 15202 10498
rect 15934 10446 15986 10498
rect 17502 10446 17554 10498
rect 22542 10446 22594 10498
rect 24670 10446 24722 10498
rect 25342 10446 25394 10498
rect 31726 10446 31778 10498
rect 5406 10334 5458 10386
rect 5742 10334 5794 10386
rect 6526 10334 6578 10386
rect 5246 10166 5298 10218
rect 5350 10166 5402 10218
rect 5454 10166 5506 10218
rect 13310 10166 13362 10218
rect 13414 10166 13466 10218
rect 13518 10166 13570 10218
rect 21374 10166 21426 10218
rect 21478 10166 21530 10218
rect 21582 10166 21634 10218
rect 29438 10166 29490 10218
rect 29542 10166 29594 10218
rect 29646 10166 29698 10218
rect 8766 9998 8818 10050
rect 5070 9886 5122 9938
rect 9998 9886 10050 9938
rect 12126 9886 12178 9938
rect 12574 9886 12626 9938
rect 13918 9886 13970 9938
rect 15150 9886 15202 9938
rect 15710 9886 15762 9938
rect 17278 9886 17330 9938
rect 19406 9886 19458 9938
rect 20078 9886 20130 9938
rect 22206 9886 22258 9938
rect 23438 9886 23490 9938
rect 26238 9886 26290 9938
rect 27134 9886 27186 9938
rect 28366 9886 28418 9938
rect 30270 9886 30322 9938
rect 2830 9774 2882 9826
rect 3166 9774 3218 9826
rect 3390 9774 3442 9826
rect 3726 9774 3778 9826
rect 4174 9774 4226 9826
rect 4734 9774 4786 9826
rect 5742 9774 5794 9826
rect 6414 9774 6466 9826
rect 7086 9774 7138 9826
rect 9214 9774 9266 9826
rect 14142 9774 14194 9826
rect 14366 9774 14418 9826
rect 16270 9774 16322 9826
rect 16606 9774 16658 9826
rect 19966 9774 20018 9826
rect 20638 9774 20690 9826
rect 22542 9774 22594 9826
rect 23550 9774 23602 9826
rect 23886 9774 23938 9826
rect 24446 9774 24498 9826
rect 24782 9774 24834 9826
rect 25454 9774 25506 9826
rect 26350 9774 26402 9826
rect 26798 9774 26850 9826
rect 27022 9774 27074 9826
rect 27246 9774 27298 9826
rect 28030 9774 28082 9826
rect 28142 9774 28194 9826
rect 28590 9774 28642 9826
rect 29150 9774 29202 9826
rect 33070 9774 33122 9826
rect 6750 9662 6802 9714
rect 7422 9662 7474 9714
rect 7646 9662 7698 9714
rect 8318 9662 8370 9714
rect 8654 9662 8706 9714
rect 13806 9662 13858 9714
rect 20190 9662 20242 9714
rect 23326 9662 23378 9714
rect 24334 9662 24386 9714
rect 25230 9662 25282 9714
rect 25790 9662 25842 9714
rect 29262 9662 29314 9714
rect 32398 9662 32450 9714
rect 2494 9550 2546 9602
rect 2718 9550 2770 9602
rect 3390 9550 3442 9602
rect 4062 9550 4114 9602
rect 4286 9550 4338 9602
rect 6078 9550 6130 9602
rect 7310 9550 7362 9602
rect 7982 9550 8034 9602
rect 8766 9550 8818 9602
rect 14814 9550 14866 9602
rect 15038 9550 15090 9602
rect 15262 9550 15314 9602
rect 15598 9550 15650 9602
rect 15822 9550 15874 9602
rect 22878 9550 22930 9602
rect 24222 9550 24274 9602
rect 25678 9550 25730 9602
rect 26126 9550 26178 9602
rect 27470 9550 27522 9602
rect 29374 9550 29426 9602
rect 29598 9550 29650 9602
rect 9278 9382 9330 9434
rect 9382 9382 9434 9434
rect 9486 9382 9538 9434
rect 17342 9382 17394 9434
rect 17446 9382 17498 9434
rect 17550 9382 17602 9434
rect 25406 9382 25458 9434
rect 25510 9382 25562 9434
rect 25614 9382 25666 9434
rect 33470 9382 33522 9434
rect 33574 9382 33626 9434
rect 33678 9382 33730 9434
rect 4958 9214 5010 9266
rect 9662 9214 9714 9266
rect 10670 9214 10722 9266
rect 11454 9214 11506 9266
rect 13134 9214 13186 9266
rect 17502 9214 17554 9266
rect 17838 9214 17890 9266
rect 17950 9214 18002 9266
rect 18174 9214 18226 9266
rect 22318 9214 22370 9266
rect 25566 9214 25618 9266
rect 29262 9214 29314 9266
rect 29374 9214 29426 9266
rect 30270 9214 30322 9266
rect 31278 9214 31330 9266
rect 31390 9214 31442 9266
rect 32286 9214 32338 9266
rect 33294 9214 33346 9266
rect 3838 9102 3890 9154
rect 8094 9102 8146 9154
rect 10222 9102 10274 9154
rect 12350 9102 12402 9154
rect 14478 9102 14530 9154
rect 18398 9102 18450 9154
rect 19742 9102 19794 9154
rect 23550 9102 23602 9154
rect 24558 9102 24610 9154
rect 25230 9102 25282 9154
rect 26686 9102 26738 9154
rect 29150 9102 29202 9154
rect 31838 9102 31890 9154
rect 4622 8990 4674 9042
rect 5182 8990 5234 9042
rect 5518 8990 5570 9042
rect 8878 8990 8930 9042
rect 9774 8990 9826 9042
rect 10110 8990 10162 9042
rect 10446 8990 10498 9042
rect 10894 8990 10946 9042
rect 11342 8990 11394 9042
rect 11566 8990 11618 9042
rect 11902 8990 11954 9042
rect 12126 8990 12178 9042
rect 12462 8990 12514 9042
rect 13694 8990 13746 9042
rect 17726 8990 17778 9042
rect 18510 8990 18562 9042
rect 19070 8990 19122 9042
rect 23774 8990 23826 9042
rect 24334 8990 24386 9042
rect 26014 8990 26066 9042
rect 29822 8990 29874 9042
rect 30606 8990 30658 9042
rect 30942 8990 30994 9042
rect 31502 8990 31554 9042
rect 32062 8990 32114 9042
rect 32398 8990 32450 9042
rect 1710 8878 1762 8930
rect 5070 8878 5122 8930
rect 5966 8878 6018 8930
rect 16606 8878 16658 8930
rect 21870 8878 21922 8930
rect 22878 8878 22930 8930
rect 23214 8878 23266 8930
rect 28814 8878 28866 8930
rect 9662 8766 9714 8818
rect 5246 8598 5298 8650
rect 5350 8598 5402 8650
rect 5454 8598 5506 8650
rect 13310 8598 13362 8650
rect 13414 8598 13466 8650
rect 13518 8598 13570 8650
rect 21374 8598 21426 8650
rect 21478 8598 21530 8650
rect 21582 8598 21634 8650
rect 29438 8598 29490 8650
rect 29542 8598 29594 8650
rect 29646 8598 29698 8650
rect 21982 8430 22034 8482
rect 22766 8430 22818 8482
rect 24782 8430 24834 8482
rect 4622 8318 4674 8370
rect 5854 8318 5906 8370
rect 8878 8318 8930 8370
rect 22318 8318 22370 8370
rect 25342 8318 25394 8370
rect 30046 8318 30098 8370
rect 30270 8318 30322 8370
rect 1822 8206 1874 8258
rect 5966 8206 6018 8258
rect 11678 8206 11730 8258
rect 12574 8206 12626 8258
rect 14926 8206 14978 8258
rect 19630 8206 19682 8258
rect 23214 8206 23266 8258
rect 23774 8206 23826 8258
rect 24334 8206 24386 8258
rect 26238 8206 26290 8258
rect 28030 8206 28082 8258
rect 28142 8206 28194 8258
rect 28254 8206 28306 8258
rect 28702 8206 28754 8258
rect 33070 8206 33122 8258
rect 2494 8094 2546 8146
rect 5742 8094 5794 8146
rect 6302 8094 6354 8146
rect 17838 8094 17890 8146
rect 20302 8094 20354 8146
rect 21870 8094 21922 8146
rect 24670 8094 24722 8146
rect 27246 8094 27298 8146
rect 27694 8094 27746 8146
rect 29486 8094 29538 8146
rect 32398 8094 32450 8146
rect 5182 7982 5234 8034
rect 12910 7982 12962 8034
rect 19406 7982 19458 8034
rect 19518 7982 19570 8034
rect 19854 7982 19906 8034
rect 20638 7982 20690 8034
rect 22766 7982 22818 8034
rect 22878 7982 22930 8034
rect 23102 7982 23154 8034
rect 23438 7982 23490 8034
rect 23662 7982 23714 8034
rect 23998 7982 24050 8034
rect 24222 7982 24274 8034
rect 24782 7982 24834 8034
rect 25902 7982 25954 8034
rect 26798 7982 26850 8034
rect 27358 7982 27410 8034
rect 27582 7982 27634 8034
rect 29150 7982 29202 8034
rect 9278 7814 9330 7866
rect 9382 7814 9434 7866
rect 9486 7814 9538 7866
rect 17342 7814 17394 7866
rect 17446 7814 17498 7866
rect 17550 7814 17602 7866
rect 25406 7814 25458 7866
rect 25510 7814 25562 7866
rect 25614 7814 25666 7866
rect 33470 7814 33522 7866
rect 33574 7814 33626 7866
rect 33678 7814 33730 7866
rect 3054 7646 3106 7698
rect 4174 7646 4226 7698
rect 4398 7646 4450 7698
rect 5854 7646 5906 7698
rect 7758 7646 7810 7698
rect 7870 7646 7922 7698
rect 13246 7646 13298 7698
rect 17502 7646 17554 7698
rect 17614 7646 17666 7698
rect 19854 7646 19906 7698
rect 20302 7646 20354 7698
rect 21646 7646 21698 7698
rect 23326 7646 23378 7698
rect 24670 7646 24722 7698
rect 27470 7646 27522 7698
rect 28366 7646 28418 7698
rect 29598 7646 29650 7698
rect 30046 7646 30098 7698
rect 31054 7646 31106 7698
rect 32062 7646 32114 7698
rect 33182 7646 33234 7698
rect 2494 7534 2546 7586
rect 3278 7534 3330 7586
rect 3502 7534 3554 7586
rect 4958 7534 5010 7586
rect 5966 7534 6018 7586
rect 8542 7534 8594 7586
rect 16718 7534 16770 7586
rect 19294 7534 19346 7586
rect 21758 7534 21810 7586
rect 22094 7534 22146 7586
rect 25566 7534 25618 7586
rect 26686 7534 26738 7586
rect 27806 7534 27858 7586
rect 28590 7534 28642 7586
rect 28926 7534 28978 7586
rect 29374 7534 29426 7586
rect 30382 7534 30434 7586
rect 2046 7422 2098 7474
rect 2382 7422 2434 7474
rect 2606 7422 2658 7474
rect 2830 7422 2882 7474
rect 3838 7422 3890 7474
rect 4286 7422 4338 7474
rect 4846 7422 4898 7474
rect 5406 7422 5458 7474
rect 5630 7422 5682 7474
rect 6078 7422 6130 7474
rect 6750 7422 6802 7474
rect 6974 7422 7026 7474
rect 7422 7422 7474 7474
rect 7646 7422 7698 7474
rect 8206 7422 8258 7474
rect 8766 7422 8818 7474
rect 12350 7422 12402 7474
rect 13134 7422 13186 7474
rect 13694 7422 13746 7474
rect 16606 7422 16658 7474
rect 16942 7422 16994 7474
rect 17390 7422 17442 7474
rect 18062 7422 18114 7474
rect 18286 7422 18338 7474
rect 18622 7422 18674 7474
rect 18846 7422 18898 7474
rect 19406 7422 19458 7474
rect 22318 7422 22370 7474
rect 22766 7422 22818 7474
rect 23102 7422 23154 7474
rect 23438 7422 23490 7474
rect 25230 7422 25282 7474
rect 27022 7422 27074 7474
rect 29262 7422 29314 7474
rect 30606 7422 30658 7474
rect 31278 7422 31330 7474
rect 31614 7422 31666 7474
rect 31950 7422 32002 7474
rect 32174 7422 32226 7474
rect 5182 7310 5234 7362
rect 6862 7310 6914 7362
rect 9550 7310 9602 7362
rect 11678 7310 11730 7362
rect 14926 7310 14978 7362
rect 18734 7310 18786 7362
rect 21310 7310 21362 7362
rect 22206 7310 22258 7362
rect 24334 7310 24386 7362
rect 26462 7310 26514 7362
rect 31166 7310 31218 7362
rect 13246 7198 13298 7250
rect 19294 7198 19346 7250
rect 21646 7198 21698 7250
rect 5246 7030 5298 7082
rect 5350 7030 5402 7082
rect 5454 7030 5506 7082
rect 13310 7030 13362 7082
rect 13414 7030 13466 7082
rect 13518 7030 13570 7082
rect 21374 7030 21426 7082
rect 21478 7030 21530 7082
rect 21582 7030 21634 7082
rect 29438 7030 29490 7082
rect 29542 7030 29594 7082
rect 29646 7030 29698 7082
rect 10894 6750 10946 6802
rect 16494 6750 16546 6802
rect 16942 6750 16994 6802
rect 20750 6750 20802 6802
rect 23550 6750 23602 6802
rect 31502 6750 31554 6802
rect 4062 6638 4114 6690
rect 4846 6638 4898 6690
rect 5854 6638 5906 6690
rect 9662 6638 9714 6690
rect 10670 6638 10722 6690
rect 11342 6638 11394 6690
rect 11902 6638 11954 6690
rect 12462 6638 12514 6690
rect 12910 6638 12962 6690
rect 13582 6638 13634 6690
rect 17054 6638 17106 6690
rect 17838 6638 17890 6690
rect 21646 6638 21698 6690
rect 22430 6638 22482 6690
rect 22766 6638 22818 6690
rect 23102 6638 23154 6690
rect 24110 6638 24162 6690
rect 24558 6638 24610 6690
rect 25678 6638 25730 6690
rect 26350 6638 26402 6690
rect 27134 6638 27186 6690
rect 28366 6638 28418 6690
rect 28702 6638 28754 6690
rect 30046 6638 30098 6690
rect 30606 6638 30658 6690
rect 30718 6638 30770 6690
rect 31390 6638 31442 6690
rect 32510 6638 32562 6690
rect 33182 6638 33234 6690
rect 9438 6526 9490 6578
rect 10222 6526 10274 6578
rect 10334 6526 10386 6578
rect 11118 6526 11170 6578
rect 11790 6526 11842 6578
rect 12798 6526 12850 6578
rect 14366 6526 14418 6578
rect 18622 6526 18674 6578
rect 21982 6526 22034 6578
rect 22206 6526 22258 6578
rect 24446 6526 24498 6578
rect 26798 6526 26850 6578
rect 27470 6526 27522 6578
rect 27806 6526 27858 6578
rect 29486 6526 29538 6578
rect 29822 6526 29874 6578
rect 31614 6526 31666 6578
rect 32174 6526 32226 6578
rect 32846 6526 32898 6578
rect 3278 6414 3330 6466
rect 5070 6414 5122 6466
rect 6862 6414 6914 6466
rect 8766 6414 8818 6466
rect 9102 6414 9154 6466
rect 10558 6414 10610 6466
rect 11566 6414 11618 6466
rect 12574 6414 12626 6466
rect 16830 6414 16882 6466
rect 17278 6414 17330 6466
rect 21758 6414 21810 6466
rect 22654 6414 22706 6466
rect 23438 6414 23490 6466
rect 23662 6414 23714 6466
rect 24222 6414 24274 6466
rect 25118 6414 25170 6466
rect 25342 6414 25394 6466
rect 26014 6414 26066 6466
rect 28478 6414 28530 6466
rect 30494 6414 30546 6466
rect 31166 6414 31218 6466
rect 9278 6246 9330 6298
rect 9382 6246 9434 6298
rect 9486 6246 9538 6298
rect 17342 6246 17394 6298
rect 17446 6246 17498 6298
rect 17550 6246 17602 6298
rect 25406 6246 25458 6298
rect 25510 6246 25562 6298
rect 25614 6246 25666 6298
rect 33470 6246 33522 6298
rect 33574 6246 33626 6298
rect 33678 6246 33730 6298
rect 5294 6078 5346 6130
rect 22206 6078 22258 6130
rect 22318 6078 22370 6130
rect 22430 6078 22482 6130
rect 23550 6078 23602 6130
rect 24110 6078 24162 6130
rect 26126 6078 26178 6130
rect 27358 6078 27410 6130
rect 28254 6078 28306 6130
rect 29150 6078 29202 6130
rect 29374 6078 29426 6130
rect 29598 6078 29650 6130
rect 31726 6078 31778 6130
rect 31950 6078 32002 6130
rect 33070 6078 33122 6130
rect 3838 5966 3890 6018
rect 5070 5966 5122 6018
rect 8094 5966 8146 6018
rect 9662 5966 9714 6018
rect 9774 5966 9826 6018
rect 10446 5966 10498 6018
rect 10782 5966 10834 6018
rect 11006 5966 11058 6018
rect 17726 5966 17778 6018
rect 17950 5966 18002 6018
rect 19742 5966 19794 6018
rect 24558 5966 24610 6018
rect 25566 5966 25618 6018
rect 27246 5966 27298 6018
rect 27918 5966 27970 6018
rect 28030 5966 28082 6018
rect 28478 5966 28530 6018
rect 28590 5966 28642 6018
rect 29038 5966 29090 6018
rect 29822 5966 29874 6018
rect 31054 5966 31106 6018
rect 4510 5854 4562 5906
rect 5406 5854 5458 5906
rect 5518 5854 5570 5906
rect 8878 5854 8930 5906
rect 11790 5854 11842 5906
rect 14254 5854 14306 5906
rect 17278 5854 17330 5906
rect 17502 5854 17554 5906
rect 19070 5854 19122 5906
rect 22766 5854 22818 5906
rect 23102 5854 23154 5906
rect 23326 5854 23378 5906
rect 24334 5854 24386 5906
rect 25230 5854 25282 5906
rect 25342 5854 25394 5906
rect 25790 5854 25842 5906
rect 26238 5854 26290 5906
rect 26350 5854 26402 5906
rect 26686 5854 26738 5906
rect 27582 5854 27634 5906
rect 28814 5854 28866 5906
rect 30158 5854 30210 5906
rect 30382 5854 30434 5906
rect 30830 5854 30882 5906
rect 31278 5854 31330 5906
rect 1710 5742 1762 5794
rect 5966 5742 6018 5794
rect 10558 5742 10610 5794
rect 18398 5742 18450 5794
rect 21870 5742 21922 5794
rect 23214 5742 23266 5794
rect 24446 5742 24498 5794
rect 29710 5742 29762 5794
rect 30942 5742 30994 5794
rect 31838 5742 31890 5794
rect 32398 5742 32450 5794
rect 33182 5742 33234 5794
rect 9774 5630 9826 5682
rect 12350 5630 12402 5682
rect 15262 5630 15314 5682
rect 32286 5630 32338 5682
rect 5246 5462 5298 5514
rect 5350 5462 5402 5514
rect 5454 5462 5506 5514
rect 13310 5462 13362 5514
rect 13414 5462 13466 5514
rect 13518 5462 13570 5514
rect 21374 5462 21426 5514
rect 21478 5462 21530 5514
rect 21582 5462 21634 5514
rect 29438 5462 29490 5514
rect 29542 5462 29594 5514
rect 29646 5462 29698 5514
rect 26798 5294 26850 5346
rect 2718 5182 2770 5234
rect 9774 5182 9826 5234
rect 11902 5182 11954 5234
rect 18734 5182 18786 5234
rect 20302 5182 20354 5234
rect 20750 5182 20802 5234
rect 22542 5182 22594 5234
rect 24558 5182 24610 5234
rect 25454 5182 25506 5234
rect 28478 5182 28530 5234
rect 30270 5182 30322 5234
rect 2270 5070 2322 5122
rect 4622 5070 4674 5122
rect 5854 5070 5906 5122
rect 8430 5070 8482 5122
rect 8990 5070 9042 5122
rect 12126 5070 12178 5122
rect 12350 5070 12402 5122
rect 12574 5070 12626 5122
rect 12798 5070 12850 5122
rect 13918 5070 13970 5122
rect 14142 5070 14194 5122
rect 14478 5070 14530 5122
rect 14814 5070 14866 5122
rect 15374 5070 15426 5122
rect 15822 5070 15874 5122
rect 18958 5070 19010 5122
rect 19966 5070 20018 5122
rect 21534 5070 21586 5122
rect 24334 5070 24386 5122
rect 24782 5070 24834 5122
rect 24894 5070 24946 5122
rect 25342 5070 25394 5122
rect 26014 5070 26066 5122
rect 26126 5070 26178 5122
rect 26462 5070 26514 5122
rect 27582 5070 27634 5122
rect 28030 5070 28082 5122
rect 28142 5070 28194 5122
rect 29038 5070 29090 5122
rect 29374 5070 29426 5122
rect 29710 5070 29762 5122
rect 32398 5070 32450 5122
rect 33070 5070 33122 5122
rect 1934 4958 1986 5010
rect 2046 4958 2098 5010
rect 7086 4958 7138 5010
rect 13582 4958 13634 5010
rect 15150 4958 15202 5010
rect 16606 4958 16658 5010
rect 19294 4958 19346 5010
rect 19630 4958 19682 5010
rect 26350 4958 26402 5010
rect 26910 4958 26962 5010
rect 27918 4958 27970 5010
rect 28590 4958 28642 5010
rect 14478 4846 14530 4898
rect 19182 4846 19234 4898
rect 19742 4846 19794 4898
rect 25566 4846 25618 4898
rect 29262 4846 29314 4898
rect 9278 4678 9330 4730
rect 9382 4678 9434 4730
rect 9486 4678 9538 4730
rect 17342 4678 17394 4730
rect 17446 4678 17498 4730
rect 17550 4678 17602 4730
rect 25406 4678 25458 4730
rect 25510 4678 25562 4730
rect 25614 4678 25666 4730
rect 33470 4678 33522 4730
rect 33574 4678 33626 4730
rect 33678 4678 33730 4730
rect 8206 4510 8258 4562
rect 8318 4510 8370 4562
rect 16606 4510 16658 4562
rect 24110 4510 24162 4562
rect 31838 4510 31890 4562
rect 33070 4510 33122 4562
rect 3838 4398 3890 4450
rect 5742 4398 5794 4450
rect 14814 4398 14866 4450
rect 18174 4398 18226 4450
rect 21646 4398 21698 4450
rect 24558 4398 24610 4450
rect 26014 4398 26066 4450
rect 29262 4398 29314 4450
rect 32062 4398 32114 4450
rect 4510 4286 4562 4338
rect 4958 4286 5010 4338
rect 8430 4286 8482 4338
rect 8766 4286 8818 4338
rect 12014 4286 12066 4338
rect 15598 4286 15650 4338
rect 16382 4286 16434 4338
rect 16606 4286 16658 4338
rect 16942 4286 16994 4338
rect 17390 4286 17442 4338
rect 20862 4286 20914 4338
rect 25342 4286 25394 4338
rect 28590 4286 28642 4338
rect 31614 4286 31666 4338
rect 32174 4286 32226 4338
rect 1710 4174 1762 4226
rect 7870 4174 7922 4226
rect 10334 4174 10386 4226
rect 12686 4174 12738 4226
rect 20302 4174 20354 4226
rect 23774 4174 23826 4226
rect 24222 4174 24274 4226
rect 24670 4174 24722 4226
rect 28142 4174 28194 4226
rect 31390 4174 31442 4226
rect 33182 4174 33234 4226
rect 5246 3894 5298 3946
rect 5350 3894 5402 3946
rect 5454 3894 5506 3946
rect 13310 3894 13362 3946
rect 13414 3894 13466 3946
rect 13518 3894 13570 3946
rect 21374 3894 21426 3946
rect 21478 3894 21530 3946
rect 21582 3894 21634 3946
rect 29438 3894 29490 3946
rect 29542 3894 29594 3946
rect 29646 3894 29698 3946
rect 26910 3726 26962 3778
rect 27918 3726 27970 3778
rect 8542 3614 8594 3666
rect 9550 3614 9602 3666
rect 11678 3614 11730 3666
rect 16158 3614 16210 3666
rect 18174 3614 18226 3666
rect 21870 3614 21922 3666
rect 25566 3614 25618 3666
rect 2382 3502 2434 3554
rect 6190 3502 6242 3554
rect 12462 3502 12514 3554
rect 13246 3502 13298 3554
rect 13582 3502 13634 3554
rect 13806 3502 13858 3554
rect 16942 3502 16994 3554
rect 17278 3502 17330 3554
rect 20078 3502 20130 3554
rect 20750 3502 20802 3554
rect 24894 3502 24946 3554
rect 26462 3502 26514 3554
rect 27022 3502 27074 3554
rect 28590 3502 28642 3554
rect 29598 3502 29650 3554
rect 30270 3502 30322 3554
rect 32286 3502 32338 3554
rect 33182 3502 33234 3554
rect 1822 3390 1874 3442
rect 4062 3390 4114 3442
rect 5742 3390 5794 3442
rect 1934 3278 1986 3330
rect 2158 3278 2210 3330
rect 5518 3278 5570 3330
rect 5854 3334 5906 3386
rect 13358 3390 13410 3442
rect 17166 3390 17218 3442
rect 23662 3390 23714 3442
rect 23998 3390 24050 3442
rect 24670 3390 24722 3442
rect 25902 3390 25954 3442
rect 26238 3390 26290 3442
rect 27470 3390 27522 3442
rect 28366 3390 28418 3442
rect 29374 3390 29426 3442
rect 30606 3390 30658 3442
rect 30942 3390 30994 3442
rect 31278 3390 31330 3442
rect 32510 3390 32562 3442
rect 32846 3390 32898 3442
rect 9278 3110 9330 3162
rect 9382 3110 9434 3162
rect 9486 3110 9538 3162
rect 17342 3110 17394 3162
rect 17446 3110 17498 3162
rect 17550 3110 17602 3162
rect 25406 3110 25458 3162
rect 25510 3110 25562 3162
rect 25614 3110 25666 3162
rect 33470 3110 33522 3162
rect 33574 3110 33626 3162
rect 33678 3110 33730 3162
<< metal2 >>
rect 448 34200 560 35000
rect 1568 34200 1680 35000
rect 2688 34200 2800 35000
rect 3808 34200 3920 35000
rect 4928 34200 5040 35000
rect 6048 34200 6160 35000
rect 7168 34200 7280 35000
rect 8288 34200 8400 35000
rect 9408 34200 9520 35000
rect 10528 34200 10640 35000
rect 10892 34300 11284 34356
rect 476 31554 532 34200
rect 1596 31948 1652 34200
rect 2716 31948 2772 34200
rect 1596 31892 1876 31948
rect 2716 31892 2996 31948
rect 476 31502 478 31554
rect 530 31502 532 31554
rect 476 31490 532 31502
rect 1820 31218 1876 31892
rect 1820 31166 1822 31218
rect 1874 31166 1876 31218
rect 1820 31154 1876 31166
rect 2268 31554 2324 31566
rect 2268 31502 2270 31554
rect 2322 31502 2324 31554
rect 2268 31218 2324 31502
rect 2268 31166 2270 31218
rect 2322 31166 2324 31218
rect 2268 31154 2324 31166
rect 2940 31218 2996 31892
rect 2940 31166 2942 31218
rect 2994 31166 2996 31218
rect 2940 31154 2996 31166
rect 3836 31220 3892 34200
rect 4956 32788 5012 34200
rect 4508 32732 5012 32788
rect 3948 31220 4004 31230
rect 3836 31218 4004 31220
rect 3836 31166 3950 31218
rect 4002 31166 4004 31218
rect 3836 31164 4004 31166
rect 3948 31154 4004 31164
rect 4508 31218 4564 32732
rect 4508 31166 4510 31218
rect 4562 31166 4564 31218
rect 4508 31154 4564 31166
rect 4956 31892 5012 31902
rect 4956 31218 5012 31836
rect 6076 31892 6132 34200
rect 6076 31826 6132 31836
rect 6860 31780 6916 31790
rect 4956 31166 4958 31218
rect 5010 31166 5012 31218
rect 4956 31154 5012 31166
rect 5068 31556 5124 31566
rect 3724 31108 3780 31118
rect 3724 31014 3780 31052
rect 5068 30548 5124 31500
rect 5852 31220 5908 31230
rect 5852 31126 5908 31164
rect 6636 30994 6692 31006
rect 6636 30942 6638 30994
rect 6690 30942 6692 30994
rect 4956 30492 5124 30548
rect 5244 30604 5508 30614
rect 5300 30548 5348 30604
rect 5404 30548 5452 30604
rect 5244 30538 5508 30548
rect 2268 30210 2324 30222
rect 2268 30158 2270 30210
rect 2322 30158 2324 30210
rect 1708 29316 1764 29326
rect 1708 28642 1764 29260
rect 2268 29316 2324 30158
rect 2940 30100 2996 30110
rect 2940 30006 2996 30044
rect 3948 30100 4004 30110
rect 4956 30100 5012 30492
rect 5068 30324 5124 30334
rect 5068 30322 5236 30324
rect 5068 30270 5070 30322
rect 5122 30270 5236 30322
rect 5068 30268 5236 30270
rect 5068 30258 5124 30268
rect 4956 30044 5124 30100
rect 3948 29650 4004 30044
rect 3948 29598 3950 29650
rect 4002 29598 4004 29650
rect 3948 29586 4004 29598
rect 5068 29650 5124 30044
rect 5068 29598 5070 29650
rect 5122 29598 5124 29650
rect 5068 29586 5124 29598
rect 2268 29250 2324 29260
rect 4060 29314 4116 29326
rect 4060 29262 4062 29314
rect 4114 29262 4116 29314
rect 4060 28756 4116 29262
rect 4508 29316 4564 29326
rect 5180 29316 5236 30268
rect 5628 30210 5684 30222
rect 5628 30158 5630 30210
rect 5682 30158 5684 30210
rect 5516 29652 5572 29662
rect 5516 29558 5572 29596
rect 5292 29316 5348 29326
rect 4564 29260 5012 29316
rect 5180 29260 5292 29316
rect 4508 29222 4564 29260
rect 4060 28690 4116 28700
rect 4620 29092 4676 29102
rect 4620 28754 4676 29036
rect 4620 28702 4622 28754
rect 4674 28702 4676 28754
rect 4620 28690 4676 28702
rect 4844 28868 4900 28878
rect 1708 28590 1710 28642
rect 1762 28590 1764 28642
rect 1708 27858 1764 28590
rect 2492 28532 2548 28542
rect 2492 28530 3332 28532
rect 2492 28478 2494 28530
rect 2546 28478 3332 28530
rect 2492 28476 3332 28478
rect 2492 28466 2548 28476
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 27794 1764 27806
rect 2492 27748 2548 27758
rect 2492 27746 2884 27748
rect 2492 27694 2494 27746
rect 2546 27694 2884 27746
rect 2492 27692 2884 27694
rect 2492 27682 2548 27692
rect 2828 27298 2884 27692
rect 2828 27246 2830 27298
rect 2882 27246 2884 27298
rect 2828 27234 2884 27246
rect 3276 27298 3332 28476
rect 4620 27746 4676 27758
rect 4620 27694 4622 27746
rect 4674 27694 4676 27746
rect 4620 27636 4676 27694
rect 4620 27570 4676 27580
rect 3276 27246 3278 27298
rect 3330 27246 3332 27298
rect 3276 27234 3332 27246
rect 2940 27188 2996 27198
rect 2940 27094 2996 27132
rect 4844 27074 4900 28812
rect 4956 28644 5012 29260
rect 5292 29250 5348 29260
rect 5244 29036 5508 29046
rect 5300 28980 5348 29036
rect 5404 28980 5452 29036
rect 5244 28970 5508 28980
rect 5180 28644 5236 28654
rect 4956 28588 5124 28644
rect 5068 28084 5124 28588
rect 5180 28550 5236 28588
rect 5516 28084 5572 28094
rect 5628 28084 5684 30158
rect 6412 30100 6468 30110
rect 6412 30006 6468 30044
rect 6076 29540 6132 29550
rect 6636 29540 6692 30942
rect 6860 29652 6916 31724
rect 7196 31220 7252 34200
rect 7196 31154 7252 31164
rect 7980 31892 8036 31902
rect 7980 31106 8036 31836
rect 7980 31054 7982 31106
rect 8034 31054 8036 31106
rect 7980 31042 8036 31054
rect 6860 29586 6916 29596
rect 7196 30324 7252 30334
rect 7196 29650 7252 30268
rect 7196 29598 7198 29650
rect 7250 29598 7252 29650
rect 7196 29586 7252 29598
rect 7644 30100 7700 30110
rect 6076 29538 6244 29540
rect 6076 29486 6078 29538
rect 6130 29486 6244 29538
rect 6076 29484 6244 29486
rect 6076 29474 6132 29484
rect 5852 29426 5908 29438
rect 5852 29374 5854 29426
rect 5906 29374 5908 29426
rect 5852 29204 5908 29374
rect 5852 29138 5908 29148
rect 6076 28756 6132 28766
rect 6076 28662 6132 28700
rect 5740 28418 5796 28430
rect 5740 28366 5742 28418
rect 5794 28366 5796 28418
rect 5740 28084 5796 28366
rect 5068 28082 5796 28084
rect 5068 28030 5070 28082
rect 5122 28030 5518 28082
rect 5570 28030 5796 28082
rect 5068 28028 5796 28030
rect 5068 28018 5124 28028
rect 5516 28018 5572 28028
rect 5244 27468 5508 27478
rect 5300 27412 5348 27468
rect 5404 27412 5452 27468
rect 5244 27402 5508 27412
rect 4844 27022 4846 27074
rect 4898 27022 4900 27074
rect 3388 26962 3444 26974
rect 3388 26910 3390 26962
rect 3442 26910 3444 26962
rect 3388 26068 3444 26910
rect 3388 26002 3444 26012
rect 4732 25732 4788 25742
rect 4172 25620 4228 25630
rect 4620 25620 4676 25630
rect 4172 25618 4676 25620
rect 4172 25566 4174 25618
rect 4226 25566 4622 25618
rect 4674 25566 4676 25618
rect 4172 25564 4676 25566
rect 4172 25554 4228 25564
rect 4620 25554 4676 25564
rect 4732 25506 4788 25676
rect 4732 25454 4734 25506
rect 4786 25454 4788 25506
rect 4732 25442 4788 25454
rect 2492 25284 2548 25294
rect 2492 24834 2548 25228
rect 2492 24782 2494 24834
rect 2546 24782 2548 24834
rect 2492 24770 2548 24782
rect 3948 25282 4004 25294
rect 3948 25230 3950 25282
rect 4002 25230 4004 25282
rect 1820 24722 1876 24734
rect 1820 24670 1822 24722
rect 1874 24670 1876 24722
rect 1820 23938 1876 24670
rect 3948 24052 4004 25230
rect 4060 25284 4116 25294
rect 4060 25190 4116 25228
rect 4508 25282 4564 25294
rect 4508 25230 4510 25282
rect 4562 25230 4564 25282
rect 4508 24836 4564 25230
rect 4508 24770 4564 24780
rect 4620 24612 4676 24622
rect 4620 24518 4676 24556
rect 3948 23986 4004 23996
rect 4732 24052 4788 24062
rect 4844 24052 4900 27022
rect 5180 26962 5236 26974
rect 5180 26910 5182 26962
rect 5234 26910 5236 26962
rect 4956 26850 5012 26862
rect 4956 26798 4958 26850
rect 5010 26798 5012 26850
rect 4956 26628 5012 26798
rect 4956 26562 5012 26572
rect 5068 26404 5124 26414
rect 4732 24050 4900 24052
rect 4732 23998 4734 24050
rect 4786 23998 4900 24050
rect 4732 23996 4900 23998
rect 4732 23986 4788 23996
rect 1820 23886 1822 23938
rect 1874 23886 1876 23938
rect 1820 22370 1876 23886
rect 4844 23940 4900 23996
rect 4844 23874 4900 23884
rect 4956 26292 5012 26302
rect 2492 23826 2548 23838
rect 2492 23774 2494 23826
rect 2546 23774 2548 23826
rect 2492 23380 2548 23774
rect 4956 23604 5012 26236
rect 5068 26290 5124 26348
rect 5068 26238 5070 26290
rect 5122 26238 5124 26290
rect 5068 26226 5124 26238
rect 5180 26178 5236 26910
rect 5180 26126 5182 26178
rect 5234 26126 5236 26178
rect 5180 26114 5236 26126
rect 5516 26180 5572 26190
rect 5516 26086 5572 26124
rect 5244 25900 5508 25910
rect 5300 25844 5348 25900
rect 5404 25844 5452 25900
rect 5244 25834 5508 25844
rect 2492 23314 2548 23324
rect 4732 23548 5012 23604
rect 5068 25732 5124 25742
rect 1820 22318 1822 22370
rect 1874 22318 1876 22370
rect 1820 22148 1876 22318
rect 4620 22482 4676 22494
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 1820 21586 1876 22092
rect 2492 22258 2548 22270
rect 2492 22206 2494 22258
rect 2546 22206 2548 22258
rect 2492 21812 2548 22206
rect 4620 21924 4676 22430
rect 4620 21858 4676 21868
rect 2492 21746 2548 21756
rect 1820 21534 1822 21586
rect 1874 21534 1876 21586
rect 1820 19234 1876 21534
rect 2492 21476 2548 21486
rect 2492 21382 2548 21420
rect 4172 21476 4228 21486
rect 4620 21476 4676 21486
rect 4172 20914 4228 21420
rect 4172 20862 4174 20914
rect 4226 20862 4228 20914
rect 4172 20850 4228 20862
rect 4508 21474 4676 21476
rect 4508 21422 4622 21474
rect 4674 21422 4676 21474
rect 4508 21420 4676 21422
rect 4284 20802 4340 20814
rect 4284 20750 4286 20802
rect 4338 20750 4340 20802
rect 4060 20690 4116 20702
rect 4060 20638 4062 20690
rect 4114 20638 4116 20690
rect 4060 19460 4116 20638
rect 4284 20242 4340 20750
rect 4284 20190 4286 20242
rect 4338 20190 4340 20242
rect 4284 20178 4340 20190
rect 4508 20580 4564 21420
rect 4620 21410 4676 21420
rect 4620 20804 4676 20814
rect 4620 20710 4676 20748
rect 4620 20580 4676 20590
rect 4508 20524 4620 20580
rect 4508 20242 4564 20524
rect 4620 20514 4676 20524
rect 4508 20190 4510 20242
rect 4562 20190 4564 20242
rect 4508 20178 4564 20190
rect 4620 20020 4676 20030
rect 4620 19926 4676 19964
rect 4060 19394 4116 19404
rect 4620 19348 4676 19358
rect 1820 19182 1822 19234
rect 1874 19182 1876 19234
rect 1820 17666 1876 19182
rect 4508 19346 4676 19348
rect 4508 19294 4622 19346
rect 4674 19294 4676 19346
rect 4508 19292 4676 19294
rect 2492 19122 2548 19134
rect 2492 19070 2494 19122
rect 2546 19070 2548 19122
rect 2492 18340 2548 19070
rect 3612 19124 3668 19134
rect 3612 18788 3668 19068
rect 4508 19012 4564 19292
rect 4620 19282 4676 19292
rect 4508 18946 4564 18956
rect 4620 19124 4676 19134
rect 3052 18676 3108 18686
rect 3052 18582 3108 18620
rect 3612 18674 3668 18732
rect 3612 18622 3614 18674
rect 3666 18622 3668 18674
rect 3612 18610 3668 18622
rect 3724 18676 3780 18686
rect 2940 18562 2996 18574
rect 2940 18510 2942 18562
rect 2994 18510 2996 18562
rect 2940 18340 2996 18510
rect 3724 18562 3780 18620
rect 3724 18510 3726 18562
rect 3778 18510 3780 18562
rect 3724 18498 3780 18510
rect 3276 18452 3332 18462
rect 3276 18358 3332 18396
rect 3948 18452 4004 18462
rect 3948 18358 4004 18396
rect 4396 18452 4452 18462
rect 4396 18358 4452 18396
rect 4508 18450 4564 18462
rect 4508 18398 4510 18450
rect 4562 18398 4564 18450
rect 4172 18340 4228 18350
rect 2940 18284 3220 18340
rect 2492 18274 2548 18284
rect 3164 18228 3220 18284
rect 4172 18246 4228 18284
rect 3500 18228 3556 18238
rect 3164 18172 3500 18228
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1820 15314 1876 17614
rect 2492 17556 2548 17566
rect 3500 17556 3556 18172
rect 3612 18228 3668 18238
rect 3612 18226 4116 18228
rect 3612 18174 3614 18226
rect 3666 18174 4116 18226
rect 3612 18172 4116 18174
rect 3612 18162 3668 18172
rect 3948 17780 4004 17790
rect 3500 17500 3892 17556
rect 2492 17462 2548 17500
rect 3836 16098 3892 17500
rect 3948 16996 4004 17724
rect 4060 17444 4116 18172
rect 4508 17780 4564 18398
rect 4508 17714 4564 17724
rect 4620 17778 4676 19068
rect 4620 17726 4622 17778
rect 4674 17726 4676 17778
rect 4620 17714 4676 17726
rect 4508 17556 4564 17566
rect 4060 17388 4452 17444
rect 4172 16996 4228 17006
rect 3948 16994 4228 16996
rect 3948 16942 4174 16994
rect 4226 16942 4228 16994
rect 3948 16940 4228 16942
rect 4172 16660 4228 16940
rect 4396 16994 4452 17388
rect 4508 17106 4564 17500
rect 4508 17054 4510 17106
rect 4562 17054 4564 17106
rect 4508 17042 4564 17054
rect 4732 17108 4788 23548
rect 4956 23380 5012 23390
rect 4844 23324 4956 23380
rect 4844 23266 4900 23324
rect 4844 23214 4846 23266
rect 4898 23214 4900 23266
rect 4844 23202 4900 23214
rect 4956 22484 5012 23324
rect 5068 23268 5124 25676
rect 5740 25618 5796 28028
rect 6188 27860 6244 29484
rect 6524 29316 6580 29326
rect 6524 28980 6580 29260
rect 6300 28644 6356 28654
rect 6300 28530 6356 28588
rect 6300 28478 6302 28530
rect 6354 28478 6356 28530
rect 6300 28084 6356 28478
rect 6300 28018 6356 28028
rect 6412 28642 6468 28654
rect 6412 28590 6414 28642
rect 6466 28590 6468 28642
rect 6300 27860 6356 27870
rect 6188 27804 6300 27860
rect 6300 27766 6356 27804
rect 6188 27524 6244 27534
rect 5964 26964 6020 27002
rect 5964 26898 6020 26908
rect 6076 26962 6132 26974
rect 6076 26910 6078 26962
rect 6130 26910 6132 26962
rect 6076 25844 6132 26910
rect 6188 26962 6244 27468
rect 6300 27188 6356 27198
rect 6412 27188 6468 28590
rect 6524 28532 6580 28924
rect 6636 28868 6692 29484
rect 7420 29538 7476 29550
rect 7420 29486 7422 29538
rect 7474 29486 7476 29538
rect 6748 29316 6804 29326
rect 6748 29222 6804 29260
rect 6636 28802 6692 28812
rect 6636 28532 6692 28542
rect 6524 28530 6692 28532
rect 6524 28478 6638 28530
rect 6690 28478 6692 28530
rect 6524 28476 6692 28478
rect 6636 28466 6692 28476
rect 6860 28418 6916 28430
rect 6860 28366 6862 28418
rect 6914 28366 6916 28418
rect 6300 27186 6468 27188
rect 6300 27134 6302 27186
rect 6354 27134 6468 27186
rect 6300 27132 6468 27134
rect 6636 27860 6692 27870
rect 6300 27122 6356 27132
rect 6188 26910 6190 26962
rect 6242 26910 6244 26962
rect 6188 26898 6244 26910
rect 6412 26852 6468 26862
rect 6300 26850 6468 26852
rect 6300 26798 6414 26850
rect 6466 26798 6468 26850
rect 6300 26796 6468 26798
rect 6300 26516 6356 26796
rect 6412 26786 6468 26796
rect 6636 26740 6692 27804
rect 6748 27748 6804 27758
rect 6748 27524 6804 27692
rect 6748 27458 6804 27468
rect 6300 26460 6580 26516
rect 6524 26402 6580 26460
rect 6524 26350 6526 26402
rect 6578 26350 6580 26402
rect 6300 26290 6356 26302
rect 6300 26238 6302 26290
rect 6354 26238 6356 26290
rect 6300 26180 6356 26238
rect 6300 26114 6356 26124
rect 6076 25778 6132 25788
rect 6188 26068 6244 26078
rect 5740 25566 5742 25618
rect 5794 25566 5796 25618
rect 5180 25506 5236 25518
rect 5180 25454 5182 25506
rect 5234 25454 5236 25506
rect 5180 24948 5236 25454
rect 5180 24882 5236 24892
rect 5292 24836 5348 24846
rect 5292 24742 5348 24780
rect 5516 24724 5572 24734
rect 5516 24630 5572 24668
rect 5404 24610 5460 24622
rect 5404 24558 5406 24610
rect 5458 24558 5460 24610
rect 5404 24500 5460 24558
rect 5404 24444 5684 24500
rect 5244 24332 5508 24342
rect 5300 24276 5348 24332
rect 5404 24276 5452 24332
rect 5244 24266 5508 24276
rect 5404 23492 5460 23502
rect 5404 23378 5460 23436
rect 5404 23326 5406 23378
rect 5458 23326 5460 23378
rect 5404 23314 5460 23326
rect 5068 23202 5124 23212
rect 5292 23266 5348 23278
rect 5292 23214 5294 23266
rect 5346 23214 5348 23266
rect 5292 23156 5348 23214
rect 5516 23268 5572 23278
rect 5628 23268 5684 24444
rect 5516 23266 5684 23268
rect 5516 23214 5518 23266
rect 5570 23214 5684 23266
rect 5516 23212 5684 23214
rect 5740 23380 5796 25566
rect 6188 25620 6244 26012
rect 6524 25844 6580 26350
rect 6524 25778 6580 25788
rect 6524 25620 6580 25630
rect 6188 25618 6580 25620
rect 6188 25566 6526 25618
rect 6578 25566 6580 25618
rect 6188 25564 6580 25566
rect 6524 25554 6580 25564
rect 6524 25450 6580 25462
rect 6300 25394 6356 25406
rect 6524 25398 6526 25450
rect 6578 25398 6580 25450
rect 6524 25396 6580 25398
rect 6300 25342 6302 25394
rect 6354 25342 6356 25394
rect 6076 25284 6132 25294
rect 5964 24948 6020 24958
rect 5964 24722 6020 24892
rect 5964 24670 5966 24722
rect 6018 24670 6020 24722
rect 5964 24658 6020 24670
rect 5964 24052 6020 24062
rect 5964 23958 6020 23996
rect 5852 23826 5908 23838
rect 5852 23774 5854 23826
rect 5906 23774 5908 23826
rect 5852 23492 5908 23774
rect 6076 23492 6132 25228
rect 6300 25284 6356 25342
rect 6300 24948 6356 25228
rect 6412 25340 6580 25396
rect 6636 25394 6692 26684
rect 6748 27186 6804 27198
rect 6748 27134 6750 27186
rect 6802 27134 6804 27186
rect 6748 26516 6804 27134
rect 6748 26450 6804 26460
rect 6748 26292 6804 26302
rect 6748 26198 6804 26236
rect 6636 25342 6638 25394
rect 6690 25342 6692 25394
rect 6412 25172 6468 25340
rect 6636 25330 6692 25342
rect 6748 26068 6804 26078
rect 6748 25284 6804 26012
rect 6860 25508 6916 28366
rect 7196 27860 7252 27870
rect 7196 27858 7364 27860
rect 7196 27806 7198 27858
rect 7250 27806 7364 27858
rect 7196 27804 7364 27806
rect 7196 27794 7252 27804
rect 7308 27634 7364 27804
rect 7308 27582 7310 27634
rect 7362 27582 7364 27634
rect 7308 27570 7364 27582
rect 7084 27076 7140 27086
rect 6972 26964 7028 27002
rect 6972 26290 7028 26908
rect 6972 26238 6974 26290
rect 7026 26238 7028 26290
rect 6972 25844 7028 26238
rect 7084 26178 7140 27020
rect 7196 26964 7252 27002
rect 7196 26898 7252 26908
rect 7308 26852 7364 26862
rect 7308 26758 7364 26796
rect 7308 26628 7364 26638
rect 7420 26628 7476 29486
rect 7644 28754 7700 30044
rect 8316 29988 8372 34200
rect 8764 32116 8820 32126
rect 8316 29922 8372 29932
rect 8540 30322 8596 30334
rect 8540 30270 8542 30322
rect 8594 30270 8596 30322
rect 8204 29538 8260 29550
rect 8204 29486 8206 29538
rect 8258 29486 8260 29538
rect 7756 29428 7812 29438
rect 7756 29334 7812 29372
rect 8092 29314 8148 29326
rect 8092 29262 8094 29314
rect 8146 29262 8148 29314
rect 8092 28980 8148 29262
rect 8092 28914 8148 28924
rect 7644 28702 7646 28754
rect 7698 28702 7700 28754
rect 7644 28690 7700 28702
rect 7868 28642 7924 28654
rect 7868 28590 7870 28642
rect 7922 28590 7924 28642
rect 7532 28532 7588 28542
rect 7532 28530 7700 28532
rect 7532 28478 7534 28530
rect 7586 28478 7700 28530
rect 7532 28476 7700 28478
rect 7532 28466 7588 28476
rect 7532 27634 7588 27646
rect 7532 27582 7534 27634
rect 7586 27582 7588 27634
rect 7532 27074 7588 27582
rect 7532 27022 7534 27074
rect 7586 27022 7588 27074
rect 7532 27010 7588 27022
rect 7364 26572 7476 26628
rect 7084 26126 7086 26178
rect 7138 26126 7140 26178
rect 7084 26114 7140 26126
rect 7196 26404 7252 26414
rect 6972 25788 7140 25844
rect 7084 25508 7140 25788
rect 6860 25452 7028 25508
rect 6860 25284 6916 25294
rect 6748 25282 6916 25284
rect 6748 25230 6862 25282
rect 6914 25230 6916 25282
rect 6748 25228 6916 25230
rect 6860 25218 6916 25228
rect 6412 25106 6468 25116
rect 6300 24882 6356 24892
rect 6636 25060 6692 25070
rect 6412 24724 6468 24734
rect 6300 24722 6468 24724
rect 6300 24670 6414 24722
rect 6466 24670 6468 24722
rect 6300 24668 6468 24670
rect 6300 24052 6356 24668
rect 6412 24658 6468 24668
rect 6636 24724 6692 25004
rect 6860 24948 6916 24958
rect 6972 24948 7028 25452
rect 7084 25442 7140 25452
rect 7196 25394 7252 26348
rect 7308 25508 7364 26572
rect 7420 26404 7476 26414
rect 7420 26310 7476 26348
rect 7420 25508 7476 25518
rect 7308 25506 7476 25508
rect 7308 25454 7422 25506
rect 7474 25454 7476 25506
rect 7308 25452 7476 25454
rect 7196 25342 7198 25394
rect 7250 25342 7252 25394
rect 7196 25330 7252 25342
rect 6860 24946 7028 24948
rect 6860 24894 6862 24946
rect 6914 24894 7028 24946
rect 6860 24892 7028 24894
rect 7084 25282 7140 25294
rect 7084 25230 7086 25282
rect 7138 25230 7140 25282
rect 6860 24882 6916 24892
rect 6524 24612 6580 24622
rect 6412 24500 6468 24510
rect 6412 24162 6468 24444
rect 6412 24110 6414 24162
rect 6466 24110 6468 24162
rect 6412 24098 6468 24110
rect 6300 23986 6356 23996
rect 5852 23426 5908 23436
rect 5964 23436 6132 23492
rect 6188 23938 6244 23950
rect 6188 23886 6190 23938
rect 6242 23886 6244 23938
rect 5516 23202 5572 23212
rect 5292 23090 5348 23100
rect 5244 22764 5508 22774
rect 5300 22708 5348 22764
rect 5404 22708 5452 22764
rect 5244 22698 5508 22708
rect 5068 22484 5124 22494
rect 4956 22482 5124 22484
rect 4956 22430 5070 22482
rect 5122 22430 5124 22482
rect 4956 22428 5124 22430
rect 5740 22484 5796 23324
rect 5852 23268 5908 23278
rect 5852 23174 5908 23212
rect 5852 22484 5908 22494
rect 5740 22482 5908 22484
rect 5740 22430 5854 22482
rect 5906 22430 5908 22482
rect 5740 22428 5908 22430
rect 5068 22148 5124 22428
rect 5852 22418 5908 22428
rect 4956 21586 5012 21598
rect 4956 21534 4958 21586
rect 5010 21534 5012 21586
rect 4956 20804 5012 21534
rect 4956 20738 5012 20748
rect 5068 20914 5124 22092
rect 5292 21812 5348 21822
rect 5292 21718 5348 21756
rect 5852 21700 5908 21710
rect 5292 21588 5348 21598
rect 5292 21494 5348 21532
rect 5628 21588 5684 21598
rect 5628 21586 5796 21588
rect 5628 21534 5630 21586
rect 5682 21534 5796 21586
rect 5628 21532 5796 21534
rect 5628 21522 5684 21532
rect 5244 21196 5508 21206
rect 5300 21140 5348 21196
rect 5404 21140 5452 21196
rect 5244 21130 5508 21140
rect 5740 21026 5796 21532
rect 5740 20974 5742 21026
rect 5794 20974 5796 21026
rect 5740 20962 5796 20974
rect 5068 20862 5070 20914
rect 5122 20862 5124 20914
rect 5068 20356 5124 20862
rect 5852 20804 5908 21644
rect 5068 20188 5124 20300
rect 4956 20132 5124 20188
rect 5404 20802 5908 20804
rect 5404 20750 5854 20802
rect 5906 20750 5908 20802
rect 5404 20748 5908 20750
rect 5404 20242 5460 20748
rect 5852 20738 5908 20748
rect 5740 20580 5796 20618
rect 5740 20514 5796 20524
rect 5404 20190 5406 20242
rect 5458 20190 5460 20242
rect 5404 20132 5460 20190
rect 4956 19796 5012 20132
rect 5404 20066 5460 20076
rect 5740 20356 5796 20366
rect 5180 20018 5236 20030
rect 5180 19966 5182 20018
rect 5234 19966 5236 20018
rect 5180 19796 5236 19966
rect 5740 20018 5796 20300
rect 5740 19966 5742 20018
rect 5794 19966 5796 20018
rect 5740 19954 5796 19966
rect 4956 19740 5124 19796
rect 5068 19346 5124 19740
rect 5180 19730 5236 19740
rect 5244 19628 5508 19638
rect 5300 19572 5348 19628
rect 5404 19572 5452 19628
rect 5244 19562 5508 19572
rect 5740 19460 5796 19470
rect 5740 19366 5796 19404
rect 5068 19294 5070 19346
rect 5122 19294 5124 19346
rect 5068 18788 5124 19294
rect 5852 19236 5908 19246
rect 5628 19234 5908 19236
rect 5628 19182 5854 19234
rect 5906 19182 5908 19234
rect 5628 19180 5908 19182
rect 4956 18732 5124 18788
rect 5292 19012 5348 19022
rect 4844 18452 4900 18462
rect 4844 18358 4900 18396
rect 4956 18340 5012 18732
rect 5180 18676 5236 18686
rect 5068 18564 5124 18574
rect 5068 18470 5124 18508
rect 5180 18562 5236 18620
rect 5180 18510 5182 18562
rect 5234 18510 5236 18562
rect 5180 18498 5236 18510
rect 5292 18564 5348 18956
rect 5292 18498 5348 18508
rect 4956 18284 5124 18340
rect 4732 17042 4788 17052
rect 5068 17778 5124 18284
rect 5628 18228 5684 19180
rect 5852 19170 5908 19180
rect 5740 19012 5796 19022
rect 5964 19012 6020 23436
rect 6188 23380 6244 23886
rect 6076 23324 6244 23380
rect 6076 22036 6132 23324
rect 6188 23156 6244 23166
rect 6524 23156 6580 24556
rect 6636 24388 6692 24668
rect 6748 24722 6804 24734
rect 6748 24670 6750 24722
rect 6802 24670 6804 24722
rect 6748 24500 6804 24670
rect 6972 24724 7028 24734
rect 6972 24630 7028 24668
rect 7084 24500 7140 25230
rect 6748 24444 7140 24500
rect 7308 24836 7364 24846
rect 7308 24722 7364 24780
rect 7308 24670 7310 24722
rect 7362 24670 7364 24722
rect 7308 24388 7364 24670
rect 6636 24332 7028 24388
rect 6636 24052 6692 24062
rect 6636 23938 6692 23996
rect 6636 23886 6638 23938
rect 6690 23886 6692 23938
rect 6636 23874 6692 23886
rect 6972 23826 7028 24332
rect 7308 24322 7364 24332
rect 7420 24276 7476 25452
rect 7644 24946 7700 28476
rect 7868 28420 7924 28590
rect 7868 28354 7924 28364
rect 8092 28084 8148 28094
rect 8092 27990 8148 28028
rect 7756 27972 7812 27982
rect 7756 27878 7812 27916
rect 7756 27524 7812 27534
rect 8204 27524 8260 29486
rect 8540 29538 8596 30270
rect 8540 29486 8542 29538
rect 8594 29486 8596 29538
rect 8540 29428 8596 29486
rect 8540 29362 8596 29372
rect 8652 29540 8708 29550
rect 8652 29426 8708 29484
rect 8652 29374 8654 29426
rect 8706 29374 8708 29426
rect 8652 29362 8708 29374
rect 8428 28866 8484 28878
rect 8428 28814 8430 28866
rect 8482 28814 8484 28866
rect 8428 28754 8484 28814
rect 8428 28702 8430 28754
rect 8482 28702 8484 28754
rect 8428 28690 8484 28702
rect 7756 26514 7812 27468
rect 8092 27468 8260 27524
rect 8540 28084 8596 28094
rect 8540 27746 8596 28028
rect 8764 27972 8820 32060
rect 9436 31892 9492 34200
rect 10556 34132 10612 34200
rect 10892 34132 10948 34300
rect 10556 34076 10948 34132
rect 9436 31826 9492 31836
rect 9276 31388 9540 31398
rect 9332 31332 9380 31388
rect 9436 31332 9484 31388
rect 9276 31322 9540 31332
rect 9436 30994 9492 31006
rect 9436 30942 9438 30994
rect 9490 30942 9492 30994
rect 9436 30212 9492 30942
rect 10108 30882 10164 30894
rect 10108 30830 10110 30882
rect 10162 30830 10164 30882
rect 9772 30212 9828 30222
rect 9436 30210 9828 30212
rect 9436 30158 9774 30210
rect 9826 30158 9828 30210
rect 9436 30156 9828 30158
rect 9324 30100 9380 30110
rect 8988 30098 9380 30100
rect 8988 30046 9326 30098
rect 9378 30046 9380 30098
rect 8988 30044 9380 30046
rect 8876 29988 8932 29998
rect 8876 29894 8932 29932
rect 8988 28644 9044 30044
rect 9324 30034 9380 30044
rect 9436 29988 9492 30026
rect 9436 29922 9492 29932
rect 9276 29820 9540 29830
rect 9332 29764 9380 29820
rect 9436 29764 9484 29820
rect 9276 29754 9540 29764
rect 9100 29652 9156 29662
rect 9100 29092 9156 29596
rect 9660 29540 9716 29550
rect 9548 29484 9660 29540
rect 9100 29026 9156 29036
rect 9324 29316 9380 29326
rect 9212 28868 9268 28878
rect 8764 27906 8820 27916
rect 8876 28588 9044 28644
rect 9100 28812 9212 28868
rect 8540 27694 8542 27746
rect 8594 27694 8596 27746
rect 7980 27188 8036 27198
rect 7980 27094 8036 27132
rect 8092 26962 8148 27468
rect 8428 27412 8484 27422
rect 8092 26910 8094 26962
rect 8146 26910 8148 26962
rect 7756 26462 7758 26514
rect 7810 26462 7812 26514
rect 7756 26450 7812 26462
rect 7868 26850 7924 26862
rect 7868 26798 7870 26850
rect 7922 26798 7924 26850
rect 7868 26516 7924 26798
rect 7868 26068 7924 26460
rect 7868 26002 7924 26012
rect 7980 26852 8036 26862
rect 7980 26180 8036 26796
rect 8092 26404 8148 26910
rect 8204 27076 8260 27086
rect 8204 26962 8260 27020
rect 8204 26910 8206 26962
rect 8258 26910 8260 26962
rect 8204 26898 8260 26910
rect 8092 26338 8148 26348
rect 7756 25506 7812 25518
rect 7756 25454 7758 25506
rect 7810 25454 7812 25506
rect 7756 25172 7812 25454
rect 7980 25396 8036 26124
rect 8428 26290 8484 27356
rect 8540 27300 8596 27694
rect 8540 27074 8596 27244
rect 8540 27022 8542 27074
rect 8594 27022 8596 27074
rect 8540 27010 8596 27022
rect 8652 27636 8708 27646
rect 8540 26740 8596 26750
rect 8652 26740 8708 27580
rect 8876 27076 8932 28588
rect 8988 28420 9044 28430
rect 9100 28420 9156 28812
rect 9212 28802 9268 28812
rect 9324 28866 9380 29260
rect 9324 28814 9326 28866
rect 9378 28814 9380 28866
rect 9324 28754 9380 28814
rect 9548 28868 9604 29484
rect 9660 29474 9716 29484
rect 9660 29316 9716 29326
rect 9772 29316 9828 30156
rect 10108 29650 10164 30830
rect 10108 29598 10110 29650
rect 10162 29598 10164 29650
rect 10108 29586 10164 29598
rect 10556 30098 10612 30110
rect 10556 30046 10558 30098
rect 10610 30046 10612 30098
rect 9716 29260 9828 29316
rect 10220 29538 10276 29550
rect 10220 29486 10222 29538
rect 10274 29486 10276 29538
rect 9660 29222 9716 29260
rect 9996 29202 10052 29214
rect 9996 29150 9998 29202
rect 10050 29150 10052 29202
rect 9772 29092 9828 29102
rect 9660 28868 9716 28878
rect 9548 28866 9716 28868
rect 9548 28814 9662 28866
rect 9714 28814 9716 28866
rect 9548 28812 9716 28814
rect 9660 28802 9716 28812
rect 9324 28702 9326 28754
rect 9378 28702 9380 28754
rect 9324 28690 9380 28702
rect 9772 28644 9828 29036
rect 9996 28756 10052 29150
rect 9996 28700 10164 28756
rect 9772 28588 9940 28644
rect 8988 28418 9156 28420
rect 8988 28366 8990 28418
rect 9042 28366 9156 28418
rect 8988 28364 9156 28366
rect 9772 28420 9828 28430
rect 8988 28354 9044 28364
rect 9772 28326 9828 28364
rect 9276 28252 9540 28262
rect 9332 28196 9380 28252
rect 9436 28196 9484 28252
rect 9276 28186 9540 28196
rect 9660 28196 9716 28206
rect 9212 27972 9268 27982
rect 9100 27746 9156 27758
rect 9100 27694 9102 27746
rect 9154 27694 9156 27746
rect 9100 27188 9156 27694
rect 9100 27122 9156 27132
rect 9212 27186 9268 27916
rect 9212 27134 9214 27186
rect 9266 27134 9268 27186
rect 9212 27122 9268 27134
rect 9548 27972 9604 27982
rect 8876 27010 8932 27020
rect 9548 27074 9604 27916
rect 9660 27970 9716 28140
rect 9660 27918 9662 27970
rect 9714 27918 9716 27970
rect 9660 27412 9716 27918
rect 9884 27970 9940 28588
rect 9996 28532 10052 28542
rect 9996 28438 10052 28476
rect 10108 28308 10164 28700
rect 10220 28420 10276 29486
rect 10556 29540 10612 30046
rect 10556 29474 10612 29484
rect 10332 29428 10388 29438
rect 10332 28642 10388 29372
rect 10892 29316 10948 29326
rect 10892 29222 10948 29260
rect 11004 29204 11060 29214
rect 11004 29202 11172 29204
rect 11004 29150 11006 29202
rect 11058 29150 11172 29202
rect 11004 29148 11172 29150
rect 11004 29138 11060 29148
rect 10332 28590 10334 28642
rect 10386 28590 10388 28642
rect 10332 28578 10388 28590
rect 11004 28756 11060 28766
rect 10220 28354 10276 28364
rect 10892 28532 10948 28542
rect 9884 27918 9886 27970
rect 9938 27918 9940 27970
rect 9884 27906 9940 27918
rect 9996 28252 10164 28308
rect 10780 28308 10836 28318
rect 9772 27858 9828 27870
rect 9772 27806 9774 27858
rect 9826 27806 9828 27858
rect 9772 27636 9828 27806
rect 9772 27570 9828 27580
rect 9660 27346 9716 27356
rect 9996 27186 10052 28252
rect 10780 27972 10836 28252
rect 10780 27878 10836 27916
rect 10668 27860 10724 27870
rect 10444 27858 10724 27860
rect 10444 27806 10670 27858
rect 10722 27806 10724 27858
rect 10444 27804 10724 27806
rect 10332 27636 10388 27646
rect 10444 27636 10500 27804
rect 10668 27794 10724 27804
rect 10780 27636 10836 27646
rect 10332 27634 10500 27636
rect 10332 27582 10334 27634
rect 10386 27582 10500 27634
rect 10332 27580 10500 27582
rect 10332 27570 10388 27580
rect 10444 27300 10500 27580
rect 9996 27134 9998 27186
rect 10050 27134 10052 27186
rect 9996 27122 10052 27134
rect 10108 27244 10500 27300
rect 10556 27634 10836 27636
rect 10556 27582 10782 27634
rect 10834 27582 10836 27634
rect 10556 27580 10836 27582
rect 9548 27022 9550 27074
rect 9602 27022 9604 27074
rect 9548 27010 9604 27022
rect 9772 26964 9828 26974
rect 9772 26852 9828 26908
rect 8596 26684 8708 26740
rect 9660 26850 9828 26852
rect 9660 26798 9774 26850
rect 9826 26798 9828 26850
rect 9660 26796 9828 26798
rect 9276 26684 9540 26694
rect 8540 26402 8596 26684
rect 9332 26628 9380 26684
rect 9436 26628 9484 26684
rect 9276 26618 9540 26628
rect 8540 26350 8542 26402
rect 8594 26350 8596 26402
rect 8540 26338 8596 26350
rect 8428 26238 8430 26290
rect 8482 26238 8484 26290
rect 8428 25732 8484 26238
rect 8988 26292 9044 26302
rect 9212 26292 9268 26302
rect 8988 26290 9212 26292
rect 8988 26238 8990 26290
rect 9042 26238 9212 26290
rect 8988 26236 9212 26238
rect 8988 26226 9044 26236
rect 9212 26226 9268 26236
rect 8764 26178 8820 26190
rect 8764 26126 8766 26178
rect 8818 26126 8820 26178
rect 8764 25956 8820 26126
rect 8764 25900 9044 25956
rect 8428 25666 8484 25676
rect 8876 25732 8932 25742
rect 7980 25340 8372 25396
rect 7756 25106 7812 25116
rect 7644 24894 7646 24946
rect 7698 24894 7700 24946
rect 7644 24882 7700 24894
rect 7756 24948 7812 24958
rect 7756 24946 7924 24948
rect 7756 24894 7758 24946
rect 7810 24894 7924 24946
rect 7756 24892 7924 24894
rect 7756 24882 7812 24892
rect 7420 24210 7476 24220
rect 7532 24722 7588 24734
rect 7532 24670 7534 24722
rect 7586 24670 7588 24722
rect 7532 24164 7588 24670
rect 7868 24276 7924 24892
rect 8316 24946 8372 25340
rect 8316 24894 8318 24946
rect 8370 24894 8372 24946
rect 8316 24882 8372 24894
rect 8540 25172 8596 25182
rect 8540 24946 8596 25116
rect 8540 24894 8542 24946
rect 8594 24894 8596 24946
rect 7532 24108 7812 24164
rect 7756 24050 7812 24108
rect 7756 23998 7758 24050
rect 7810 23998 7812 24050
rect 7756 23986 7812 23998
rect 7196 23940 7252 23950
rect 7196 23846 7252 23884
rect 7868 23938 7924 24220
rect 7868 23886 7870 23938
rect 7922 23886 7924 23938
rect 7868 23874 7924 23886
rect 7980 24722 8036 24734
rect 7980 24670 7982 24722
rect 8034 24670 8036 24722
rect 7980 24500 8036 24670
rect 8428 24610 8484 24622
rect 8428 24558 8430 24610
rect 8482 24558 8484 24610
rect 8428 24500 8484 24558
rect 7980 24444 8484 24500
rect 6972 23774 6974 23826
rect 7026 23774 7028 23826
rect 6972 23762 7028 23774
rect 7644 23716 7700 23726
rect 7644 23622 7700 23660
rect 6188 23154 6580 23156
rect 6188 23102 6190 23154
rect 6242 23102 6580 23154
rect 6188 23100 6580 23102
rect 6636 23492 6692 23502
rect 6636 23154 6692 23436
rect 6972 23380 7028 23390
rect 6972 23286 7028 23324
rect 6636 23102 6638 23154
rect 6690 23102 6692 23154
rect 6188 23090 6244 23100
rect 6636 23044 6692 23102
rect 6636 22978 6692 22988
rect 6748 23266 6804 23278
rect 6748 23214 6750 23266
rect 6802 23214 6804 23266
rect 6076 21980 6356 22036
rect 6188 21812 6244 21822
rect 6188 21718 6244 21756
rect 6076 21700 6132 21710
rect 6076 21606 6132 21644
rect 6188 21362 6244 21374
rect 6188 21310 6190 21362
rect 6242 21310 6244 21362
rect 6188 20802 6244 21310
rect 6188 20750 6190 20802
rect 6242 20750 6244 20802
rect 6188 20738 6244 20750
rect 5740 18918 5796 18956
rect 5852 18956 6020 19012
rect 6076 20020 6132 20030
rect 5852 18788 5908 18956
rect 5244 18060 5508 18070
rect 5300 18004 5348 18060
rect 5404 18004 5452 18060
rect 5244 17994 5508 18004
rect 5068 17726 5070 17778
rect 5122 17726 5124 17778
rect 4396 16942 4398 16994
rect 4450 16942 4452 16994
rect 4396 16930 4452 16942
rect 4956 16994 5012 17006
rect 4956 16942 4958 16994
rect 5010 16942 5012 16994
rect 4844 16884 4900 16894
rect 4956 16884 5012 16942
rect 4844 16882 5012 16884
rect 4844 16830 4846 16882
rect 4898 16830 5012 16882
rect 4844 16828 5012 16830
rect 4844 16818 4900 16828
rect 4172 16594 4228 16604
rect 4844 16660 4900 16670
rect 4900 16604 5012 16660
rect 4844 16594 4900 16604
rect 3836 16046 3838 16098
rect 3890 16046 3892 16098
rect 3836 16034 3892 16046
rect 4956 16100 5012 16604
rect 4956 16006 5012 16044
rect 4172 15988 4228 15998
rect 4396 15988 4452 15998
rect 4172 15986 4452 15988
rect 4172 15934 4174 15986
rect 4226 15934 4398 15986
rect 4450 15934 4452 15986
rect 4172 15932 4452 15934
rect 4172 15922 4228 15932
rect 4396 15922 4452 15932
rect 4732 15988 4788 15998
rect 4732 15986 4900 15988
rect 4732 15934 4734 15986
rect 4786 15934 4900 15986
rect 4732 15932 4900 15934
rect 4732 15922 4788 15932
rect 2492 15876 2548 15886
rect 2492 15426 2548 15820
rect 2492 15374 2494 15426
rect 2546 15374 2548 15426
rect 2492 15362 2548 15374
rect 3948 15874 4004 15886
rect 3948 15822 3950 15874
rect 4002 15822 4004 15874
rect 3948 15764 4004 15822
rect 4508 15876 4564 15886
rect 4508 15782 4564 15820
rect 1820 15262 1822 15314
rect 1874 15262 1876 15314
rect 1820 14530 1876 15262
rect 2492 15204 2548 15214
rect 2492 14642 2548 15148
rect 3948 15148 4004 15708
rect 4844 15652 4900 15932
rect 5068 15764 5124 17726
rect 5628 17556 5684 18172
rect 5292 17554 5684 17556
rect 5292 17502 5630 17554
rect 5682 17502 5684 17554
rect 5292 17500 5684 17502
rect 5180 17220 5236 17230
rect 5180 17106 5236 17164
rect 5180 17054 5182 17106
rect 5234 17054 5236 17106
rect 5180 17042 5236 17054
rect 5292 16994 5348 17500
rect 5628 17490 5684 17500
rect 5740 18732 5908 18788
rect 5404 17220 5460 17230
rect 5460 17164 5572 17220
rect 5404 17154 5460 17164
rect 5292 16942 5294 16994
rect 5346 16942 5348 16994
rect 5292 16930 5348 16942
rect 5516 16660 5572 17164
rect 5628 17108 5684 17118
rect 5740 17108 5796 18732
rect 5964 18676 6020 18686
rect 6076 18676 6132 19964
rect 6300 19124 6356 21980
rect 6748 21812 6804 23214
rect 7756 23268 7812 23278
rect 7980 23268 8036 24444
rect 8540 24276 8596 24894
rect 8540 24210 8596 24220
rect 8652 24948 8708 24958
rect 7756 23266 8036 23268
rect 7756 23214 7758 23266
rect 7810 23214 8036 23266
rect 7756 23212 8036 23214
rect 8204 23938 8260 23950
rect 8652 23940 8708 24892
rect 8204 23886 8206 23938
rect 8258 23886 8260 23938
rect 7756 23202 7812 23212
rect 7196 23154 7252 23166
rect 7196 23102 7198 23154
rect 7250 23102 7252 23154
rect 7196 23044 7252 23102
rect 7308 23156 7364 23166
rect 7308 23062 7364 23100
rect 7420 23154 7476 23166
rect 7420 23102 7422 23154
rect 7474 23102 7476 23154
rect 7196 22978 7252 22988
rect 6748 21718 6804 21756
rect 6636 21588 6692 21598
rect 6412 21586 6692 21588
rect 6412 21534 6638 21586
rect 6690 21534 6692 21586
rect 6412 21532 6692 21534
rect 6412 20020 6468 21532
rect 6636 21522 6692 21532
rect 6972 21588 7028 21598
rect 6972 21494 7028 21532
rect 7308 21586 7364 21598
rect 7308 21534 7310 21586
rect 7362 21534 7364 21586
rect 6636 21028 6692 21038
rect 6636 20802 6692 20972
rect 7308 21028 7364 21534
rect 7308 20962 7364 20972
rect 6636 20750 6638 20802
rect 6690 20750 6692 20802
rect 6636 20738 6692 20750
rect 6860 20804 6916 20814
rect 6860 20710 6916 20748
rect 7196 20802 7252 20814
rect 7196 20750 7198 20802
rect 7250 20750 7252 20802
rect 6524 20578 6580 20590
rect 6524 20526 6526 20578
rect 6578 20526 6580 20578
rect 6524 20130 6580 20526
rect 7196 20356 7252 20750
rect 7196 20290 7252 20300
rect 7308 20804 7364 20814
rect 6524 20078 6526 20130
rect 6578 20078 6580 20130
rect 6524 20066 6580 20078
rect 6412 19954 6468 19964
rect 6300 19058 6356 19068
rect 6020 18620 6132 18676
rect 5964 18582 6020 18620
rect 7308 18564 7364 20748
rect 7420 19012 7476 23102
rect 7532 21698 7588 21710
rect 7532 21646 7534 21698
rect 7586 21646 7588 21698
rect 7532 21476 7588 21646
rect 7644 21700 7700 21710
rect 7644 21698 7812 21700
rect 7644 21646 7646 21698
rect 7698 21646 7812 21698
rect 7644 21644 7812 21646
rect 7644 21634 7700 21644
rect 7532 21420 7700 21476
rect 7644 19908 7700 21420
rect 7644 19842 7700 19852
rect 7532 19796 7588 19806
rect 7532 19124 7588 19740
rect 7532 19068 7700 19124
rect 7420 18956 7588 19012
rect 7420 18564 7476 18574
rect 7308 18562 7476 18564
rect 7308 18510 7422 18562
rect 7474 18510 7476 18562
rect 7308 18508 7476 18510
rect 7420 18498 7476 18508
rect 6300 18452 6356 18462
rect 6300 18358 6356 18396
rect 6748 18452 6804 18462
rect 6804 18396 7028 18452
rect 6748 18358 6804 18396
rect 6748 17780 6804 17790
rect 5852 17668 5908 17678
rect 5852 17574 5908 17612
rect 6748 17554 6804 17724
rect 6748 17502 6750 17554
rect 6802 17502 6804 17554
rect 6748 17490 6804 17502
rect 5628 17106 5796 17108
rect 5628 17054 5630 17106
rect 5682 17054 5796 17106
rect 5628 17052 5796 17054
rect 6636 17108 6692 17118
rect 5628 17042 5684 17052
rect 6636 17014 6692 17052
rect 5852 16994 5908 17006
rect 5852 16942 5854 16994
rect 5906 16942 5908 16994
rect 5516 16604 5796 16660
rect 5244 16492 5508 16502
rect 5300 16436 5348 16492
rect 5404 16436 5452 16492
rect 5244 16426 5508 16436
rect 5628 16100 5684 16110
rect 5628 16006 5684 16044
rect 5068 15708 5684 15764
rect 4844 15596 5124 15652
rect 4620 15540 4676 15550
rect 4620 15202 4676 15484
rect 5068 15538 5124 15596
rect 5068 15486 5070 15538
rect 5122 15486 5124 15538
rect 5068 15474 5124 15486
rect 5292 15540 5348 15550
rect 5292 15446 5348 15484
rect 5404 15316 5460 15326
rect 5404 15222 5460 15260
rect 5628 15316 5684 15708
rect 5740 15540 5796 16604
rect 5852 15764 5908 16942
rect 5964 16996 6020 17006
rect 6300 16996 6356 17006
rect 5964 16994 6300 16996
rect 5964 16942 5966 16994
rect 6018 16942 6300 16994
rect 5964 16940 6300 16942
rect 5964 16930 6020 16940
rect 6300 16902 6356 16940
rect 6412 16996 6468 17006
rect 6412 16994 6580 16996
rect 6412 16942 6414 16994
rect 6466 16942 6580 16994
rect 6412 16940 6580 16942
rect 6412 16930 6468 16940
rect 5964 16156 6356 16212
rect 5964 16098 6020 16156
rect 5964 16046 5966 16098
rect 6018 16046 6020 16098
rect 5964 16034 6020 16046
rect 6300 16100 6356 16156
rect 6412 16100 6468 16110
rect 6300 16098 6468 16100
rect 6300 16046 6414 16098
rect 6466 16046 6468 16098
rect 6300 16044 6468 16046
rect 6412 16034 6468 16044
rect 6188 15986 6244 15998
rect 6188 15934 6190 15986
rect 6242 15934 6244 15986
rect 5852 15698 5908 15708
rect 5964 15874 6020 15886
rect 5964 15822 5966 15874
rect 6018 15822 6020 15874
rect 5740 15474 5796 15484
rect 5852 15316 5908 15326
rect 5628 15314 5908 15316
rect 5628 15262 5854 15314
rect 5906 15262 5908 15314
rect 5628 15260 5908 15262
rect 4620 15150 4622 15202
rect 4674 15150 4676 15202
rect 3948 15092 4564 15148
rect 4620 15138 4676 15150
rect 2492 14590 2494 14642
rect 2546 14590 2548 14642
rect 2492 14578 2548 14590
rect 4508 14644 4564 15092
rect 5244 14924 5508 14934
rect 5300 14868 5348 14924
rect 5404 14868 5452 14924
rect 5244 14858 5508 14868
rect 5628 14756 5684 15260
rect 5852 15250 5908 15260
rect 5964 15204 6020 15822
rect 6188 15540 6244 15934
rect 6524 15876 6580 16940
rect 6860 16994 6916 17006
rect 6860 16942 6862 16994
rect 6914 16942 6916 16994
rect 6748 15988 6804 15998
rect 6860 15988 6916 16942
rect 6972 16884 7028 18396
rect 7196 17892 7252 17902
rect 7252 17836 7364 17892
rect 7196 17826 7252 17836
rect 7084 17666 7140 17678
rect 7084 17614 7086 17666
rect 7138 17614 7140 17666
rect 7084 17444 7140 17614
rect 7308 17666 7364 17836
rect 7532 17668 7588 18956
rect 7644 18676 7700 19068
rect 7756 18788 7812 21644
rect 7868 21586 7924 21598
rect 7868 21534 7870 21586
rect 7922 21534 7924 21586
rect 7868 19234 7924 21534
rect 8092 21474 8148 21486
rect 8092 21422 8094 21474
rect 8146 21422 8148 21474
rect 7980 20916 8036 20926
rect 8092 20916 8148 21422
rect 7980 20914 8148 20916
rect 7980 20862 7982 20914
rect 8034 20862 8148 20914
rect 7980 20860 8148 20862
rect 7980 20850 8036 20860
rect 7980 20132 8036 20142
rect 8036 20076 8148 20132
rect 7980 20066 8036 20076
rect 7868 19182 7870 19234
rect 7922 19182 7924 19234
rect 7868 19170 7924 19182
rect 7980 19908 8036 19918
rect 7980 19012 8036 19852
rect 8092 19236 8148 20076
rect 8204 19348 8260 23886
rect 8540 23884 8708 23940
rect 8764 24836 8820 24846
rect 8764 23938 8820 24780
rect 8876 24722 8932 25676
rect 8988 24948 9044 25900
rect 9548 25732 9604 25742
rect 9660 25732 9716 26796
rect 9772 26758 9828 26796
rect 9996 26852 10052 26862
rect 9996 26758 10052 26796
rect 9772 26404 9828 26414
rect 9772 26310 9828 26348
rect 9996 26292 10052 26302
rect 9548 25730 9716 25732
rect 9548 25678 9550 25730
rect 9602 25678 9716 25730
rect 9548 25676 9716 25678
rect 9884 26068 9940 26078
rect 9884 25730 9940 26012
rect 9884 25678 9886 25730
rect 9938 25678 9940 25730
rect 9548 25666 9604 25676
rect 9884 25666 9940 25678
rect 9996 25732 10052 26236
rect 9996 25666 10052 25676
rect 9212 25620 9268 25630
rect 9212 25526 9268 25564
rect 10108 25508 10164 27244
rect 10220 27076 10276 27086
rect 10220 27074 10500 27076
rect 10220 27022 10222 27074
rect 10274 27022 10500 27074
rect 10220 27020 10500 27022
rect 10220 27010 10276 27020
rect 10332 26740 10388 26750
rect 10220 25508 10276 25518
rect 9772 25506 10276 25508
rect 9772 25454 10222 25506
rect 10274 25454 10276 25506
rect 9772 25452 10276 25454
rect 9660 25396 9716 25406
rect 9548 25284 9604 25322
rect 9660 25302 9716 25340
rect 9548 25218 9604 25228
rect 9276 25116 9540 25126
rect 9332 25060 9380 25116
rect 9436 25060 9484 25116
rect 9276 25050 9540 25060
rect 8988 24892 9604 24948
rect 8876 24670 8878 24722
rect 8930 24670 8932 24722
rect 8876 24658 8932 24670
rect 9548 24722 9604 24892
rect 9548 24670 9550 24722
rect 9602 24670 9604 24722
rect 9548 24658 9604 24670
rect 9772 24722 9828 25452
rect 10220 25442 10276 25452
rect 9996 25284 10052 25294
rect 9996 24836 10052 25228
rect 9996 24770 10052 24780
rect 9772 24670 9774 24722
rect 9826 24670 9828 24722
rect 9772 24658 9828 24670
rect 9996 24498 10052 24510
rect 9996 24446 9998 24498
rect 10050 24446 10052 24498
rect 8764 23886 8766 23938
rect 8818 23886 8820 23938
rect 8428 23716 8484 23726
rect 8428 23622 8484 23660
rect 8540 23380 8596 23884
rect 8764 23874 8820 23886
rect 8876 24276 8932 24286
rect 8652 23716 8708 23726
rect 8876 23716 8932 24220
rect 9996 23940 10052 24446
rect 10108 24500 10164 24510
rect 10108 24406 10164 24444
rect 10108 23940 10164 23950
rect 8652 23714 8932 23716
rect 8652 23662 8654 23714
rect 8706 23662 8932 23714
rect 8652 23660 8932 23662
rect 9660 23938 10164 23940
rect 9660 23886 10110 23938
rect 10162 23886 10164 23938
rect 9660 23884 10164 23886
rect 8652 23650 8708 23660
rect 9276 23548 9540 23558
rect 9332 23492 9380 23548
rect 9436 23492 9484 23548
rect 9276 23482 9540 23492
rect 8652 23380 8708 23390
rect 8540 23378 8708 23380
rect 8540 23326 8654 23378
rect 8706 23326 8708 23378
rect 8540 23324 8708 23326
rect 8652 23314 8708 23324
rect 8876 23266 8932 23278
rect 8876 23214 8878 23266
rect 8930 23214 8932 23266
rect 8316 21586 8372 21598
rect 8316 21534 8318 21586
rect 8370 21534 8372 21586
rect 8316 20188 8372 21534
rect 8428 21586 8484 21598
rect 8428 21534 8430 21586
rect 8482 21534 8484 21586
rect 8428 20804 8484 21534
rect 8428 20738 8484 20748
rect 8316 20132 8820 20188
rect 8652 19908 8708 19918
rect 8652 19814 8708 19852
rect 8204 19292 8372 19348
rect 8092 19180 8260 19236
rect 8204 19122 8260 19180
rect 8204 19070 8206 19122
rect 8258 19070 8260 19122
rect 8204 19058 8260 19070
rect 8092 19012 8148 19022
rect 7980 19010 8148 19012
rect 7980 18958 8094 19010
rect 8146 18958 8148 19010
rect 7980 18956 8148 18958
rect 8092 18946 8148 18956
rect 8204 18788 8260 18798
rect 7756 18732 8204 18788
rect 7644 18620 7924 18676
rect 7308 17614 7310 17666
rect 7362 17614 7364 17666
rect 7308 17602 7364 17614
rect 7420 17612 7588 17668
rect 7756 18450 7812 18462
rect 7756 18398 7758 18450
rect 7810 18398 7812 18450
rect 7420 17444 7476 17612
rect 7644 17554 7700 17566
rect 7644 17502 7646 17554
rect 7698 17502 7700 17554
rect 7084 17378 7140 17388
rect 7308 17388 7476 17444
rect 7532 17442 7588 17454
rect 7532 17390 7534 17442
rect 7586 17390 7588 17442
rect 7084 16884 7140 16894
rect 6972 16828 7084 16884
rect 7084 16790 7140 16828
rect 6748 15986 6916 15988
rect 6748 15934 6750 15986
rect 6802 15934 6916 15986
rect 6748 15932 6916 15934
rect 6748 15922 6804 15932
rect 6188 15474 6244 15484
rect 6412 15820 6580 15876
rect 6636 15876 6692 15886
rect 6412 15428 6468 15820
rect 6636 15782 6692 15820
rect 6748 15540 6804 15550
rect 6748 15446 6804 15484
rect 6300 15316 6356 15354
rect 6300 15250 6356 15260
rect 6412 15148 6468 15372
rect 5964 15138 6020 15148
rect 5180 14700 5684 14756
rect 6076 15092 6468 15148
rect 6524 15316 6580 15326
rect 4620 14644 4676 14654
rect 4508 14642 4676 14644
rect 4508 14590 4622 14642
rect 4674 14590 4676 14642
rect 4508 14588 4676 14590
rect 4620 14578 4676 14588
rect 5180 14642 5236 14700
rect 5180 14590 5182 14642
rect 5234 14590 5236 14642
rect 5180 14578 5236 14590
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 14466 1876 14478
rect 6076 14196 6132 15092
rect 6524 14530 6580 15260
rect 6524 14478 6526 14530
rect 6578 14478 6580 14530
rect 6524 14466 6580 14478
rect 6636 15314 6692 15326
rect 6636 15262 6638 15314
rect 6690 15262 6692 15314
rect 6636 14532 6692 15262
rect 6748 15204 6804 15214
rect 6860 15204 6916 15932
rect 6972 15428 7028 15438
rect 7196 15428 7252 15438
rect 6972 15334 7028 15372
rect 7084 15372 7196 15428
rect 7084 15314 7140 15372
rect 7196 15362 7252 15372
rect 7084 15262 7086 15314
rect 7138 15262 7140 15314
rect 7084 15250 7140 15262
rect 6804 15148 6916 15204
rect 6748 15138 6804 15148
rect 6860 14532 6916 14542
rect 6636 14530 6916 14532
rect 6636 14478 6862 14530
rect 6914 14478 6916 14530
rect 6636 14476 6916 14478
rect 6860 14466 6916 14476
rect 7196 14532 7252 14542
rect 7196 14438 7252 14476
rect 5628 14140 6132 14196
rect 6748 14306 6804 14318
rect 6748 14254 6750 14306
rect 6802 14254 6804 14306
rect 5244 13356 5508 13366
rect 5300 13300 5348 13356
rect 5404 13300 5452 13356
rect 5244 13290 5508 13300
rect 5628 13074 5684 14140
rect 5628 13022 5630 13074
rect 5682 13022 5684 13074
rect 5628 13010 5684 13022
rect 6188 13746 6244 13758
rect 6188 13694 6190 13746
rect 6242 13694 6244 13746
rect 6188 12964 6244 13694
rect 5244 11788 5508 11798
rect 5300 11732 5348 11788
rect 5404 11732 5452 11788
rect 5244 11722 5508 11732
rect 6188 11394 6244 12908
rect 6748 12852 6804 14254
rect 7308 14308 7364 17388
rect 7532 17220 7588 17390
rect 7532 17154 7588 17164
rect 7644 16996 7700 17502
rect 7756 17444 7812 18398
rect 7756 17378 7812 17388
rect 7868 17220 7924 18620
rect 8204 18674 8260 18732
rect 8204 18622 8206 18674
rect 8258 18622 8260 18674
rect 8204 18610 8260 18622
rect 8204 17444 8260 17454
rect 8204 17350 8260 17388
rect 7644 16930 7700 16940
rect 7756 17164 7924 17220
rect 7532 16884 7588 16894
rect 7532 16210 7588 16828
rect 7532 16158 7534 16210
rect 7586 16158 7588 16210
rect 7532 16146 7588 16158
rect 7756 15988 7812 17164
rect 8204 17108 8260 17118
rect 8316 17108 8372 19292
rect 8764 19234 8820 20132
rect 8764 19182 8766 19234
rect 8818 19182 8820 19234
rect 8764 19170 8820 19182
rect 8876 19012 8932 23214
rect 8988 23268 9044 23278
rect 9548 23268 9604 23278
rect 9660 23268 9716 23884
rect 10108 23828 10164 23884
rect 10108 23762 10164 23772
rect 8988 23266 9716 23268
rect 8988 23214 8990 23266
rect 9042 23214 9550 23266
rect 9602 23214 9716 23266
rect 8988 23212 9716 23214
rect 9884 23714 9940 23726
rect 9884 23662 9886 23714
rect 9938 23662 9940 23714
rect 8988 23202 9044 23212
rect 9548 23202 9604 23212
rect 9772 23156 9828 23166
rect 9884 23156 9940 23662
rect 9772 23154 9940 23156
rect 9772 23102 9774 23154
rect 9826 23102 9940 23154
rect 9772 23100 9940 23102
rect 10220 23714 10276 23726
rect 10220 23662 10222 23714
rect 10274 23662 10276 23714
rect 9276 21980 9540 21990
rect 9332 21924 9380 21980
rect 9436 21924 9484 21980
rect 9276 21914 9540 21924
rect 9548 21700 9604 21710
rect 9548 21606 9604 21644
rect 9660 21698 9716 21710
rect 9660 21646 9662 21698
rect 9714 21646 9716 21698
rect 8988 20916 9044 20926
rect 8988 19122 9044 20860
rect 9660 20916 9716 21646
rect 9660 20850 9716 20860
rect 9772 20468 9828 23100
rect 9884 21588 9940 21598
rect 9884 21586 10052 21588
rect 9884 21534 9886 21586
rect 9938 21534 10052 21586
rect 9884 21532 10052 21534
rect 9884 21522 9940 21532
rect 9884 20468 9940 20478
rect 9276 20412 9540 20422
rect 9772 20412 9884 20468
rect 9332 20356 9380 20412
rect 9436 20356 9484 20412
rect 9276 20346 9540 20356
rect 9548 20244 9604 20254
rect 9548 19346 9604 20188
rect 9548 19294 9550 19346
rect 9602 19294 9604 19346
rect 9548 19282 9604 19294
rect 9772 20020 9828 20030
rect 9660 19236 9716 19246
rect 8988 19070 8990 19122
rect 9042 19070 9044 19122
rect 8988 19058 9044 19070
rect 9100 19124 9156 19134
rect 8876 18946 8932 18956
rect 9100 18788 9156 19068
rect 9276 18844 9540 18854
rect 9332 18788 9380 18844
rect 9436 18788 9484 18844
rect 9276 18778 9540 18788
rect 9100 18722 9156 18732
rect 9212 18676 9268 18686
rect 8540 18564 8596 18574
rect 8540 18450 8596 18508
rect 8540 18398 8542 18450
rect 8594 18398 8596 18450
rect 8540 18386 8596 18398
rect 8988 18564 9044 18574
rect 8988 18450 9044 18508
rect 8988 18398 8990 18450
rect 9042 18398 9044 18450
rect 8988 18386 9044 18398
rect 9212 17666 9268 18620
rect 9660 18564 9716 19180
rect 9772 18788 9828 19964
rect 9772 18722 9828 18732
rect 9884 18564 9940 20412
rect 9996 19908 10052 21532
rect 10108 20916 10164 20926
rect 10220 20916 10276 23662
rect 10332 22596 10388 26684
rect 10444 25284 10500 27020
rect 10556 26290 10612 27580
rect 10780 27570 10836 27580
rect 10892 27412 10948 28476
rect 10668 27356 10948 27412
rect 10668 27186 10724 27356
rect 11004 27188 11060 28700
rect 10668 27134 10670 27186
rect 10722 27134 10724 27186
rect 10668 27122 10724 27134
rect 10780 27132 11060 27188
rect 10780 27074 10836 27132
rect 10780 27022 10782 27074
rect 10834 27022 10836 27074
rect 10668 26964 10724 27002
rect 10668 26898 10724 26908
rect 10780 26404 10836 27022
rect 11004 26962 11060 26974
rect 11004 26910 11006 26962
rect 11058 26910 11060 26962
rect 11004 26628 11060 26910
rect 11116 26852 11172 29148
rect 11228 28868 11284 34300
rect 11648 34200 11760 35000
rect 12768 34200 12880 35000
rect 13888 34200 14000 35000
rect 15008 34200 15120 35000
rect 16128 34200 16240 35000
rect 17248 34200 17360 35000
rect 18368 34200 18480 35000
rect 19488 34200 19600 35000
rect 20608 34200 20720 35000
rect 21728 34200 21840 35000
rect 22848 34200 22960 35000
rect 23968 34200 24080 35000
rect 25088 34200 25200 35000
rect 26208 34200 26320 35000
rect 27328 34200 27440 35000
rect 28448 34200 28560 35000
rect 29568 34200 29680 35000
rect 30688 34200 30800 35000
rect 30940 34300 31556 34356
rect 11676 32564 11732 34200
rect 11564 32508 11732 32564
rect 11340 29540 11396 29550
rect 11340 29538 11508 29540
rect 11340 29486 11342 29538
rect 11394 29486 11508 29538
rect 11340 29484 11508 29486
rect 11340 29474 11396 29484
rect 11340 28868 11396 28878
rect 11228 28866 11396 28868
rect 11228 28814 11342 28866
rect 11394 28814 11396 28866
rect 11228 28812 11396 28814
rect 11340 28802 11396 28812
rect 11228 27858 11284 27870
rect 11228 27806 11230 27858
rect 11282 27806 11284 27858
rect 11228 27524 11284 27806
rect 11452 27636 11508 29484
rect 11564 29204 11620 32508
rect 12236 30996 12292 31006
rect 12236 30882 12292 30940
rect 12236 30830 12238 30882
rect 12290 30830 12292 30882
rect 11676 29652 11732 29662
rect 11676 29558 11732 29596
rect 12124 29428 12180 29438
rect 11564 29148 11732 29204
rect 11452 27570 11508 27580
rect 11564 28644 11620 28654
rect 11228 27458 11284 27468
rect 11228 26964 11284 26974
rect 11228 26870 11284 26908
rect 11116 26786 11172 26796
rect 11004 26572 11284 26628
rect 11116 26404 11172 26414
rect 10780 26402 11172 26404
rect 10780 26350 11118 26402
rect 11170 26350 11172 26402
rect 10780 26348 11172 26350
rect 11116 26338 11172 26348
rect 10556 26238 10558 26290
rect 10610 26238 10612 26290
rect 10556 25508 10612 26238
rect 10668 26180 10724 26190
rect 10668 26068 10724 26124
rect 10780 26068 10836 26078
rect 10668 26066 10836 26068
rect 10668 26014 10782 26066
rect 10834 26014 10836 26066
rect 10668 26012 10836 26014
rect 10780 26002 10836 26012
rect 10892 26068 10948 26078
rect 10948 26012 11060 26068
rect 10892 26002 10948 26012
rect 10556 25414 10612 25452
rect 11004 25506 11060 26012
rect 11228 26066 11284 26572
rect 11228 26014 11230 26066
rect 11282 26014 11284 26066
rect 11228 26002 11284 26014
rect 11340 26066 11396 26078
rect 11340 26014 11342 26066
rect 11394 26014 11396 26066
rect 11340 25732 11396 26014
rect 11004 25454 11006 25506
rect 11058 25454 11060 25506
rect 11004 25442 11060 25454
rect 11116 25676 11396 25732
rect 10668 25284 10724 25294
rect 10444 25282 10724 25284
rect 10444 25230 10670 25282
rect 10722 25230 10724 25282
rect 10444 25228 10724 25230
rect 10668 25218 10724 25228
rect 10892 25282 10948 25294
rect 10892 25230 10894 25282
rect 10946 25230 10948 25282
rect 10556 25060 10612 25070
rect 10556 24946 10612 25004
rect 10556 24894 10558 24946
rect 10610 24894 10612 24946
rect 10556 24882 10612 24894
rect 10892 24948 10948 25230
rect 10892 24882 10948 24892
rect 11004 24836 11060 24846
rect 11116 24836 11172 25676
rect 11340 25508 11396 25546
rect 11340 25442 11396 25452
rect 11452 25338 11508 25350
rect 11452 25286 11454 25338
rect 11506 25286 11508 25338
rect 11452 25172 11508 25286
rect 11340 25116 11508 25172
rect 11340 25060 11396 25116
rect 11340 24994 11396 25004
rect 11564 24948 11620 28588
rect 11676 28084 11732 29148
rect 12124 28644 12180 29372
rect 12124 28578 12180 28588
rect 12236 28308 12292 30830
rect 12796 30212 12852 34200
rect 13916 31220 13972 34200
rect 13692 31164 13972 31220
rect 13356 30884 13412 30894
rect 13356 30790 13412 30828
rect 13468 30772 13524 30810
rect 13468 30706 13524 30716
rect 13308 30604 13572 30614
rect 13364 30548 13412 30604
rect 13468 30548 13516 30604
rect 13308 30538 13572 30548
rect 12796 30156 13188 30212
rect 12236 28242 12292 28252
rect 12348 30100 12404 30110
rect 12236 28084 12292 28094
rect 11676 28082 12292 28084
rect 11676 28030 12238 28082
rect 12290 28030 12292 28082
rect 11676 28028 12292 28030
rect 12236 28018 12292 28028
rect 11788 27860 11844 27870
rect 12348 27860 12404 30044
rect 12684 29988 12740 29998
rect 12684 29540 12740 29932
rect 12796 29988 12852 29998
rect 12796 29986 12964 29988
rect 12796 29934 12798 29986
rect 12850 29934 12964 29986
rect 12796 29932 12964 29934
rect 12796 29922 12852 29932
rect 12796 29540 12852 29550
rect 12684 29538 12852 29540
rect 12684 29486 12798 29538
rect 12850 29486 12852 29538
rect 12684 29484 12852 29486
rect 12796 29474 12852 29484
rect 11788 27074 11844 27804
rect 11788 27022 11790 27074
rect 11842 27022 11844 27074
rect 11788 27010 11844 27022
rect 12012 27804 12404 27860
rect 12572 29428 12628 29438
rect 12012 27300 12068 27804
rect 11900 26964 11956 26974
rect 11900 26870 11956 26908
rect 11900 26290 11956 26302
rect 11900 26238 11902 26290
rect 11954 26238 11956 26290
rect 11900 26068 11956 26238
rect 11900 26002 11956 26012
rect 12012 25844 12068 27244
rect 12348 27636 12404 27646
rect 12348 27186 12404 27580
rect 12572 27298 12628 29372
rect 12572 27246 12574 27298
rect 12626 27246 12628 27298
rect 12572 27234 12628 27246
rect 12796 28980 12852 28990
rect 12348 27134 12350 27186
rect 12402 27134 12404 27186
rect 12348 27122 12404 27134
rect 12460 26964 12516 26974
rect 12124 26850 12180 26862
rect 12124 26798 12126 26850
rect 12178 26798 12180 26850
rect 12124 26740 12180 26798
rect 12124 26674 12180 26684
rect 12460 26514 12516 26908
rect 12796 26908 12852 28924
rect 12908 28756 12964 29932
rect 12908 28690 12964 28700
rect 13132 28532 13188 30156
rect 13308 29036 13572 29046
rect 13364 28980 13412 29036
rect 13468 28980 13516 29036
rect 13308 28970 13572 28980
rect 13468 28756 13524 28766
rect 13692 28756 13748 31164
rect 13804 30996 13860 31006
rect 13804 30902 13860 30940
rect 14812 30548 14868 30558
rect 14028 30436 14084 30446
rect 13804 30210 13860 30222
rect 13804 30158 13806 30210
rect 13858 30158 13860 30210
rect 13804 29764 13860 30158
rect 14028 29986 14084 30380
rect 14812 30210 14868 30492
rect 15036 30324 15092 34200
rect 16156 30882 16212 34200
rect 17276 31556 17332 34200
rect 17164 31500 17332 31556
rect 16940 31108 16996 31118
rect 16940 31106 17108 31108
rect 16940 31054 16942 31106
rect 16994 31054 17108 31106
rect 16940 31052 17108 31054
rect 16940 31042 16996 31052
rect 16156 30830 16158 30882
rect 16210 30830 16212 30882
rect 16156 30818 16212 30830
rect 15260 30772 15316 30782
rect 15036 30268 15204 30324
rect 14812 30158 14814 30210
rect 14866 30158 14868 30210
rect 14812 30146 14868 30158
rect 14924 30212 14980 30250
rect 14924 30146 14980 30156
rect 15036 30100 15092 30110
rect 15036 30006 15092 30044
rect 14028 29934 14030 29986
rect 14082 29934 14084 29986
rect 14028 29922 14084 29934
rect 14364 29986 14420 29998
rect 14364 29934 14366 29986
rect 14418 29934 14420 29986
rect 14364 29764 14420 29934
rect 15148 29876 15204 30268
rect 13804 29708 14420 29764
rect 15036 29820 15204 29876
rect 15036 29540 15092 29820
rect 15036 29474 15092 29484
rect 14364 29428 14420 29438
rect 13468 28662 13524 28700
rect 13580 28700 13748 28756
rect 14140 29204 14196 29214
rect 13132 28466 13188 28476
rect 13580 28420 13636 28700
rect 14140 28642 14196 29148
rect 14140 28590 14142 28642
rect 14194 28590 14196 28642
rect 13580 28354 13636 28364
rect 13692 28530 13748 28542
rect 13692 28478 13694 28530
rect 13746 28478 13748 28530
rect 13692 28308 13748 28478
rect 13692 28242 13748 28252
rect 13804 28530 13860 28542
rect 13804 28478 13806 28530
rect 13858 28478 13860 28530
rect 13804 28196 13860 28478
rect 13804 28130 13860 28140
rect 14028 28532 14084 28542
rect 13692 27972 13748 27982
rect 13308 27468 13572 27478
rect 13364 27412 13412 27468
rect 13468 27412 13516 27468
rect 13308 27402 13572 27412
rect 12908 27300 12964 27310
rect 12908 27206 12964 27244
rect 13692 27076 13748 27916
rect 13468 27020 13748 27076
rect 13468 26964 13524 27020
rect 12796 26852 13076 26908
rect 13468 26870 13524 26908
rect 12460 26462 12462 26514
rect 12514 26462 12516 26514
rect 12460 26450 12516 26462
rect 12572 26516 12628 26554
rect 12572 26450 12628 26460
rect 12236 26292 12292 26302
rect 11788 25788 12068 25844
rect 12124 26290 12292 26292
rect 12124 26238 12238 26290
rect 12290 26238 12292 26290
rect 12124 26236 12292 26238
rect 11676 25396 11732 25406
rect 11676 25302 11732 25340
rect 11676 24948 11732 24958
rect 11564 24946 11732 24948
rect 11564 24894 11678 24946
rect 11730 24894 11732 24946
rect 11564 24892 11732 24894
rect 11116 24780 11396 24836
rect 10892 24722 10948 24734
rect 10892 24670 10894 24722
rect 10946 24670 10948 24722
rect 10444 24164 10500 24174
rect 10444 23938 10500 24108
rect 10444 23886 10446 23938
rect 10498 23886 10500 23938
rect 10444 23874 10500 23886
rect 10668 23828 10724 23838
rect 10668 23734 10724 23772
rect 10332 22530 10388 22540
rect 10780 23714 10836 23726
rect 10780 23662 10782 23714
rect 10834 23662 10836 23714
rect 10164 20860 10276 20916
rect 10332 21474 10388 21486
rect 10332 21422 10334 21474
rect 10386 21422 10388 21474
rect 10108 20822 10164 20860
rect 10332 20244 10388 21422
rect 10332 20178 10388 20188
rect 10668 20578 10724 20590
rect 10668 20526 10670 20578
rect 10722 20526 10724 20578
rect 9996 19852 10388 19908
rect 10332 19234 10388 19852
rect 10444 19906 10500 19918
rect 10444 19854 10446 19906
rect 10498 19854 10500 19906
rect 10444 19348 10500 19854
rect 10556 19348 10612 19358
rect 10444 19346 10612 19348
rect 10444 19294 10558 19346
rect 10610 19294 10612 19346
rect 10444 19292 10612 19294
rect 10556 19282 10612 19292
rect 10332 19182 10334 19234
rect 10386 19182 10388 19234
rect 10332 19170 10388 19182
rect 10668 19234 10724 20526
rect 10780 19908 10836 23662
rect 10892 23716 10948 24670
rect 11004 23938 11060 24780
rect 11004 23886 11006 23938
rect 11058 23886 11060 23938
rect 11004 23874 11060 23886
rect 11228 23716 11284 23726
rect 10892 23660 11228 23716
rect 11228 23622 11284 23660
rect 10892 23156 10948 23166
rect 10892 22370 10948 23100
rect 11340 22594 11396 24780
rect 11564 23828 11620 23838
rect 11452 23772 11564 23828
rect 11452 22932 11508 23772
rect 11564 23734 11620 23772
rect 11676 23268 11732 24892
rect 11788 23492 11844 25788
rect 12124 25618 12180 26236
rect 12236 26226 12292 26236
rect 12572 26292 12628 26302
rect 12348 26180 12404 26190
rect 12404 26124 12516 26180
rect 12348 26114 12404 26124
rect 12124 25566 12126 25618
rect 12178 25566 12180 25618
rect 12124 25554 12180 25566
rect 12236 26068 12292 26078
rect 11900 25172 11956 25182
rect 11900 24388 11956 25116
rect 12236 24836 12292 26012
rect 12460 25508 12516 26124
rect 11900 23826 11956 24332
rect 11900 23774 11902 23826
rect 11954 23774 11956 23826
rect 11900 23762 11956 23774
rect 12124 24780 12292 24836
rect 12348 25394 12404 25406
rect 12348 25342 12350 25394
rect 12402 25342 12404 25394
rect 12124 23548 12180 24780
rect 12236 24610 12292 24622
rect 12236 24558 12238 24610
rect 12290 24558 12292 24610
rect 12236 23940 12292 24558
rect 12348 24164 12404 25342
rect 12460 24612 12516 25452
rect 12572 25394 12628 26236
rect 12684 26290 12740 26302
rect 12684 26238 12686 26290
rect 12738 26238 12740 26290
rect 12684 25844 12740 26238
rect 13020 26290 13076 26852
rect 13804 26850 13860 26862
rect 13804 26798 13806 26850
rect 13858 26798 13860 26850
rect 13804 26628 13860 26798
rect 13804 26562 13860 26572
rect 14028 26514 14084 28476
rect 14140 27858 14196 28590
rect 14364 28644 14420 29372
rect 14924 29316 14980 29326
rect 14812 29314 14980 29316
rect 14812 29262 14926 29314
rect 14978 29262 14980 29314
rect 14812 29260 14980 29262
rect 14700 28868 14756 28878
rect 14476 28644 14532 28654
rect 14364 28642 14532 28644
rect 14364 28590 14478 28642
rect 14530 28590 14532 28642
rect 14364 28588 14532 28590
rect 14476 28578 14532 28588
rect 14140 27806 14142 27858
rect 14194 27806 14196 27858
rect 14140 27794 14196 27806
rect 14700 28530 14756 28812
rect 14700 28478 14702 28530
rect 14754 28478 14756 28530
rect 14140 27412 14196 27422
rect 14140 27298 14196 27356
rect 14140 27246 14142 27298
rect 14194 27246 14196 27298
rect 14140 27234 14196 27246
rect 14252 27300 14308 27310
rect 14252 27076 14308 27244
rect 14700 27188 14756 28478
rect 14812 27412 14868 29260
rect 14924 29250 14980 29260
rect 15036 28756 15092 28766
rect 15036 28642 15092 28700
rect 15036 28590 15038 28642
rect 15090 28590 15092 28642
rect 15036 28578 15092 28590
rect 15148 28084 15204 28094
rect 15148 27990 15204 28028
rect 14812 27346 14868 27356
rect 14588 27132 15204 27188
rect 14252 27010 14308 27020
rect 14476 27074 14532 27086
rect 14476 27022 14478 27074
rect 14530 27022 14532 27074
rect 14476 26852 14532 27022
rect 14588 27074 14644 27132
rect 14588 27022 14590 27074
rect 14642 27022 14644 27074
rect 14588 27010 14644 27022
rect 14812 26964 14868 27002
rect 14812 26898 14868 26908
rect 14700 26852 14756 26862
rect 14476 26796 14644 26852
rect 14028 26462 14030 26514
rect 14082 26462 14084 26514
rect 14028 26450 14084 26462
rect 14140 26740 14196 26750
rect 13020 26238 13022 26290
rect 13074 26238 13076 26290
rect 13020 26226 13076 26238
rect 14028 26292 14084 26302
rect 13308 25900 13572 25910
rect 13364 25844 13412 25900
rect 13468 25844 13516 25900
rect 13308 25834 13572 25844
rect 13916 25844 13972 25854
rect 12684 25778 12740 25788
rect 12572 25342 12574 25394
rect 12626 25342 12628 25394
rect 12684 25620 12740 25630
rect 12684 25450 12740 25564
rect 12684 25398 12686 25450
rect 12738 25398 12740 25450
rect 13916 25506 13972 25788
rect 13916 25454 13918 25506
rect 13970 25454 13972 25506
rect 13916 25442 13972 25454
rect 12684 25386 12740 25398
rect 12908 25394 12964 25406
rect 12572 25330 12628 25342
rect 12908 25342 12910 25394
rect 12962 25342 12964 25394
rect 12908 25284 12964 25342
rect 12684 25228 12964 25284
rect 13692 25394 13748 25406
rect 13692 25342 13694 25394
rect 13746 25342 13748 25394
rect 12572 24948 12628 24958
rect 12572 24854 12628 24892
rect 12684 24946 12740 25228
rect 13244 25060 13300 25070
rect 13020 24948 13076 24958
rect 12684 24894 12686 24946
rect 12738 24894 12740 24946
rect 12684 24882 12740 24894
rect 12796 24892 13020 24948
rect 12796 24834 12852 24892
rect 13020 24882 13076 24892
rect 13244 24946 13300 25004
rect 13244 24894 13246 24946
rect 13298 24894 13300 24946
rect 13244 24882 13300 24894
rect 13356 24948 13412 24958
rect 13356 24854 13412 24892
rect 12796 24782 12798 24834
rect 12850 24782 12852 24834
rect 12796 24770 12852 24782
rect 13468 24836 13524 24874
rect 13468 24770 13524 24780
rect 13132 24722 13188 24734
rect 13132 24670 13134 24722
rect 13186 24670 13188 24722
rect 13132 24612 13188 24670
rect 12460 24556 12628 24612
rect 12348 24098 12404 24108
rect 12236 23884 12516 23940
rect 12236 23716 12292 23726
rect 12236 23622 12292 23660
rect 11788 23426 11844 23436
rect 11900 23492 12180 23548
rect 12236 23492 12292 23502
rect 11900 23268 11956 23492
rect 11676 23202 11732 23212
rect 11788 23212 11956 23268
rect 11564 23156 11620 23166
rect 11564 23062 11620 23100
rect 11452 22866 11508 22876
rect 11340 22542 11342 22594
rect 11394 22542 11396 22594
rect 11340 22530 11396 22542
rect 10892 22318 10894 22370
rect 10946 22318 10948 22370
rect 10892 22306 10948 22318
rect 11452 22258 11508 22270
rect 11452 22206 11454 22258
rect 11506 22206 11508 22258
rect 11340 22148 11396 22158
rect 11228 22146 11396 22148
rect 11228 22094 11342 22146
rect 11394 22094 11396 22146
rect 11228 22092 11396 22094
rect 11116 21588 11172 21598
rect 11004 20690 11060 20702
rect 11004 20638 11006 20690
rect 11058 20638 11060 20690
rect 10892 20578 10948 20590
rect 10892 20526 10894 20578
rect 10946 20526 10948 20578
rect 10892 20132 10948 20526
rect 10892 20066 10948 20076
rect 10780 19842 10836 19852
rect 10668 19182 10670 19234
rect 10722 19182 10724 19234
rect 10668 19170 10724 19182
rect 10892 19234 10948 19246
rect 10892 19182 10894 19234
rect 10946 19182 10948 19234
rect 9660 18498 9716 18508
rect 9772 18508 9940 18564
rect 9212 17614 9214 17666
rect 9266 17614 9268 17666
rect 9212 17602 9268 17614
rect 8204 17106 8372 17108
rect 8204 17054 8206 17106
rect 8258 17054 8372 17106
rect 8204 17052 8372 17054
rect 8540 17556 8596 17566
rect 8204 17042 8260 17052
rect 7868 16996 7924 17006
rect 7868 16902 7924 16940
rect 7980 16996 8036 17006
rect 8428 16996 8484 17006
rect 7980 16994 8148 16996
rect 7980 16942 7982 16994
rect 8034 16942 8148 16994
rect 7980 16940 8148 16942
rect 7980 16930 8036 16940
rect 7308 14242 7364 14252
rect 7420 15932 7812 15988
rect 7196 14196 7252 14206
rect 6860 14140 7196 14196
rect 6860 13858 6916 14140
rect 7196 14130 7252 14140
rect 6860 13806 6862 13858
rect 6914 13806 6916 13858
rect 6860 13794 6916 13806
rect 6748 12786 6804 12796
rect 7308 12180 7364 12190
rect 6748 12178 7364 12180
rect 6748 12126 7310 12178
rect 7362 12126 7364 12178
rect 6748 12124 7364 12126
rect 6188 11342 6190 11394
rect 6242 11342 6244 11394
rect 3724 11060 3780 11070
rect 3612 10722 3668 10734
rect 3612 10670 3614 10722
rect 3666 10670 3668 10722
rect 2828 10612 2884 10622
rect 3388 10612 3444 10622
rect 2828 9826 2884 10556
rect 2828 9774 2830 9826
rect 2882 9774 2884 9826
rect 2828 9762 2884 9774
rect 3164 10610 3444 10612
rect 3164 10558 3390 10610
rect 3442 10558 3444 10610
rect 3164 10556 3444 10558
rect 3164 9826 3220 10556
rect 3388 10546 3444 10556
rect 3388 9828 3444 9838
rect 3164 9774 3166 9826
rect 3218 9774 3220 9826
rect 3164 9762 3220 9774
rect 3276 9826 3444 9828
rect 3276 9774 3390 9826
rect 3442 9774 3444 9826
rect 3276 9772 3444 9774
rect 3276 9716 3332 9772
rect 3388 9762 3444 9772
rect 2492 9602 2548 9614
rect 2492 9550 2494 9602
rect 2546 9550 2548 9602
rect 1708 8930 1764 8942
rect 1708 8878 1710 8930
rect 1762 8878 1764 8930
rect 1708 8820 1764 8878
rect 1708 8754 1764 8764
rect 2492 8428 2548 9550
rect 2156 8372 2212 8382
rect 1820 8260 1876 8270
rect 1820 8166 1876 8204
rect 2044 7924 2100 7934
rect 2044 7474 2100 7868
rect 2044 7422 2046 7474
rect 2098 7422 2100 7474
rect 2044 7410 2100 7422
rect 2156 7700 2212 8316
rect 2380 8372 2548 8428
rect 2716 9602 2772 9614
rect 2716 9550 2718 9602
rect 2770 9550 2772 9602
rect 2716 8372 2772 9550
rect 2380 7812 2436 8372
rect 2716 8306 2772 8316
rect 2492 8148 2548 8158
rect 3164 8148 3220 8158
rect 2492 8146 3108 8148
rect 2492 8094 2494 8146
rect 2546 8094 3108 8146
rect 2492 8092 3108 8094
rect 2492 8082 2548 8092
rect 2380 7756 2884 7812
rect 1708 5794 1764 5806
rect 1708 5742 1710 5794
rect 1762 5742 1764 5794
rect 1708 5684 1764 5742
rect 2156 5684 2212 7644
rect 2492 7588 2548 7598
rect 2492 7494 2548 7532
rect 1708 5628 2212 5684
rect 1708 5460 1764 5470
rect 1708 4226 1764 5404
rect 2044 5460 2100 5470
rect 1708 4174 1710 4226
rect 1762 4174 1764 4226
rect 1708 4162 1764 4174
rect 1932 5012 1988 5022
rect 924 3556 980 3566
rect 1932 3556 1988 4956
rect 2044 5010 2100 5404
rect 2044 4958 2046 5010
rect 2098 4958 2100 5010
rect 2044 4946 2100 4958
rect 924 800 980 3500
rect 1820 3500 1988 3556
rect 2156 3556 2212 5628
rect 2380 7474 2436 7486
rect 2380 7422 2382 7474
rect 2434 7422 2436 7474
rect 2380 6580 2436 7422
rect 2604 7474 2660 7486
rect 2604 7422 2606 7474
rect 2658 7422 2660 7474
rect 2604 7252 2660 7422
rect 2828 7474 2884 7756
rect 3052 7698 3108 8092
rect 3052 7646 3054 7698
rect 3106 7646 3108 7698
rect 3052 7634 3108 7646
rect 2828 7422 2830 7474
rect 2882 7422 2884 7474
rect 2828 7410 2884 7422
rect 2604 7186 2660 7196
rect 2380 5460 2436 6524
rect 2380 5394 2436 5404
rect 2268 5348 2324 5358
rect 2268 5122 2324 5292
rect 2716 5236 2772 5246
rect 2268 5070 2270 5122
rect 2322 5070 2324 5122
rect 2268 5058 2324 5070
rect 2492 5234 2772 5236
rect 2492 5182 2718 5234
rect 2770 5182 2772 5234
rect 2492 5180 2772 5182
rect 2380 3556 2436 3566
rect 2156 3554 2436 3556
rect 2156 3502 2382 3554
rect 2434 3502 2436 3554
rect 2156 3500 2436 3502
rect 1820 3442 1876 3500
rect 2380 3490 2436 3500
rect 2044 3444 2100 3454
rect 1820 3390 1822 3442
rect 1874 3390 1876 3442
rect 1820 3378 1876 3390
rect 1932 3388 2044 3444
rect 1932 3330 1988 3388
rect 2044 3378 2100 3388
rect 1932 3278 1934 3330
rect 1986 3278 1988 3330
rect 1932 3266 1988 3278
rect 2156 3332 2212 3342
rect 2156 3238 2212 3276
rect 2492 800 2548 5180
rect 2716 5170 2772 5180
rect 3164 3332 3220 8092
rect 3276 7586 3332 9660
rect 3388 9602 3444 9614
rect 3388 9550 3390 9602
rect 3442 9550 3444 9602
rect 3388 9156 3444 9550
rect 3612 9380 3668 10670
rect 3724 10612 3780 11004
rect 4508 10836 4564 10846
rect 4508 10742 4564 10780
rect 5404 10836 5460 10846
rect 5964 10836 6020 10846
rect 5404 10834 5684 10836
rect 5404 10782 5406 10834
rect 5458 10782 5684 10834
rect 5404 10780 5684 10782
rect 5404 10770 5460 10780
rect 3724 10518 3780 10556
rect 5516 10610 5572 10622
rect 5516 10558 5518 10610
rect 5570 10558 5572 10610
rect 4844 10498 4900 10510
rect 4844 10446 4846 10498
rect 4898 10446 4900 10498
rect 4844 10052 4900 10446
rect 5516 10500 5572 10558
rect 5628 10612 5684 10780
rect 5964 10742 6020 10780
rect 5628 10556 5908 10612
rect 5516 10444 5796 10500
rect 5404 10388 5460 10426
rect 5404 10322 5460 10332
rect 5740 10386 5796 10444
rect 5740 10334 5742 10386
rect 5794 10334 5796 10386
rect 5740 10322 5796 10334
rect 5244 10220 5508 10230
rect 5300 10164 5348 10220
rect 5404 10164 5452 10220
rect 5244 10154 5508 10164
rect 5516 10052 5572 10062
rect 4900 9996 5124 10052
rect 3724 9828 3780 9838
rect 4172 9828 4228 9838
rect 3724 9826 4228 9828
rect 3724 9774 3726 9826
rect 3778 9774 4174 9826
rect 4226 9774 4228 9826
rect 3724 9772 4228 9774
rect 3724 9762 3780 9772
rect 4172 9762 4228 9772
rect 4732 9828 4788 9838
rect 4844 9828 4900 9996
rect 5068 9938 5124 9996
rect 5068 9886 5070 9938
rect 5122 9886 5124 9938
rect 5068 9874 5124 9886
rect 4732 9826 4900 9828
rect 4732 9774 4734 9826
rect 4786 9774 4900 9826
rect 4732 9772 4900 9774
rect 4732 9762 4788 9772
rect 4060 9604 4116 9614
rect 4060 9510 4116 9548
rect 4284 9602 4340 9614
rect 4284 9550 4286 9602
rect 4338 9550 4340 9602
rect 3612 9324 4004 9380
rect 3836 9156 3892 9166
rect 3388 9154 3892 9156
rect 3388 9102 3838 9154
rect 3890 9102 3892 9154
rect 3388 9100 3892 9102
rect 3836 9090 3892 9100
rect 3276 7534 3278 7586
rect 3330 7534 3332 7586
rect 3276 7522 3332 7534
rect 3500 8932 3556 8942
rect 3500 7586 3556 8876
rect 3948 8708 4004 9324
rect 3948 8642 4004 8652
rect 4284 8820 4340 9550
rect 4956 9604 5012 9614
rect 4956 9266 5012 9548
rect 4956 9214 4958 9266
rect 5010 9214 5012 9266
rect 4956 9202 5012 9214
rect 4620 9156 4676 9166
rect 4620 9044 4676 9100
rect 4284 8372 4340 8764
rect 4060 8316 4340 8372
rect 4508 9042 4676 9044
rect 4508 8990 4622 9042
rect 4674 8990 4676 9042
rect 4508 8988 4676 8990
rect 3500 7534 3502 7586
rect 3554 7534 3556 7586
rect 3500 7522 3556 7534
rect 3836 7924 3892 7934
rect 3836 7474 3892 7868
rect 3836 7422 3838 7474
rect 3890 7422 3892 7474
rect 3836 6916 3892 7422
rect 3836 6850 3892 6860
rect 4060 6690 4116 8316
rect 4508 8260 4564 8988
rect 4620 8978 4676 8988
rect 5180 9042 5236 9054
rect 5180 8990 5182 9042
rect 5234 8990 5236 9042
rect 5068 8932 5124 8942
rect 5068 8838 5124 8876
rect 4396 8036 4452 8046
rect 4172 7700 4228 7710
rect 4172 7606 4228 7644
rect 4396 7698 4452 7980
rect 4396 7646 4398 7698
rect 4450 7646 4452 7698
rect 4284 7476 4340 7486
rect 4284 7382 4340 7420
rect 4396 7252 4452 7646
rect 4396 7186 4452 7196
rect 4060 6638 4062 6690
rect 4114 6638 4116 6690
rect 4060 6626 4116 6638
rect 3276 6466 3332 6478
rect 3276 6414 3278 6466
rect 3330 6414 3332 6466
rect 3276 3556 3332 6414
rect 3836 6468 3892 6478
rect 3836 6018 3892 6412
rect 3836 5966 3838 6018
rect 3890 5966 3892 6018
rect 3836 5954 3892 5966
rect 4508 5906 4564 8204
rect 4508 5854 4510 5906
rect 4562 5854 4564 5906
rect 3836 5684 3892 5694
rect 3836 4450 3892 5628
rect 3836 4398 3838 4450
rect 3890 4398 3892 4450
rect 3836 4386 3892 4398
rect 4508 4340 4564 5854
rect 4620 8820 4676 8830
rect 4620 8370 4676 8764
rect 5180 8820 5236 8990
rect 5516 9042 5572 9996
rect 5740 9828 5796 9838
rect 5740 9734 5796 9772
rect 5516 8990 5518 9042
rect 5570 8990 5572 9042
rect 5516 8978 5572 8990
rect 5852 8932 5908 10556
rect 6076 9604 6132 9614
rect 6076 9510 6132 9548
rect 6188 9156 6244 11342
rect 6412 11396 6468 11406
rect 6412 10836 6468 11340
rect 6412 9828 6468 10780
rect 6748 10722 6804 12124
rect 7308 12114 7364 12124
rect 6860 11282 6916 11294
rect 6860 11230 6862 11282
rect 6914 11230 6916 11282
rect 6860 10834 6916 11230
rect 7420 10948 7476 15932
rect 7644 15540 7700 15550
rect 8092 15540 8148 16940
rect 8428 16902 8484 16940
rect 8204 15540 8260 15550
rect 7644 15538 8260 15540
rect 7644 15486 7646 15538
rect 7698 15486 8206 15538
rect 8258 15486 8260 15538
rect 7644 15484 8260 15486
rect 7644 15474 7700 15484
rect 7532 15314 7588 15326
rect 7532 15262 7534 15314
rect 7586 15262 7588 15314
rect 7532 15204 7588 15262
rect 7532 15138 7588 15148
rect 7868 15314 7924 15326
rect 7868 15262 7870 15314
rect 7922 15262 7924 15314
rect 7644 14532 7700 14542
rect 7644 14438 7700 14476
rect 7868 14530 7924 15262
rect 7980 15316 8036 15326
rect 7980 15222 8036 15260
rect 8204 15148 8260 15484
rect 8316 15428 8372 15438
rect 8316 15334 8372 15372
rect 8204 15092 8484 15148
rect 7868 14478 7870 14530
rect 7922 14478 7924 14530
rect 7868 14466 7924 14478
rect 8092 14420 8148 14430
rect 8316 14420 8372 14430
rect 8092 14418 8372 14420
rect 8092 14366 8094 14418
rect 8146 14366 8318 14418
rect 8370 14366 8372 14418
rect 8092 14364 8372 14366
rect 8092 14354 8148 14364
rect 8316 14354 8372 14364
rect 7868 14306 7924 14318
rect 7868 14254 7870 14306
rect 7922 14254 7924 14306
rect 7868 14196 7924 14254
rect 7868 14130 7924 14140
rect 8428 13636 8484 15092
rect 8540 14532 8596 17500
rect 9276 17276 9540 17286
rect 9332 17220 9380 17276
rect 9436 17220 9484 17276
rect 9276 17210 9540 17220
rect 8764 17108 8820 17118
rect 9660 17108 9716 17118
rect 9772 17108 9828 18508
rect 10892 18450 10948 19182
rect 11004 19124 11060 20638
rect 11116 20468 11172 21532
rect 11228 20580 11284 22092
rect 11340 22082 11396 22092
rect 11452 22036 11508 22206
rect 11788 22258 11844 23212
rect 12012 23156 12068 23166
rect 11788 22206 11790 22258
rect 11842 22206 11844 22258
rect 11788 22194 11844 22206
rect 11900 23100 12012 23156
rect 11340 21812 11396 21822
rect 11452 21812 11508 21980
rect 11340 21810 11508 21812
rect 11340 21758 11342 21810
rect 11394 21758 11508 21810
rect 11340 21756 11508 21758
rect 11340 21746 11396 21756
rect 11900 20916 11956 23100
rect 12012 23090 12068 23100
rect 12124 22146 12180 22158
rect 12124 22094 12126 22146
rect 12178 22094 12180 22146
rect 12124 21586 12180 22094
rect 12236 21700 12292 23436
rect 12348 23268 12404 23278
rect 12348 23174 12404 23212
rect 12236 21634 12292 21644
rect 12124 21534 12126 21586
rect 12178 21534 12180 21586
rect 12012 20916 12068 20926
rect 11900 20914 12068 20916
rect 11900 20862 12014 20914
rect 12066 20862 12068 20914
rect 11900 20860 12068 20862
rect 12012 20850 12068 20860
rect 11228 20514 11284 20524
rect 11564 20578 11620 20590
rect 11564 20526 11566 20578
rect 11618 20526 11620 20578
rect 11116 20402 11172 20412
rect 11564 20468 11620 20526
rect 11564 20402 11620 20412
rect 11004 19058 11060 19068
rect 11452 20132 11508 20142
rect 11452 19122 11508 20076
rect 11452 19070 11454 19122
rect 11506 19070 11508 19122
rect 11452 19058 11508 19070
rect 11564 19124 11620 19134
rect 11564 19030 11620 19068
rect 11228 19010 11284 19022
rect 11228 18958 11230 19010
rect 11282 18958 11284 19010
rect 11228 18564 11284 18958
rect 11676 19012 11732 19022
rect 11340 18564 11396 18574
rect 11228 18562 11396 18564
rect 11228 18510 11342 18562
rect 11394 18510 11396 18562
rect 11228 18508 11396 18510
rect 11340 18498 11396 18508
rect 11676 18562 11732 18956
rect 12124 18900 12180 21534
rect 12460 21476 12516 23884
rect 12572 23826 12628 24556
rect 12572 23774 12574 23826
rect 12626 23774 12628 23826
rect 12572 23762 12628 23774
rect 12684 24556 13188 24612
rect 12684 23044 12740 24556
rect 13308 24332 13572 24342
rect 13364 24276 13412 24332
rect 13468 24276 13516 24332
rect 13308 24266 13572 24276
rect 13692 23940 13748 25342
rect 13804 24724 13860 24734
rect 13804 24276 13860 24668
rect 13916 24722 13972 24734
rect 13916 24670 13918 24722
rect 13970 24670 13972 24722
rect 13916 24500 13972 24670
rect 13916 24434 13972 24444
rect 13804 24210 13860 24220
rect 13468 23884 13748 23940
rect 12572 22260 12628 22270
rect 12684 22260 12740 22988
rect 12908 23714 12964 23726
rect 12908 23662 12910 23714
rect 12962 23662 12964 23714
rect 12908 22484 12964 23662
rect 13468 23380 13524 23884
rect 13916 23828 13972 23838
rect 14028 23828 14084 26236
rect 14140 25956 14196 26684
rect 14140 25900 14420 25956
rect 14140 25732 14196 25742
rect 14140 25284 14196 25676
rect 14252 25508 14308 25518
rect 14364 25508 14420 25900
rect 14588 25732 14644 26796
rect 14700 26758 14756 26796
rect 14588 25666 14644 25676
rect 14812 26740 14868 26750
rect 14476 25508 14532 25518
rect 14364 25506 14532 25508
rect 14364 25454 14478 25506
rect 14530 25454 14532 25506
rect 14364 25452 14532 25454
rect 14252 25414 14308 25452
rect 14140 25228 14308 25284
rect 14252 24836 14308 25228
rect 14476 24948 14532 25452
rect 14588 25396 14644 25406
rect 14588 25282 14644 25340
rect 14588 25230 14590 25282
rect 14642 25230 14644 25282
rect 14588 25218 14644 25230
rect 14476 24882 14532 24892
rect 14364 24836 14420 24846
rect 14252 24834 14420 24836
rect 14252 24782 14366 24834
rect 14418 24782 14420 24834
rect 14252 24780 14420 24782
rect 13916 23826 14084 23828
rect 13916 23774 13918 23826
rect 13970 23774 14084 23826
rect 13916 23772 14084 23774
rect 14140 24724 14196 24734
rect 13916 23762 13972 23772
rect 13580 23716 13636 23726
rect 14140 23716 14196 24668
rect 14364 24388 14420 24780
rect 14364 24322 14420 24332
rect 14588 24722 14644 24734
rect 14588 24670 14590 24722
rect 14642 24670 14644 24722
rect 13580 23714 13748 23716
rect 13580 23662 13582 23714
rect 13634 23662 13748 23714
rect 13580 23660 13748 23662
rect 13580 23650 13636 23660
rect 12908 22370 12964 22428
rect 12908 22318 12910 22370
rect 12962 22318 12964 22370
rect 12908 22306 12964 22318
rect 13132 23324 13524 23380
rect 12572 22258 12740 22260
rect 12572 22206 12574 22258
rect 12626 22206 12740 22258
rect 12572 22204 12740 22206
rect 12572 22194 12628 22204
rect 12908 21812 12964 21822
rect 13132 21812 13188 23324
rect 13692 23156 13748 23660
rect 13308 22764 13572 22774
rect 13364 22708 13412 22764
rect 13468 22708 13516 22764
rect 13308 22698 13572 22708
rect 13580 22596 13636 22606
rect 13468 22258 13524 22270
rect 13468 22206 13470 22258
rect 13522 22206 13524 22258
rect 13244 21812 13300 21822
rect 13132 21810 13300 21812
rect 13132 21758 13246 21810
rect 13298 21758 13300 21810
rect 13132 21756 13300 21758
rect 12572 21700 12628 21710
rect 12572 21586 12628 21644
rect 12908 21698 12964 21756
rect 13244 21746 13300 21756
rect 12908 21646 12910 21698
rect 12962 21646 12964 21698
rect 12908 21634 12964 21646
rect 13020 21698 13076 21710
rect 13020 21646 13022 21698
rect 13074 21646 13076 21698
rect 12572 21534 12574 21586
rect 12626 21534 12628 21586
rect 12572 21522 12628 21534
rect 12460 21410 12516 21420
rect 12124 18834 12180 18844
rect 12236 20580 12292 20590
rect 11788 18676 11844 18686
rect 11788 18582 11844 18620
rect 12012 18676 12068 18686
rect 12068 18620 12180 18676
rect 12012 18610 12068 18620
rect 11676 18510 11678 18562
rect 11730 18510 11732 18562
rect 11676 18498 11732 18510
rect 10892 18398 10894 18450
rect 10946 18398 10948 18450
rect 9884 18340 9940 18350
rect 9884 17778 9940 18284
rect 9884 17726 9886 17778
rect 9938 17726 9940 17778
rect 9884 17714 9940 17726
rect 10892 18228 10948 18398
rect 11116 18452 11172 18462
rect 11116 18358 11172 18396
rect 12012 18452 12068 18462
rect 12012 18358 12068 18396
rect 11228 18340 11284 18350
rect 11228 18246 11284 18284
rect 8764 17106 9828 17108
rect 8764 17054 8766 17106
rect 8818 17054 9662 17106
rect 9714 17054 9828 17106
rect 8764 17052 9828 17054
rect 10668 17444 10724 17454
rect 8764 17042 8820 17052
rect 9660 17042 9716 17052
rect 10668 16884 10724 17388
rect 10892 17106 10948 18172
rect 12012 17780 12068 17790
rect 12124 17780 12180 18620
rect 12012 17778 12180 17780
rect 12012 17726 12014 17778
rect 12066 17726 12180 17778
rect 12012 17724 12180 17726
rect 12012 17714 12068 17724
rect 10892 17054 10894 17106
rect 10946 17054 10948 17106
rect 10892 17042 10948 17054
rect 11340 17668 11396 17678
rect 11228 16996 11284 17006
rect 11004 16994 11284 16996
rect 11004 16942 11230 16994
rect 11282 16942 11284 16994
rect 11004 16940 11284 16942
rect 11004 16884 11060 16940
rect 11228 16930 11284 16940
rect 10668 16882 11060 16884
rect 10668 16830 10670 16882
rect 10722 16830 11060 16882
rect 10668 16828 11060 16830
rect 10668 16818 10724 16828
rect 10892 16100 10948 16110
rect 10892 16006 10948 16044
rect 11340 15986 11396 17612
rect 12236 17556 12292 20524
rect 13020 20356 13076 21646
rect 13468 21588 13524 22206
rect 13580 21812 13636 22540
rect 13692 21924 13748 23100
rect 13804 22484 13860 22494
rect 13804 22258 13860 22428
rect 13804 22206 13806 22258
rect 13858 22206 13860 22258
rect 13804 22194 13860 22206
rect 14140 22258 14196 23660
rect 14252 23714 14308 23726
rect 14252 23662 14254 23714
rect 14306 23662 14308 23714
rect 14252 23548 14308 23662
rect 14252 23492 14532 23548
rect 14140 22206 14142 22258
rect 14194 22206 14196 22258
rect 14140 22194 14196 22206
rect 14252 23156 14308 23166
rect 13692 21858 13748 21868
rect 14028 22148 14084 22158
rect 13580 21746 13636 21756
rect 13468 21522 13524 21532
rect 13692 21476 13748 21486
rect 14028 21476 14084 22092
rect 14140 21586 14196 21598
rect 14140 21534 14142 21586
rect 14194 21534 14196 21586
rect 14140 21476 14196 21534
rect 13692 21474 14196 21476
rect 13692 21422 13694 21474
rect 13746 21422 14196 21474
rect 13692 21420 14196 21422
rect 13692 21410 13748 21420
rect 13308 21196 13572 21206
rect 13364 21140 13412 21196
rect 13468 21140 13516 21196
rect 13308 21130 13572 21140
rect 13804 21028 13860 21038
rect 12572 20300 13076 20356
rect 13468 20916 13524 20926
rect 13468 20802 13524 20860
rect 13468 20750 13470 20802
rect 13522 20750 13524 20802
rect 12572 20132 12628 20300
rect 13468 20188 13524 20750
rect 13020 20132 13524 20188
rect 13692 20132 13748 20142
rect 12572 19906 12628 20076
rect 12572 19854 12574 19906
rect 12626 19854 12628 19906
rect 12572 19842 12628 19854
rect 12908 20130 13076 20132
rect 12908 20078 13022 20130
rect 13074 20078 13076 20130
rect 12908 20076 13076 20078
rect 12908 20020 12964 20076
rect 13020 20066 13076 20076
rect 13692 20038 13748 20076
rect 12908 19348 12964 19964
rect 13580 20018 13636 20030
rect 13580 19966 13582 20018
rect 13634 19966 13636 20018
rect 13580 19796 13636 19966
rect 13580 19740 13748 19796
rect 13308 19628 13572 19638
rect 13364 19572 13412 19628
rect 13468 19572 13516 19628
rect 13308 19562 13572 19572
rect 12236 17490 12292 17500
rect 12348 19124 12404 19134
rect 12348 17554 12404 19068
rect 12348 17502 12350 17554
rect 12402 17502 12404 17554
rect 12348 17490 12404 17502
rect 12460 17668 12516 17678
rect 12460 17332 12516 17612
rect 12908 17668 12964 19292
rect 13580 19236 13636 19246
rect 13692 19236 13748 19740
rect 13020 19234 13748 19236
rect 13020 19182 13582 19234
rect 13634 19182 13748 19234
rect 13020 19180 13748 19182
rect 13020 19124 13076 19180
rect 13580 19170 13636 19180
rect 13020 18562 13076 19068
rect 13692 19010 13748 19022
rect 13692 18958 13694 19010
rect 13746 18958 13748 19010
rect 13692 18900 13748 18958
rect 13692 18834 13748 18844
rect 13132 18676 13188 18686
rect 13132 18582 13188 18620
rect 13804 18676 13860 20972
rect 14140 20188 14196 21420
rect 14252 20916 14308 23100
rect 14476 22260 14532 23492
rect 14588 22484 14644 24670
rect 14812 24724 14868 26684
rect 15148 25956 15204 27132
rect 15260 26516 15316 30716
rect 15372 30548 15428 30558
rect 15372 27300 15428 30492
rect 16492 30436 16548 30446
rect 15708 30212 15764 30222
rect 15484 30210 15764 30212
rect 15484 30158 15710 30210
rect 15762 30158 15764 30210
rect 15484 30156 15764 30158
rect 15484 28644 15540 30156
rect 15708 30146 15764 30156
rect 16492 30210 16548 30380
rect 16492 30158 16494 30210
rect 16546 30158 16548 30210
rect 16492 30146 16548 30158
rect 16940 29988 16996 29998
rect 15932 29652 15988 29662
rect 15708 29540 15764 29550
rect 15708 29426 15764 29484
rect 15932 29538 15988 29596
rect 15932 29486 15934 29538
rect 15986 29486 15988 29538
rect 15932 29474 15988 29486
rect 16492 29652 16548 29662
rect 15708 29374 15710 29426
rect 15762 29374 15764 29426
rect 15708 29204 15764 29374
rect 15708 29138 15764 29148
rect 15820 29426 15876 29438
rect 15820 29374 15822 29426
rect 15874 29374 15876 29426
rect 15820 28868 15876 29374
rect 16156 29428 16212 29438
rect 16156 29334 16212 29372
rect 15820 28802 15876 28812
rect 16044 29092 16100 29102
rect 15484 28550 15540 28588
rect 15372 27244 15652 27300
rect 15260 26450 15316 26460
rect 15372 26068 15428 26078
rect 15428 26012 15540 26068
rect 15372 26002 15428 26012
rect 15148 25890 15204 25900
rect 15372 25844 15428 25854
rect 15260 25620 15316 25630
rect 14924 25394 14980 25406
rect 14924 25342 14926 25394
rect 14978 25342 14980 25394
rect 14924 24948 14980 25342
rect 15036 25396 15092 25406
rect 15148 25396 15204 25406
rect 15092 25394 15204 25396
rect 15092 25342 15150 25394
rect 15202 25342 15204 25394
rect 15092 25340 15204 25342
rect 15036 25330 15092 25340
rect 15148 25330 15204 25340
rect 14924 24892 15092 24948
rect 14924 24724 14980 24734
rect 14812 24722 14980 24724
rect 14812 24670 14926 24722
rect 14978 24670 14980 24722
rect 14812 24668 14980 24670
rect 14924 24658 14980 24668
rect 15036 24500 15092 24892
rect 14812 24444 15092 24500
rect 15148 24836 15204 24846
rect 14588 22418 14644 22428
rect 14700 23714 14756 23726
rect 14700 23662 14702 23714
rect 14754 23662 14756 23714
rect 14700 23380 14756 23662
rect 14476 22166 14532 22204
rect 14700 22148 14756 23324
rect 14812 22932 14868 24444
rect 15036 24276 15092 24286
rect 14812 22866 14868 22876
rect 14924 24164 14980 24174
rect 14812 22708 14868 22718
rect 14812 22482 14868 22652
rect 14812 22430 14814 22482
rect 14866 22430 14868 22482
rect 14812 22418 14868 22430
rect 14700 22082 14756 22092
rect 14364 21812 14420 21822
rect 14924 21812 14980 24108
rect 15036 23940 15092 24220
rect 15036 23826 15092 23884
rect 15036 23774 15038 23826
rect 15090 23774 15092 23826
rect 15036 23762 15092 23774
rect 15036 23156 15092 23166
rect 15036 22594 15092 23100
rect 15036 22542 15038 22594
rect 15090 22542 15092 22594
rect 15036 22036 15092 22542
rect 15148 22596 15204 24780
rect 15260 24612 15316 25564
rect 15372 25506 15428 25788
rect 15484 25618 15540 26012
rect 15484 25566 15486 25618
rect 15538 25566 15540 25618
rect 15484 25554 15540 25566
rect 15372 25454 15374 25506
rect 15426 25454 15428 25506
rect 15372 25442 15428 25454
rect 15484 25282 15540 25294
rect 15484 25230 15486 25282
rect 15538 25230 15540 25282
rect 15484 25172 15540 25230
rect 15484 25106 15540 25116
rect 15484 24948 15540 24958
rect 15596 24948 15652 27244
rect 15708 27074 15764 27086
rect 15708 27022 15710 27074
rect 15762 27022 15764 27074
rect 15708 25620 15764 27022
rect 15708 25554 15764 25564
rect 15820 26964 15876 26974
rect 15820 25506 15876 26908
rect 15932 26740 15988 26750
rect 15932 26402 15988 26684
rect 15932 26350 15934 26402
rect 15986 26350 15988 26402
rect 15932 26338 15988 26350
rect 15820 25454 15822 25506
rect 15874 25454 15876 25506
rect 15820 25442 15876 25454
rect 15932 25732 15988 25742
rect 15932 25284 15988 25676
rect 16044 25508 16100 29036
rect 16492 29092 16548 29596
rect 16604 29202 16660 29214
rect 16604 29150 16606 29202
rect 16658 29150 16660 29202
rect 16604 29092 16660 29150
rect 16940 29092 16996 29932
rect 16604 29036 16996 29092
rect 16492 29026 16548 29036
rect 16156 28530 16212 28542
rect 16156 28478 16158 28530
rect 16210 28478 16212 28530
rect 16156 26516 16212 28478
rect 16828 28532 16884 28542
rect 16828 27186 16884 28476
rect 16828 27134 16830 27186
rect 16882 27134 16884 27186
rect 16828 27122 16884 27134
rect 16940 27076 16996 29036
rect 17052 27860 17108 31052
rect 17164 28084 17220 31500
rect 17340 31388 17604 31398
rect 17396 31332 17444 31388
rect 17500 31332 17548 31388
rect 17340 31322 17604 31332
rect 18396 31220 18452 34200
rect 18620 31220 18676 31230
rect 18396 31218 18676 31220
rect 18396 31166 18622 31218
rect 18674 31166 18676 31218
rect 18396 31164 18676 31166
rect 18620 31154 18676 31164
rect 19516 31220 19572 34200
rect 20636 33124 20692 34200
rect 20636 33058 20692 33068
rect 20748 32116 20804 32126
rect 20804 32060 20916 32116
rect 20748 32050 20804 32060
rect 19516 31154 19572 31164
rect 19628 32004 19684 32014
rect 19628 31556 19684 31948
rect 17276 30994 17332 31006
rect 17276 30942 17278 30994
rect 17330 30942 17332 30994
rect 17276 29988 17332 30942
rect 17948 30994 18004 31006
rect 17948 30942 17950 30994
rect 18002 30942 18004 30994
rect 17836 30212 17892 30222
rect 17276 29922 17332 29932
rect 17724 30156 17836 30212
rect 17340 29820 17604 29830
rect 17396 29764 17444 29820
rect 17500 29764 17548 29820
rect 17340 29754 17604 29764
rect 17724 29426 17780 30156
rect 17836 30146 17892 30156
rect 17724 29374 17726 29426
rect 17778 29374 17780 29426
rect 17724 29362 17780 29374
rect 17388 29314 17444 29326
rect 17388 29262 17390 29314
rect 17442 29262 17444 29314
rect 17388 29092 17444 29262
rect 17836 29316 17892 29326
rect 17388 29026 17444 29036
rect 17500 29202 17556 29214
rect 17500 29150 17502 29202
rect 17554 29150 17556 29202
rect 17500 28420 17556 29150
rect 17500 28354 17556 28364
rect 17724 28980 17780 28990
rect 17340 28252 17604 28262
rect 17396 28196 17444 28252
rect 17500 28196 17548 28252
rect 17340 28186 17604 28196
rect 17276 28084 17332 28094
rect 17164 28028 17276 28084
rect 17276 28018 17332 28028
rect 17052 27794 17108 27804
rect 17724 27858 17780 28924
rect 17724 27806 17726 27858
rect 17778 27806 17780 27858
rect 17724 27794 17780 27806
rect 17052 27076 17108 27086
rect 16940 27020 17052 27076
rect 17052 27010 17108 27020
rect 17340 26684 17604 26694
rect 17396 26628 17444 26684
rect 17500 26628 17548 26684
rect 17340 26618 17604 26628
rect 16268 26516 16324 26526
rect 16156 26514 16324 26516
rect 16156 26462 16270 26514
rect 16322 26462 16324 26514
rect 16156 26460 16324 26462
rect 16268 26450 16324 26460
rect 17052 26516 17108 26526
rect 16156 26290 16212 26302
rect 16156 26238 16158 26290
rect 16210 26238 16212 26290
rect 16156 26180 16212 26238
rect 16828 26290 16884 26302
rect 16828 26238 16830 26290
rect 16882 26238 16884 26290
rect 16156 26114 16212 26124
rect 16604 26180 16660 26190
rect 16604 26086 16660 26124
rect 16380 26066 16436 26078
rect 16380 26014 16382 26066
rect 16434 26014 16436 26066
rect 16156 25956 16212 25966
rect 16212 25900 16324 25956
rect 16156 25890 16212 25900
rect 16044 25452 16212 25508
rect 16044 25284 16100 25294
rect 15484 24946 15652 24948
rect 15484 24894 15486 24946
rect 15538 24894 15652 24946
rect 15484 24892 15652 24894
rect 15708 25282 16100 25284
rect 15708 25230 16046 25282
rect 16098 25230 16100 25282
rect 15708 25228 16100 25230
rect 15484 24882 15540 24892
rect 15260 24546 15316 24556
rect 15372 24722 15428 24734
rect 15372 24670 15374 24722
rect 15426 24670 15428 24722
rect 15260 24276 15316 24286
rect 15260 23938 15316 24220
rect 15372 24052 15428 24670
rect 15596 24724 15652 24734
rect 15708 24724 15764 25228
rect 16044 25218 16100 25228
rect 15596 24722 15764 24724
rect 15596 24670 15598 24722
rect 15650 24670 15764 24722
rect 15596 24668 15764 24670
rect 15932 24724 15988 24734
rect 15596 24658 15652 24668
rect 15932 24630 15988 24668
rect 16156 24052 16212 25452
rect 16268 25506 16324 25900
rect 16268 25454 16270 25506
rect 16322 25454 16324 25506
rect 16268 25442 16324 25454
rect 16380 25508 16436 26014
rect 16828 25730 16884 26238
rect 16828 25678 16830 25730
rect 16882 25678 16884 25730
rect 16828 25666 16884 25678
rect 16940 25956 16996 25966
rect 16940 25618 16996 25900
rect 16940 25566 16942 25618
rect 16994 25566 16996 25618
rect 16940 25554 16996 25566
rect 16380 25442 16436 25452
rect 16492 25396 16548 25406
rect 16828 25396 16884 25406
rect 16492 25394 16660 25396
rect 16492 25342 16494 25394
rect 16546 25342 16660 25394
rect 16492 25340 16660 25342
rect 16492 25330 16548 25340
rect 16268 25172 16324 25182
rect 16324 25116 16548 25172
rect 16268 25106 16324 25116
rect 16492 24946 16548 25116
rect 16492 24894 16494 24946
rect 16546 24894 16548 24946
rect 16492 24882 16548 24894
rect 16268 24836 16324 24846
rect 16268 24742 16324 24780
rect 16604 24276 16660 25340
rect 16716 24836 16772 24846
rect 16716 24742 16772 24780
rect 16828 24834 16884 25340
rect 16828 24782 16830 24834
rect 16882 24782 16884 24834
rect 16828 24612 16884 24782
rect 16828 24546 16884 24556
rect 16604 24220 16772 24276
rect 15372 23986 15428 23996
rect 15932 23996 16212 24052
rect 16604 24052 16660 24062
rect 15596 23940 15652 23950
rect 15260 23886 15262 23938
rect 15314 23886 15316 23938
rect 15260 23874 15316 23886
rect 15484 23938 15652 23940
rect 15484 23886 15598 23938
rect 15650 23886 15652 23938
rect 15484 23884 15652 23886
rect 15148 22530 15204 22540
rect 15372 22596 15428 22606
rect 15484 22596 15540 23884
rect 15596 23874 15652 23884
rect 15708 23380 15764 23390
rect 15708 22820 15764 23324
rect 15820 22932 15876 22942
rect 15820 22838 15876 22876
rect 15708 22754 15764 22764
rect 15372 22594 15540 22596
rect 15372 22542 15374 22594
rect 15426 22542 15540 22594
rect 15372 22540 15540 22542
rect 15372 22530 15428 22540
rect 15036 21970 15092 21980
rect 15820 22146 15876 22158
rect 15820 22094 15822 22146
rect 15874 22094 15876 22146
rect 14364 21476 14420 21756
rect 14700 21756 14980 21812
rect 15820 21924 15876 22094
rect 14364 21420 14644 21476
rect 14252 20850 14308 20860
rect 14252 20692 14308 20702
rect 14252 20690 14420 20692
rect 14252 20638 14254 20690
rect 14306 20638 14420 20690
rect 14252 20636 14420 20638
rect 14252 20626 14308 20636
rect 14364 20242 14420 20636
rect 14364 20190 14366 20242
rect 14418 20190 14420 20242
rect 14140 20132 14308 20188
rect 14364 20178 14420 20190
rect 13916 20020 13972 20030
rect 14140 20020 14196 20030
rect 13916 20018 14196 20020
rect 13916 19966 13918 20018
rect 13970 19966 14142 20018
rect 14194 19966 14196 20018
rect 13916 19964 14196 19966
rect 13916 19954 13972 19964
rect 14140 19954 14196 19964
rect 14252 19796 14308 20132
rect 14476 20132 14532 20142
rect 14364 20020 14420 20030
rect 14364 19926 14420 19964
rect 14252 19740 14420 19796
rect 14140 19348 14196 19358
rect 14140 19234 14196 19292
rect 14140 19182 14142 19234
rect 14194 19182 14196 19234
rect 14140 19170 14196 19182
rect 13916 19010 13972 19022
rect 13916 18958 13918 19010
rect 13970 18958 13972 19010
rect 13916 18788 13972 18958
rect 13916 18722 13972 18732
rect 13804 18610 13860 18620
rect 13020 18510 13022 18562
rect 13074 18510 13076 18562
rect 13020 18498 13076 18510
rect 13356 18562 13412 18574
rect 13356 18510 13358 18562
rect 13410 18510 13412 18562
rect 13356 18452 13412 18510
rect 13468 18452 13524 18462
rect 13356 18450 13524 18452
rect 13356 18398 13470 18450
rect 13522 18398 13524 18450
rect 13356 18396 13524 18398
rect 13468 18386 13524 18396
rect 13916 18452 13972 18462
rect 13916 18358 13972 18396
rect 14028 18450 14084 18462
rect 14028 18398 14030 18450
rect 14082 18398 14084 18450
rect 13692 18338 13748 18350
rect 13692 18286 13694 18338
rect 13746 18286 13748 18338
rect 13308 18060 13572 18070
rect 13364 18004 13412 18060
rect 13468 18004 13516 18060
rect 13308 17994 13572 18004
rect 13692 18004 13748 18286
rect 14028 18228 14084 18398
rect 14028 18162 14084 18172
rect 13692 17948 14308 18004
rect 14252 17778 14308 17948
rect 14252 17726 14254 17778
rect 14306 17726 14308 17778
rect 14252 17714 14308 17726
rect 12908 17602 12964 17612
rect 13580 17668 13636 17678
rect 13580 17574 13636 17612
rect 14364 17556 14420 19740
rect 14476 18676 14532 20076
rect 14588 20018 14644 21420
rect 14588 19966 14590 20018
rect 14642 19966 14644 20018
rect 14588 19954 14644 19966
rect 14476 18610 14532 18620
rect 14476 18450 14532 18462
rect 14476 18398 14478 18450
rect 14530 18398 14532 18450
rect 14476 18228 14532 18398
rect 14476 18162 14532 18172
rect 14140 17500 14420 17556
rect 12348 17276 12516 17332
rect 12684 17442 12740 17454
rect 12684 17390 12686 17442
rect 12738 17390 12740 17442
rect 11788 17220 11844 17230
rect 11564 16884 11620 16894
rect 11564 16790 11620 16828
rect 11676 16100 11732 16110
rect 11788 16100 11844 17164
rect 12348 17106 12404 17276
rect 12684 17220 12740 17390
rect 12684 17154 12740 17164
rect 12348 17054 12350 17106
rect 12402 17054 12404 17106
rect 12348 17042 12404 17054
rect 12572 16996 12628 17006
rect 12460 16884 12516 16894
rect 11732 16044 11844 16100
rect 12348 16828 12460 16884
rect 11676 16006 11732 16044
rect 11340 15934 11342 15986
rect 11394 15934 11396 15986
rect 10556 15876 10612 15886
rect 10220 15874 10612 15876
rect 10220 15822 10558 15874
rect 10610 15822 10612 15874
rect 10220 15820 10612 15822
rect 9276 15708 9540 15718
rect 9332 15652 9380 15708
rect 9436 15652 9484 15708
rect 9276 15642 9540 15652
rect 8540 14466 8596 14476
rect 8652 15428 8708 15438
rect 8652 14530 8708 15372
rect 10220 15428 10276 15820
rect 10556 15810 10612 15820
rect 10444 15540 10500 15550
rect 10444 15538 11172 15540
rect 10444 15486 10446 15538
rect 10498 15486 11172 15538
rect 10444 15484 11172 15486
rect 10444 15474 10500 15484
rect 10220 15334 10276 15372
rect 10556 15316 10612 15326
rect 10556 15222 10612 15260
rect 10668 15314 10724 15326
rect 10668 15262 10670 15314
rect 10722 15262 10724 15314
rect 10556 14980 10612 14990
rect 8652 14478 8654 14530
rect 8706 14478 8708 14530
rect 8652 14466 8708 14478
rect 8988 14642 9044 14654
rect 8988 14590 8990 14642
rect 9042 14590 9044 14642
rect 8540 14308 8596 14318
rect 8988 14308 9044 14590
rect 8596 14252 9044 14308
rect 8540 14214 8596 14252
rect 8988 13972 9044 14252
rect 9276 14140 9540 14150
rect 9332 14084 9380 14140
rect 9436 14084 9484 14140
rect 9276 14074 9540 14084
rect 8988 13906 9044 13916
rect 10556 13970 10612 14924
rect 10556 13918 10558 13970
rect 10610 13918 10612 13970
rect 10556 13906 10612 13918
rect 10668 13970 10724 15262
rect 11116 14642 11172 15484
rect 11228 15316 11284 15326
rect 11228 15222 11284 15260
rect 11340 14980 11396 15934
rect 12348 15538 12404 16828
rect 12460 16818 12516 16828
rect 12348 15486 12350 15538
rect 12402 15486 12404 15538
rect 12348 15474 12404 15486
rect 11340 14914 11396 14924
rect 11452 15316 11508 15326
rect 11116 14590 11118 14642
rect 11170 14590 11172 14642
rect 11116 14578 11172 14590
rect 10668 13918 10670 13970
rect 10722 13918 10724 13970
rect 10668 13906 10724 13918
rect 10780 13972 10836 13982
rect 10780 13878 10836 13916
rect 11004 13858 11060 13870
rect 11004 13806 11006 13858
rect 11058 13806 11060 13858
rect 11004 13748 11060 13806
rect 10668 13692 11060 13748
rect 8988 13636 9044 13646
rect 8428 13634 9044 13636
rect 8428 13582 8990 13634
rect 9042 13582 9044 13634
rect 8428 13580 9044 13582
rect 8988 13570 9044 13580
rect 10220 13636 10276 13646
rect 10668 13636 10724 13692
rect 10220 13634 10724 13636
rect 10220 13582 10222 13634
rect 10274 13582 10724 13634
rect 10220 13580 10724 13582
rect 8540 12964 8596 12974
rect 9212 12964 9268 12974
rect 8540 12870 8596 12908
rect 9100 12908 9212 12964
rect 7756 12852 7812 12862
rect 7756 12758 7812 12796
rect 7532 12290 7588 12302
rect 7532 12238 7534 12290
rect 7586 12238 7588 12290
rect 7532 12068 7588 12238
rect 7532 12002 7588 12012
rect 7644 12178 7700 12190
rect 7644 12126 7646 12178
rect 7698 12126 7700 12178
rect 7644 11060 7700 12126
rect 8092 12068 8148 12078
rect 8092 11974 8148 12012
rect 8540 12066 8596 12078
rect 8540 12014 8542 12066
rect 8594 12014 8596 12066
rect 8540 11620 8596 12014
rect 8204 11564 8596 11620
rect 7644 10994 7700 11004
rect 7868 11508 7924 11518
rect 6860 10782 6862 10834
rect 6914 10782 6916 10834
rect 6860 10770 6916 10782
rect 7196 10892 7476 10948
rect 6748 10670 6750 10722
rect 6802 10670 6804 10722
rect 6748 10658 6804 10670
rect 6972 10610 7028 10622
rect 6972 10558 6974 10610
rect 7026 10558 7028 10610
rect 6412 9734 6468 9772
rect 6524 10386 6580 10398
rect 6524 10334 6526 10386
rect 6578 10334 6580 10386
rect 6188 9090 6244 9100
rect 5964 8932 6020 8942
rect 5852 8930 6244 8932
rect 5852 8878 5966 8930
rect 6018 8878 6244 8930
rect 5852 8876 6244 8878
rect 5964 8866 6020 8876
rect 5180 8754 5236 8764
rect 5244 8652 5508 8662
rect 5300 8596 5348 8652
rect 5404 8596 5452 8652
rect 5244 8586 5508 8596
rect 4620 8318 4622 8370
rect 4674 8318 4676 8370
rect 4620 5122 4676 8318
rect 5852 8428 6132 8484
rect 5852 8370 5908 8428
rect 5852 8318 5854 8370
rect 5906 8318 5908 8370
rect 5852 8306 5908 8318
rect 5964 8258 6020 8270
rect 5964 8206 5966 8258
rect 6018 8206 6020 8258
rect 5740 8148 5796 8158
rect 5740 8054 5796 8092
rect 5180 8034 5236 8046
rect 5180 7982 5182 8034
rect 5234 7982 5236 8034
rect 5180 7924 5236 7982
rect 5180 7858 5236 7868
rect 5516 7812 5572 7822
rect 4956 7700 5012 7710
rect 4956 7586 5012 7644
rect 4956 7534 4958 7586
rect 5010 7534 5012 7586
rect 4844 7474 4900 7486
rect 4844 7422 4846 7474
rect 4898 7422 4900 7474
rect 4844 7252 4900 7422
rect 4844 7186 4900 7196
rect 4844 6690 4900 6702
rect 4844 6638 4846 6690
rect 4898 6638 4900 6690
rect 4844 6580 4900 6638
rect 4844 6514 4900 6524
rect 4956 6468 5012 7534
rect 5404 7476 5460 7486
rect 5516 7476 5572 7756
rect 5852 7698 5908 7710
rect 5852 7646 5854 7698
rect 5906 7646 5908 7698
rect 5404 7474 5572 7476
rect 5404 7422 5406 7474
rect 5458 7422 5572 7474
rect 5404 7420 5572 7422
rect 5628 7476 5684 7486
rect 5628 7474 5796 7476
rect 5628 7422 5630 7474
rect 5682 7422 5796 7474
rect 5628 7420 5796 7422
rect 5404 7410 5460 7420
rect 5628 7410 5684 7420
rect 5180 7364 5236 7374
rect 5068 7362 5236 7364
rect 5068 7310 5182 7362
rect 5234 7310 5236 7362
rect 5068 7308 5236 7310
rect 5068 6692 5124 7308
rect 5180 7298 5236 7308
rect 5740 7252 5796 7420
rect 5628 7196 5796 7252
rect 5244 7084 5508 7094
rect 5300 7028 5348 7084
rect 5404 7028 5452 7084
rect 5244 7018 5508 7028
rect 5516 6804 5572 6814
rect 5068 6636 5236 6692
rect 5068 6468 5124 6478
rect 4956 6466 5124 6468
rect 4956 6414 5070 6466
rect 5122 6414 5124 6466
rect 4956 6412 5124 6414
rect 4956 5796 5012 6412
rect 5068 6402 5124 6412
rect 5180 6132 5236 6636
rect 5180 6066 5236 6076
rect 5292 6244 5348 6254
rect 5292 6130 5348 6188
rect 5292 6078 5294 6130
rect 5346 6078 5348 6130
rect 5292 6066 5348 6078
rect 5068 6020 5124 6030
rect 5068 5926 5124 5964
rect 5404 5906 5460 5918
rect 5404 5854 5406 5906
rect 5458 5854 5460 5906
rect 5404 5796 5460 5854
rect 5516 5906 5572 6748
rect 5516 5854 5518 5906
rect 5570 5854 5572 5906
rect 5516 5842 5572 5854
rect 4956 5740 5460 5796
rect 5244 5516 5508 5526
rect 5300 5460 5348 5516
rect 5404 5460 5452 5516
rect 5244 5450 5508 5460
rect 5628 5348 5684 7196
rect 5852 6916 5908 7646
rect 5964 7700 6020 8206
rect 6076 7700 6132 8428
rect 6188 8372 6244 8876
rect 6188 8306 6244 8316
rect 6300 8146 6356 8158
rect 6300 8094 6302 8146
rect 6354 8094 6356 8146
rect 6076 7644 6244 7700
rect 5964 7586 6020 7644
rect 5964 7534 5966 7586
rect 6018 7534 6020 7586
rect 5964 7522 6020 7534
rect 6076 7476 6132 7486
rect 6076 7382 6132 7420
rect 5740 6860 5908 6916
rect 5964 7364 6020 7374
rect 5740 6468 5796 6860
rect 5852 6692 5908 6702
rect 5852 6598 5908 6636
rect 5740 6402 5796 6412
rect 5628 5282 5684 5292
rect 5740 6132 5796 6142
rect 4620 5070 4622 5122
rect 4674 5070 4676 5122
rect 4620 5058 4676 5070
rect 5740 4450 5796 6076
rect 5964 5796 6020 7308
rect 6188 7140 6244 7644
rect 6300 7588 6356 8094
rect 6300 7522 6356 7532
rect 6188 7084 6356 7140
rect 5964 5794 6244 5796
rect 5964 5742 5966 5794
rect 6018 5742 6244 5794
rect 5964 5740 6244 5742
rect 5964 5730 6020 5740
rect 5964 5236 6020 5246
rect 5852 5180 5964 5236
rect 5852 5122 5908 5180
rect 5964 5170 6020 5180
rect 5852 5070 5854 5122
rect 5906 5070 5908 5122
rect 5852 5058 5908 5070
rect 6076 5124 6132 5134
rect 5740 4398 5742 4450
rect 5794 4398 5796 4450
rect 5740 4386 5796 4398
rect 4956 4340 5012 4350
rect 4508 4338 5012 4340
rect 4508 4286 4510 4338
rect 4562 4286 4958 4338
rect 5010 4286 5012 4338
rect 4508 4284 5012 4286
rect 4508 4274 4564 4284
rect 4956 4274 5012 4284
rect 5244 3948 5508 3958
rect 5300 3892 5348 3948
rect 5404 3892 5452 3948
rect 5244 3882 5508 3892
rect 6076 3668 6132 5068
rect 3276 3490 3332 3500
rect 5628 3612 6132 3668
rect 3164 3266 3220 3276
rect 4060 3442 4116 3454
rect 4060 3390 4062 3442
rect 4114 3390 4116 3442
rect 4060 800 4116 3390
rect 5516 3332 5572 3342
rect 5516 3238 5572 3276
rect 5628 800 5684 3612
rect 6188 3556 6244 5740
rect 6300 5684 6356 7084
rect 6524 6916 6580 10334
rect 6748 9716 6804 9726
rect 6972 9716 7028 10558
rect 7196 10052 7252 10892
rect 7756 10836 7812 10846
rect 7308 10834 7812 10836
rect 7308 10782 7758 10834
rect 7810 10782 7812 10834
rect 7308 10780 7812 10782
rect 7308 10722 7364 10780
rect 7756 10770 7812 10780
rect 7868 10834 7924 11452
rect 7868 10782 7870 10834
rect 7922 10782 7924 10834
rect 7868 10770 7924 10782
rect 8204 10836 8260 11564
rect 8652 11508 8708 11518
rect 8540 11452 8652 11508
rect 8428 11396 8484 11406
rect 7308 10670 7310 10722
rect 7362 10670 7364 10722
rect 7308 10658 7364 10670
rect 7644 10612 7700 10622
rect 7196 9986 7252 9996
rect 7532 10610 7700 10612
rect 7532 10558 7646 10610
rect 7698 10558 7700 10610
rect 7532 10556 7700 10558
rect 7084 9828 7140 9838
rect 7084 9734 7140 9772
rect 6804 9660 7028 9716
rect 7420 9716 7476 9726
rect 6748 9622 6804 9660
rect 7420 9622 7476 9660
rect 7308 9602 7364 9614
rect 7308 9550 7310 9602
rect 7362 9550 7364 9602
rect 7308 9380 7364 9550
rect 7308 9314 7364 9324
rect 7532 9604 7588 10556
rect 7644 10546 7700 10556
rect 8204 10610 8260 10780
rect 8204 10558 8206 10610
rect 8258 10558 8260 10610
rect 6748 8036 6804 8046
rect 6748 7476 6804 7980
rect 6748 7382 6804 7420
rect 6972 7474 7028 7486
rect 6972 7422 6974 7474
rect 7026 7422 7028 7474
rect 6300 5618 6356 5628
rect 6412 6692 6468 6702
rect 6412 5236 6468 6636
rect 6412 5170 6468 5180
rect 5740 3554 6244 3556
rect 5740 3502 6190 3554
rect 6242 3502 6244 3554
rect 5740 3500 6244 3502
rect 5740 3442 5796 3500
rect 6188 3490 6244 3500
rect 6524 5012 6580 6860
rect 6860 7362 6916 7374
rect 6860 7310 6862 7362
rect 6914 7310 6916 7362
rect 6860 6804 6916 7310
rect 6972 7364 7028 7422
rect 6972 7298 7028 7308
rect 7420 7474 7476 7486
rect 7420 7422 7422 7474
rect 7474 7422 7476 7474
rect 6860 6738 6916 6748
rect 7420 7028 7476 7422
rect 7532 7476 7588 9548
rect 7644 9714 7700 9726
rect 7644 9662 7646 9714
rect 7698 9662 7700 9714
rect 7644 7700 7700 9662
rect 7980 9604 8036 9614
rect 7980 9510 8036 9548
rect 7756 9380 7812 9390
rect 7812 9324 8148 9380
rect 7756 9314 7812 9324
rect 8092 9154 8148 9324
rect 8092 9102 8094 9154
rect 8146 9102 8148 9154
rect 8092 9090 8148 9102
rect 7868 8372 7924 8382
rect 7756 7700 7812 7710
rect 7644 7698 7812 7700
rect 7644 7646 7758 7698
rect 7810 7646 7812 7698
rect 7644 7644 7812 7646
rect 7756 7634 7812 7644
rect 7868 7698 7924 8316
rect 7868 7646 7870 7698
rect 7922 7646 7924 7698
rect 7868 7634 7924 7646
rect 7644 7476 7700 7486
rect 7532 7474 7700 7476
rect 7532 7422 7646 7474
rect 7698 7422 7700 7474
rect 7532 7420 7700 7422
rect 7644 7410 7700 7420
rect 8204 7474 8260 10558
rect 8316 11060 8372 11070
rect 8316 9716 8372 11004
rect 8316 9622 8372 9660
rect 8428 9380 8484 11340
rect 8540 9492 8596 11452
rect 8652 11442 8708 11452
rect 8988 11508 9044 11518
rect 8988 11414 9044 11452
rect 8652 10836 8708 10846
rect 8652 10742 8708 10780
rect 8764 10050 8820 10062
rect 8764 9998 8766 10050
rect 8818 9998 8820 10050
rect 8764 9828 8820 9998
rect 9100 9828 9156 12908
rect 9212 12898 9268 12908
rect 9996 12964 10052 12974
rect 9996 12870 10052 12908
rect 9276 12572 9540 12582
rect 9332 12516 9380 12572
rect 9436 12516 9484 12572
rect 9276 12506 9540 12516
rect 9436 11508 9492 11518
rect 9436 11414 9492 11452
rect 10220 11396 10276 13580
rect 10780 13524 10836 13534
rect 10780 13074 10836 13468
rect 10780 13022 10782 13074
rect 10834 13022 10836 13074
rect 10780 13010 10836 13022
rect 11452 12404 11508 15260
rect 12012 15204 12068 15214
rect 12236 15204 12292 15214
rect 12572 15204 12628 16940
rect 13132 16884 13188 16894
rect 13132 15316 13188 16828
rect 13916 16884 13972 16894
rect 13916 16790 13972 16828
rect 13308 16492 13572 16502
rect 13364 16436 13412 16492
rect 13468 16436 13516 16492
rect 13308 16426 13572 16436
rect 13356 15428 13412 15438
rect 13356 15334 13412 15372
rect 14028 15428 14084 15438
rect 14140 15428 14196 17500
rect 14700 17444 14756 21756
rect 14812 21588 14868 21598
rect 14812 20468 14868 21532
rect 15484 21474 15540 21486
rect 15484 21422 15486 21474
rect 15538 21422 15540 21474
rect 15484 21364 15540 21422
rect 15484 21298 15540 21308
rect 14812 20402 14868 20412
rect 15260 20244 15316 20254
rect 15260 20150 15316 20188
rect 15820 20132 15876 21868
rect 15932 21812 15988 23996
rect 16268 23940 16324 23950
rect 16156 23828 16212 23838
rect 16156 23734 16212 23772
rect 16044 23714 16100 23726
rect 16044 23662 16046 23714
rect 16098 23662 16100 23714
rect 16044 22036 16100 23662
rect 16268 23604 16324 23884
rect 16604 23826 16660 23996
rect 16604 23774 16606 23826
rect 16658 23774 16660 23826
rect 16604 23762 16660 23774
rect 16156 23548 16324 23604
rect 16380 23716 16436 23726
rect 16156 23380 16212 23548
rect 16156 22370 16212 23324
rect 16380 23268 16436 23660
rect 16380 23202 16436 23212
rect 16716 23268 16772 24220
rect 17052 24164 17108 26460
rect 17724 26516 17780 26526
rect 17724 26422 17780 26460
rect 17388 26404 17444 26414
rect 17388 25508 17444 26348
rect 17836 26178 17892 29260
rect 17948 28756 18004 30942
rect 18620 30996 18676 31006
rect 18620 30322 18676 30940
rect 18620 30270 18622 30322
rect 18674 30270 18676 30322
rect 18508 30212 18564 30222
rect 18396 29652 18452 29662
rect 18396 29558 18452 29596
rect 18172 29426 18228 29438
rect 18172 29374 18174 29426
rect 18226 29374 18228 29426
rect 18172 28980 18228 29374
rect 18284 29314 18340 29326
rect 18284 29262 18286 29314
rect 18338 29262 18340 29314
rect 18284 29204 18340 29262
rect 18284 29138 18340 29148
rect 18508 29092 18564 30156
rect 18620 29540 18676 30270
rect 19068 30212 19124 30222
rect 18956 30210 19124 30212
rect 18956 30158 19070 30210
rect 19122 30158 19124 30210
rect 18956 30156 19124 30158
rect 18620 29474 18676 29484
rect 18732 30100 18788 30110
rect 18508 29036 18676 29092
rect 18172 28924 18564 28980
rect 17948 28690 18004 28700
rect 18284 28756 18340 28766
rect 18284 28662 18340 28700
rect 18396 28644 18452 28654
rect 18396 28532 18452 28588
rect 18284 28476 18452 28532
rect 18172 26962 18228 26974
rect 18172 26910 18174 26962
rect 18226 26910 18228 26962
rect 18172 26908 18228 26910
rect 18060 26852 18228 26908
rect 18060 26292 18116 26852
rect 18284 26516 18340 28476
rect 18508 28308 18564 28924
rect 18620 28644 18676 29036
rect 18732 28866 18788 30044
rect 18844 29428 18900 29438
rect 18844 29334 18900 29372
rect 18732 28814 18734 28866
rect 18786 28814 18788 28866
rect 18732 28802 18788 28814
rect 18620 28588 18788 28644
rect 18732 28530 18788 28588
rect 18732 28478 18734 28530
rect 18786 28478 18788 28530
rect 18732 28466 18788 28478
rect 18844 28532 18900 28542
rect 18844 28438 18900 28476
rect 18508 28242 18564 28252
rect 18620 28420 18676 28430
rect 18508 28084 18564 28094
rect 18508 27990 18564 28028
rect 18396 26962 18452 26974
rect 18396 26910 18398 26962
rect 18450 26910 18452 26962
rect 18396 26852 18452 26910
rect 18396 26796 18564 26852
rect 18396 26516 18452 26526
rect 18284 26514 18452 26516
rect 18284 26462 18398 26514
rect 18450 26462 18452 26514
rect 18284 26460 18452 26462
rect 18396 26450 18452 26460
rect 18508 26404 18564 26796
rect 18620 26514 18676 28364
rect 18956 28308 19012 30156
rect 19068 30146 19124 30156
rect 19628 30210 19684 31500
rect 20860 31332 20916 32060
rect 21756 31444 21812 34200
rect 20748 30996 20804 31006
rect 20748 30902 20804 30940
rect 20412 30436 20468 30446
rect 19628 30158 19630 30210
rect 19682 30158 19684 30210
rect 19628 30146 19684 30158
rect 20076 30324 20132 30334
rect 20076 30212 20132 30268
rect 20300 30212 20356 30222
rect 20076 30156 20244 30212
rect 20076 29988 20132 29998
rect 19516 29316 19572 29326
rect 19516 29222 19572 29260
rect 20076 29092 20132 29932
rect 20188 29876 20244 30156
rect 20300 30098 20356 30156
rect 20300 30046 20302 30098
rect 20354 30046 20356 30098
rect 20300 30034 20356 30046
rect 20412 30098 20468 30380
rect 20636 30324 20692 30334
rect 20636 30230 20692 30268
rect 20412 30046 20414 30098
rect 20466 30046 20468 30098
rect 20412 30034 20468 30046
rect 20524 29986 20580 29998
rect 20524 29934 20526 29986
rect 20578 29934 20580 29986
rect 20524 29876 20580 29934
rect 20188 29820 20580 29876
rect 20524 29316 20580 29820
rect 20524 29250 20580 29260
rect 20748 29986 20804 29998
rect 20748 29934 20750 29986
rect 20802 29934 20804 29986
rect 19964 28756 20020 28766
rect 19292 28644 19348 28654
rect 19628 28644 19684 28654
rect 19292 28550 19348 28588
rect 19516 28588 19628 28644
rect 18844 28252 19012 28308
rect 19180 28418 19236 28430
rect 19180 28366 19182 28418
rect 19234 28366 19236 28418
rect 18732 27300 18788 27338
rect 18732 27234 18788 27244
rect 18620 26462 18622 26514
rect 18674 26462 18676 26514
rect 18620 26450 18676 26462
rect 18732 27074 18788 27086
rect 18732 27022 18734 27074
rect 18786 27022 18788 27074
rect 18732 26516 18788 27022
rect 18844 26628 18900 28252
rect 18956 27748 19012 27758
rect 18956 26850 19012 27692
rect 19180 27636 19236 28366
rect 19404 28420 19460 28430
rect 19404 27636 19460 28364
rect 19516 27748 19572 28588
rect 19628 28578 19684 28588
rect 19964 28642 20020 28700
rect 19964 28590 19966 28642
rect 20018 28590 20020 28642
rect 19964 28578 20020 28590
rect 19628 28420 19684 28430
rect 19628 28418 19796 28420
rect 19628 28366 19630 28418
rect 19682 28366 19796 28418
rect 19628 28364 19796 28366
rect 19628 28354 19684 28364
rect 19516 27692 19684 27748
rect 19404 27580 19572 27636
rect 19180 26908 19236 27580
rect 19292 27076 19348 27086
rect 19292 26982 19348 27020
rect 18956 26798 18958 26850
rect 19010 26798 19012 26850
rect 18956 26786 19012 26798
rect 19068 26852 19236 26908
rect 18844 26562 18900 26572
rect 18732 26450 18788 26460
rect 18508 26338 18564 26348
rect 17836 26126 17838 26178
rect 17890 26126 17892 26178
rect 17836 26114 17892 26126
rect 17948 26236 18116 26292
rect 18172 26292 18228 26302
rect 17500 26068 17556 26078
rect 17500 25974 17556 26012
rect 17724 25620 17780 25630
rect 17724 25526 17780 25564
rect 17500 25508 17556 25518
rect 17388 25506 17556 25508
rect 17388 25454 17502 25506
rect 17554 25454 17556 25506
rect 17388 25452 17556 25454
rect 17500 25442 17556 25452
rect 17836 25508 17892 25518
rect 17276 25396 17332 25406
rect 17052 24098 17108 24108
rect 17164 25394 17332 25396
rect 17164 25342 17278 25394
rect 17330 25342 17332 25394
rect 17164 25340 17332 25342
rect 16716 23202 16772 23212
rect 16940 24052 16996 24062
rect 16940 23714 16996 23996
rect 16940 23662 16942 23714
rect 16994 23662 16996 23714
rect 16716 23042 16772 23054
rect 16716 22990 16718 23042
rect 16770 22990 16772 23042
rect 16268 22932 16324 22942
rect 16268 22930 16436 22932
rect 16268 22878 16270 22930
rect 16322 22878 16436 22930
rect 16268 22876 16436 22878
rect 16268 22866 16324 22876
rect 16380 22484 16436 22876
rect 16492 22930 16548 22942
rect 16492 22878 16494 22930
rect 16546 22878 16548 22930
rect 16492 22708 16548 22878
rect 16604 22932 16660 22942
rect 16716 22932 16772 22990
rect 16828 22932 16884 22942
rect 16716 22876 16828 22932
rect 16604 22708 16660 22876
rect 16828 22866 16884 22876
rect 16604 22652 16772 22708
rect 16492 22642 16548 22652
rect 16380 22418 16436 22428
rect 16156 22318 16158 22370
rect 16210 22318 16212 22370
rect 16156 22306 16212 22318
rect 16268 22372 16324 22382
rect 16268 22278 16324 22316
rect 16716 22370 16772 22652
rect 16716 22318 16718 22370
rect 16770 22318 16772 22370
rect 16716 22306 16772 22318
rect 16044 21970 16100 21980
rect 16380 22146 16436 22158
rect 16380 22094 16382 22146
rect 16434 22094 16436 22146
rect 16044 21812 16100 21822
rect 15932 21810 16100 21812
rect 15932 21758 16046 21810
rect 16098 21758 16100 21810
rect 15932 21756 16100 21758
rect 16044 21746 16100 21756
rect 16380 20916 16436 22094
rect 16716 22148 16772 22158
rect 16940 22148 16996 23662
rect 17052 23940 17108 23950
rect 17052 22372 17108 23884
rect 17164 23716 17220 25340
rect 17276 25330 17332 25340
rect 17836 25284 17892 25452
rect 17724 25228 17892 25284
rect 17340 25116 17604 25126
rect 17396 25060 17444 25116
rect 17500 25060 17548 25116
rect 17340 25050 17604 25060
rect 17388 24948 17444 24958
rect 17388 24834 17444 24892
rect 17388 24782 17390 24834
rect 17442 24782 17444 24834
rect 17388 24770 17444 24782
rect 17500 24836 17556 24846
rect 17500 24834 17668 24836
rect 17500 24782 17502 24834
rect 17554 24782 17668 24834
rect 17500 24780 17668 24782
rect 17500 24770 17556 24780
rect 17500 24612 17556 24622
rect 17500 24498 17556 24556
rect 17500 24446 17502 24498
rect 17554 24446 17556 24498
rect 17500 24434 17556 24446
rect 17612 24500 17668 24780
rect 17500 24276 17556 24286
rect 17612 24276 17668 24444
rect 17556 24220 17668 24276
rect 17500 24210 17556 24220
rect 17164 23650 17220 23660
rect 17612 23716 17668 23754
rect 17612 23650 17668 23660
rect 17340 23548 17604 23558
rect 17396 23492 17444 23548
rect 17500 23492 17548 23548
rect 17340 23482 17604 23492
rect 17500 23044 17556 23054
rect 17724 23044 17780 25228
rect 17948 23828 18004 26236
rect 18172 26198 18228 26236
rect 18732 26292 18788 26302
rect 18620 26180 18676 26190
rect 18060 26068 18116 26078
rect 18060 25282 18116 26012
rect 18060 25230 18062 25282
rect 18114 25230 18116 25282
rect 18060 25218 18116 25230
rect 18172 25564 18564 25620
rect 18172 24948 18228 25564
rect 18508 25508 18564 25564
rect 18508 25414 18564 25452
rect 17948 23762 18004 23772
rect 18060 24892 18228 24948
rect 18284 25396 18340 25406
rect 17500 23042 17780 23044
rect 17500 22990 17502 23042
rect 17554 22990 17780 23042
rect 17500 22988 17780 22990
rect 17836 23714 17892 23726
rect 17836 23662 17838 23714
rect 17890 23662 17892 23714
rect 17836 23604 17892 23662
rect 17500 22820 17556 22988
rect 17500 22754 17556 22764
rect 17836 22708 17892 23548
rect 17836 22642 17892 22652
rect 18060 23716 18116 24892
rect 18284 24834 18340 25340
rect 18508 25060 18564 25070
rect 18396 24948 18452 24958
rect 18396 24854 18452 24892
rect 18284 24782 18286 24834
rect 18338 24782 18340 24834
rect 18284 24770 18340 24782
rect 18172 24724 18228 24734
rect 18172 23938 18228 24668
rect 18172 23886 18174 23938
rect 18226 23886 18228 23938
rect 18172 23874 18228 23886
rect 18508 24388 18564 25004
rect 18508 23938 18564 24332
rect 18508 23886 18510 23938
rect 18562 23886 18564 23938
rect 18508 23874 18564 23886
rect 18060 22594 18116 23660
rect 18620 23492 18676 26124
rect 18732 26178 18788 26236
rect 18844 26292 18900 26302
rect 19068 26292 19124 26852
rect 19404 26850 19460 26862
rect 19404 26798 19406 26850
rect 19458 26798 19460 26850
rect 19292 26404 19348 26414
rect 18844 26290 19124 26292
rect 18844 26238 18846 26290
rect 18898 26238 19124 26290
rect 18844 26236 19124 26238
rect 19180 26290 19236 26302
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 18844 26226 18900 26236
rect 18732 26126 18734 26178
rect 18786 26126 18788 26178
rect 18732 26114 18788 26126
rect 19180 26180 19236 26238
rect 19180 26114 19236 26124
rect 19292 25844 19348 26348
rect 18844 25788 19348 25844
rect 18844 25506 18900 25788
rect 18956 25620 19012 25630
rect 18956 25526 19012 25564
rect 18844 25454 18846 25506
rect 18898 25454 18900 25506
rect 18844 25442 18900 25454
rect 18844 25284 18900 25294
rect 18844 25172 18900 25228
rect 18732 25116 18900 25172
rect 19068 25172 19124 25788
rect 19180 25506 19236 25518
rect 19180 25454 19182 25506
rect 19234 25454 19236 25506
rect 19180 25284 19236 25454
rect 19404 25284 19460 26798
rect 19516 26290 19572 27580
rect 19628 26404 19684 27692
rect 19740 26908 19796 28364
rect 19964 27076 20020 27086
rect 20076 27076 20132 29036
rect 20412 28756 20468 28766
rect 20300 28644 20356 28654
rect 20300 28550 20356 28588
rect 20188 28418 20244 28430
rect 20412 28420 20468 28700
rect 20636 28532 20692 28542
rect 20636 28438 20692 28476
rect 20188 28366 20190 28418
rect 20242 28366 20244 28418
rect 20188 27300 20244 28366
rect 20188 27234 20244 27244
rect 20300 28364 20468 28420
rect 19964 27074 20132 27076
rect 19964 27022 19966 27074
rect 20018 27022 20132 27074
rect 19964 27020 20132 27022
rect 19964 27010 20020 27020
rect 20300 26908 20356 28364
rect 20524 28084 20580 28094
rect 20580 28028 20692 28084
rect 20524 27990 20580 28028
rect 20412 27860 20468 27870
rect 20412 27766 20468 27804
rect 20524 27636 20580 27646
rect 20524 27542 20580 27580
rect 20524 27076 20580 27114
rect 20524 27010 20580 27020
rect 20412 26964 20468 26984
rect 20636 26962 20692 28028
rect 20636 26910 20638 26962
rect 20690 26910 20692 26962
rect 19740 26852 19908 26908
rect 20300 26852 20580 26908
rect 20636 26898 20692 26910
rect 20748 26908 20804 29934
rect 20860 28868 20916 31276
rect 21196 31388 21812 31444
rect 20972 31108 21028 31118
rect 21028 31052 21140 31108
rect 20972 31042 21028 31052
rect 20860 28802 20916 28812
rect 20972 29428 21028 29438
rect 20860 28532 20916 28542
rect 20860 27860 20916 28476
rect 20860 27076 20916 27804
rect 20972 27860 21028 29372
rect 21084 28532 21140 31052
rect 21084 28466 21140 28476
rect 21196 28420 21252 31388
rect 21756 31220 21812 31230
rect 21756 31126 21812 31164
rect 22876 31220 22932 34200
rect 22876 31154 22932 31164
rect 23884 33460 23940 33470
rect 23884 31668 23940 33404
rect 23660 31108 23716 31118
rect 23660 31014 23716 31052
rect 23884 30994 23940 31612
rect 23884 30942 23886 30994
rect 23938 30942 23940 30994
rect 23884 30930 23940 30942
rect 21868 30772 21924 30782
rect 21372 30604 21636 30614
rect 21428 30548 21476 30604
rect 21532 30548 21580 30604
rect 21372 30538 21636 30548
rect 21308 30210 21364 30222
rect 21308 30158 21310 30210
rect 21362 30158 21364 30210
rect 21308 29428 21364 30158
rect 21308 29362 21364 29372
rect 21756 29314 21812 29326
rect 21756 29262 21758 29314
rect 21810 29262 21812 29314
rect 21372 29036 21636 29046
rect 21428 28980 21476 29036
rect 21532 28980 21580 29036
rect 21372 28970 21636 28980
rect 21308 28868 21364 28878
rect 21308 28532 21364 28812
rect 21644 28756 21700 28766
rect 21756 28756 21812 29262
rect 21700 28700 21812 28756
rect 21868 28754 21924 30716
rect 23436 30436 23492 30446
rect 23436 30212 23492 30380
rect 21868 28702 21870 28754
rect 21922 28702 21924 28754
rect 21644 28690 21700 28700
rect 21868 28690 21924 28702
rect 22092 30098 22148 30110
rect 22092 30046 22094 30098
rect 22146 30046 22148 30098
rect 21308 28476 21476 28532
rect 21420 28420 21476 28476
rect 21532 28530 21588 28542
rect 21532 28478 21534 28530
rect 21586 28478 21588 28530
rect 21532 28420 21588 28478
rect 21420 28364 21588 28420
rect 21644 28532 21700 28542
rect 21644 28420 21700 28476
rect 21868 28532 21924 28542
rect 21868 28438 21924 28476
rect 21756 28420 21812 28430
rect 21644 28418 21812 28420
rect 21644 28366 21758 28418
rect 21810 28366 21812 28418
rect 21644 28364 21812 28366
rect 21196 28354 21252 28364
rect 21756 28308 21812 28364
rect 21756 28252 21924 28308
rect 20972 27858 21252 27860
rect 20972 27806 20974 27858
rect 21026 27806 21252 27858
rect 20972 27804 21252 27806
rect 20972 27794 21028 27804
rect 21196 27300 21252 27804
rect 21756 27748 21812 27758
rect 21756 27654 21812 27692
rect 21372 27468 21636 27478
rect 21428 27412 21476 27468
rect 21532 27412 21580 27468
rect 21372 27402 21636 27412
rect 21196 27244 21812 27300
rect 20860 27010 20916 27020
rect 21308 26962 21364 26974
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 20748 26852 20916 26908
rect 19628 26338 19684 26348
rect 19740 26516 19796 26526
rect 19516 26238 19518 26290
rect 19570 26238 19572 26290
rect 19516 26226 19572 26238
rect 19740 26290 19796 26460
rect 19740 26238 19742 26290
rect 19794 26238 19796 26290
rect 19628 26180 19684 26190
rect 19628 26086 19684 26124
rect 19740 25508 19796 26238
rect 19740 25442 19796 25452
rect 19180 25218 19236 25228
rect 19292 25282 19460 25284
rect 19292 25230 19406 25282
rect 19458 25230 19460 25282
rect 19292 25228 19460 25230
rect 18732 24834 18788 25116
rect 19068 25106 19124 25116
rect 18844 24948 18900 24958
rect 18844 24946 19236 24948
rect 18844 24894 18846 24946
rect 18898 24894 19236 24946
rect 18844 24892 19236 24894
rect 18844 24882 18900 24892
rect 18732 24782 18734 24834
rect 18786 24782 18788 24834
rect 18732 24724 18788 24782
rect 18732 24668 19012 24724
rect 18844 24498 18900 24510
rect 18844 24446 18846 24498
rect 18898 24446 18900 24498
rect 18732 23940 18788 23950
rect 18732 23846 18788 23884
rect 18508 23380 18564 23390
rect 18508 23266 18564 23324
rect 18508 23214 18510 23266
rect 18562 23214 18564 23266
rect 18508 23202 18564 23214
rect 18060 22542 18062 22594
rect 18114 22542 18116 22594
rect 18060 22530 18116 22542
rect 18284 23154 18340 23166
rect 18284 23102 18286 23154
rect 18338 23102 18340 23154
rect 17388 22372 17444 22382
rect 17052 22316 17220 22372
rect 17052 22148 17108 22158
rect 16940 22146 17108 22148
rect 16940 22094 17054 22146
rect 17106 22094 17108 22146
rect 16940 22092 17108 22094
rect 16492 21810 16548 21822
rect 16492 21758 16494 21810
rect 16546 21758 16548 21810
rect 16492 21700 16548 21758
rect 16492 21634 16548 21644
rect 16268 20914 16436 20916
rect 16268 20862 16382 20914
rect 16434 20862 16436 20914
rect 16268 20860 16436 20862
rect 16156 20244 16212 20254
rect 16268 20244 16324 20860
rect 16380 20850 16436 20860
rect 16604 20804 16660 20814
rect 16212 20188 16324 20244
rect 16492 20748 16604 20804
rect 16156 20150 16212 20188
rect 15820 20066 15876 20076
rect 15036 20020 15092 20030
rect 15036 19926 15092 19964
rect 15372 20018 15428 20030
rect 15372 19966 15374 20018
rect 15426 19966 15428 20018
rect 15036 19572 15092 19582
rect 15036 19236 15092 19516
rect 15372 19348 15428 19966
rect 16044 20018 16100 20030
rect 16044 19966 16046 20018
rect 16098 19966 16100 20018
rect 15372 19292 15652 19348
rect 15036 19180 15204 19236
rect 14924 19122 14980 19134
rect 14924 19070 14926 19122
rect 14978 19070 14980 19122
rect 14924 18674 14980 19070
rect 14924 18622 14926 18674
rect 14978 18622 14980 18674
rect 14924 18610 14980 18622
rect 15036 18788 15092 18798
rect 15036 18562 15092 18732
rect 15036 18510 15038 18562
rect 15090 18510 15092 18562
rect 15036 18498 15092 18510
rect 14812 18452 14868 18462
rect 14812 18358 14868 18396
rect 15148 18340 15204 19180
rect 15484 18676 15540 18686
rect 15484 18582 15540 18620
rect 15596 18564 15652 19292
rect 16044 18900 16100 19966
rect 16380 20020 16436 20030
rect 16492 20020 16548 20748
rect 16604 20738 16660 20748
rect 16380 20018 16548 20020
rect 16380 19966 16382 20018
rect 16434 19966 16548 20018
rect 16380 19964 16548 19966
rect 16380 19954 16436 19964
rect 15596 18470 15652 18508
rect 15932 18844 16100 18900
rect 16156 19124 16212 19134
rect 15260 18452 15316 18462
rect 15260 18358 15316 18396
rect 15820 18452 15876 18462
rect 15820 18358 15876 18396
rect 14252 17388 14756 17444
rect 15036 18284 15204 18340
rect 14252 17106 14308 17388
rect 14252 17054 14254 17106
rect 14306 17054 14308 17106
rect 14252 17042 14308 17054
rect 15036 16324 15092 18284
rect 15932 17780 15988 18844
rect 16044 18562 16100 18574
rect 16044 18510 16046 18562
rect 16098 18510 16100 18562
rect 16044 18452 16100 18510
rect 16156 18564 16212 19068
rect 16156 18470 16212 18508
rect 16044 18340 16100 18396
rect 16044 18284 16436 18340
rect 15932 17714 15988 17724
rect 16380 17778 16436 18284
rect 16380 17726 16382 17778
rect 16434 17726 16436 17778
rect 16380 17714 16436 17726
rect 16716 17556 16772 22092
rect 17052 22082 17108 22092
rect 16940 21476 16996 21486
rect 16940 21474 17108 21476
rect 16940 21422 16942 21474
rect 16994 21422 17108 21474
rect 16940 21420 17108 21422
rect 16940 21410 16996 21420
rect 16940 20916 16996 20926
rect 16828 20578 16884 20590
rect 16828 20526 16830 20578
rect 16882 20526 16884 20578
rect 16828 19236 16884 20526
rect 16940 20242 16996 20860
rect 16940 20190 16942 20242
rect 16994 20190 16996 20242
rect 16940 20178 16996 20190
rect 17052 19572 17108 21420
rect 17052 19506 17108 19516
rect 16828 17778 16884 19180
rect 17052 19348 17108 19358
rect 17164 19348 17220 22316
rect 17388 22258 17444 22316
rect 17388 22206 17390 22258
rect 17442 22206 17444 22258
rect 17388 22194 17444 22206
rect 17948 22260 18004 22270
rect 17340 21980 17604 21990
rect 17396 21924 17444 21980
rect 17500 21924 17548 21980
rect 17340 21914 17604 21924
rect 17612 21474 17668 21486
rect 17612 21422 17614 21474
rect 17666 21422 17668 21474
rect 17388 21364 17444 21374
rect 17388 20914 17444 21308
rect 17612 21252 17668 21422
rect 17948 21474 18004 22204
rect 17948 21422 17950 21474
rect 18002 21422 18004 21474
rect 17948 21410 18004 21422
rect 18172 22146 18228 22158
rect 18172 22094 18174 22146
rect 18226 22094 18228 22146
rect 18172 21252 18228 22094
rect 18284 21924 18340 23102
rect 18284 21858 18340 21868
rect 18396 23154 18452 23166
rect 18396 23102 18398 23154
rect 18450 23102 18452 23154
rect 18396 21812 18452 23102
rect 18620 23044 18676 23436
rect 18732 23268 18788 23278
rect 18732 23174 18788 23212
rect 18844 23156 18900 24446
rect 18956 23380 19012 24668
rect 19068 24612 19124 24622
rect 19068 24162 19124 24556
rect 19180 24500 19236 24892
rect 19292 24724 19348 25228
rect 19404 25218 19460 25228
rect 19516 25282 19572 25294
rect 19516 25230 19518 25282
rect 19570 25230 19572 25282
rect 19516 25172 19572 25230
rect 19516 25106 19572 25116
rect 19628 25282 19684 25294
rect 19628 25230 19630 25282
rect 19682 25230 19684 25282
rect 19628 24948 19684 25230
rect 19852 25282 19908 26852
rect 19964 26516 20020 26526
rect 19964 26422 20020 26460
rect 19852 25230 19854 25282
rect 19906 25230 19908 25282
rect 19852 24948 19908 25230
rect 20188 26290 20244 26302
rect 20188 26238 20190 26290
rect 20242 26238 20244 26290
rect 20188 25060 20244 26238
rect 20412 26180 20468 26190
rect 20412 26086 20468 26124
rect 20524 25844 20580 26852
rect 20524 25778 20580 25788
rect 20636 26290 20692 26302
rect 20636 26238 20638 26290
rect 20690 26238 20692 26290
rect 20524 25620 20580 25630
rect 20636 25620 20692 26238
rect 20748 26292 20804 26302
rect 20748 26198 20804 26236
rect 20636 25564 20804 25620
rect 20300 25508 20356 25518
rect 20356 25452 20468 25508
rect 20300 25442 20356 25452
rect 20188 24994 20244 25004
rect 20300 25282 20356 25294
rect 20300 25230 20302 25282
rect 20354 25230 20356 25282
rect 19684 24892 19796 24948
rect 19628 24882 19684 24892
rect 19292 24630 19348 24668
rect 19516 24836 19572 24846
rect 19516 24722 19572 24780
rect 19516 24670 19518 24722
rect 19570 24670 19572 24722
rect 19404 24610 19460 24622
rect 19404 24558 19406 24610
rect 19458 24558 19460 24610
rect 19404 24500 19460 24558
rect 19180 24444 19460 24500
rect 19068 24110 19070 24162
rect 19122 24110 19124 24162
rect 19068 24098 19124 24110
rect 19404 24164 19460 24174
rect 18956 23314 19012 23324
rect 19180 24052 19236 24062
rect 19180 23938 19236 23996
rect 19180 23886 19182 23938
rect 19234 23886 19236 23938
rect 19068 23156 19124 23166
rect 18844 23154 19124 23156
rect 18844 23102 19070 23154
rect 19122 23102 19124 23154
rect 18844 23100 19124 23102
rect 19180 23156 19236 23886
rect 19292 23940 19348 23950
rect 19292 23714 19348 23884
rect 19292 23662 19294 23714
rect 19346 23662 19348 23714
rect 19292 23650 19348 23662
rect 19292 23156 19348 23166
rect 19180 23100 19292 23156
rect 19404 23156 19460 24108
rect 19516 23604 19572 24670
rect 19740 24724 19796 24892
rect 19852 24882 19908 24892
rect 20188 24836 20244 24846
rect 19964 24834 20244 24836
rect 19964 24782 20190 24834
rect 20242 24782 20244 24834
rect 19964 24780 20244 24782
rect 19740 23940 19796 24668
rect 19852 24722 19908 24734
rect 19852 24670 19854 24722
rect 19906 24670 19908 24722
rect 19852 24164 19908 24670
rect 19852 24098 19908 24108
rect 19852 23940 19908 23950
rect 19740 23938 19908 23940
rect 19740 23886 19854 23938
rect 19906 23886 19908 23938
rect 19740 23884 19908 23886
rect 19852 23874 19908 23884
rect 19628 23826 19684 23838
rect 19628 23774 19630 23826
rect 19682 23774 19684 23826
rect 19628 23716 19684 23774
rect 19628 23660 19908 23716
rect 19516 23548 19796 23604
rect 19404 23100 19684 23156
rect 19068 23090 19124 23100
rect 19292 23090 19348 23100
rect 18620 22988 18900 23044
rect 18396 21746 18452 21756
rect 18508 22820 18564 22830
rect 18396 21476 18452 21486
rect 18396 21382 18452 21420
rect 17612 21196 18228 21252
rect 18172 21140 18228 21196
rect 18172 21084 18452 21140
rect 17388 20862 17390 20914
rect 17442 20862 17444 20914
rect 17388 20850 17444 20862
rect 17836 20804 17892 20814
rect 17836 20710 17892 20748
rect 18284 20802 18340 20814
rect 18284 20750 18286 20802
rect 18338 20750 18340 20802
rect 17612 20690 17668 20702
rect 17612 20638 17614 20690
rect 17666 20638 17668 20690
rect 17612 20580 17668 20638
rect 17612 20514 17668 20524
rect 18060 20578 18116 20590
rect 18060 20526 18062 20578
rect 18114 20526 18116 20578
rect 17340 20412 17604 20422
rect 17396 20356 17444 20412
rect 17500 20356 17548 20412
rect 17340 20346 17604 20356
rect 17500 20244 17556 20254
rect 17500 20018 17556 20188
rect 18060 20132 18116 20526
rect 18284 20580 18340 20750
rect 18284 20514 18340 20524
rect 18172 20132 18228 20142
rect 18060 20130 18228 20132
rect 18060 20078 18174 20130
rect 18226 20078 18228 20130
rect 18060 20076 18228 20078
rect 18172 20066 18228 20076
rect 17500 19966 17502 20018
rect 17554 19966 17556 20018
rect 17500 19954 17556 19966
rect 17052 19346 17220 19348
rect 17052 19294 17054 19346
rect 17106 19294 17220 19346
rect 17052 19292 17220 19294
rect 17052 18676 17108 19292
rect 17500 19234 17556 19246
rect 17500 19182 17502 19234
rect 17554 19182 17556 19234
rect 17500 19012 17556 19182
rect 17724 19124 17780 19134
rect 17724 19030 17780 19068
rect 17500 18946 17556 18956
rect 18284 19012 18340 19022
rect 18284 18918 18340 18956
rect 18396 18900 18452 21084
rect 17340 18844 17604 18854
rect 17396 18788 17444 18844
rect 17500 18788 17548 18844
rect 18396 18834 18452 18844
rect 17340 18778 17604 18788
rect 17052 18610 17108 18620
rect 16828 17726 16830 17778
rect 16882 17726 16884 17778
rect 16828 17714 16884 17726
rect 17612 17892 17668 17902
rect 18508 17892 18564 22764
rect 18620 22594 18676 22606
rect 18620 22542 18622 22594
rect 18674 22542 18676 22594
rect 18620 22482 18676 22542
rect 18620 22430 18622 22482
rect 18674 22430 18676 22482
rect 18620 20020 18676 22430
rect 18844 22372 18900 22988
rect 19180 22932 19236 22942
rect 19516 22932 19572 22942
rect 19180 22930 19572 22932
rect 19180 22878 19182 22930
rect 19234 22878 19518 22930
rect 19570 22878 19572 22930
rect 19180 22876 19572 22878
rect 19180 22866 19236 22876
rect 19516 22866 19572 22876
rect 19628 22930 19684 23100
rect 19628 22878 19630 22930
rect 19682 22878 19684 22930
rect 18844 22278 18900 22316
rect 19068 22820 19124 22830
rect 19068 21700 19124 22764
rect 19180 22596 19236 22606
rect 19180 22370 19236 22540
rect 19628 22484 19684 22878
rect 19740 22932 19796 23548
rect 19852 23492 19908 23660
rect 19852 23426 19908 23436
rect 19964 23604 20020 24780
rect 20188 24770 20244 24780
rect 20300 24836 20356 25230
rect 20412 25060 20468 25452
rect 20524 25394 20580 25564
rect 20524 25342 20526 25394
rect 20578 25342 20580 25394
rect 20524 25330 20580 25342
rect 20636 25396 20692 25406
rect 20636 25302 20692 25340
rect 20636 25172 20692 25182
rect 20412 25004 20580 25060
rect 20300 24770 20356 24780
rect 20412 24724 20468 24734
rect 20412 24630 20468 24668
rect 20300 24612 20356 24622
rect 20300 24518 20356 24556
rect 20188 24500 20244 24510
rect 20076 23940 20132 23950
rect 20076 23846 20132 23884
rect 20076 23716 20132 23726
rect 20076 23622 20132 23660
rect 19964 23154 20020 23548
rect 19964 23102 19966 23154
rect 20018 23102 20020 23154
rect 19964 23090 20020 23102
rect 20188 23156 20244 24444
rect 20412 23940 20468 23950
rect 20524 23940 20580 25004
rect 20636 24722 20692 25116
rect 20636 24670 20638 24722
rect 20690 24670 20692 24722
rect 20636 24658 20692 24670
rect 20412 23938 20580 23940
rect 20412 23886 20414 23938
rect 20466 23886 20580 23938
rect 20412 23884 20580 23886
rect 20412 23874 20468 23884
rect 20636 23828 20692 23838
rect 20524 23772 20636 23828
rect 20412 23380 20468 23390
rect 20412 23286 20468 23324
rect 19852 22932 19908 22942
rect 19740 22876 19852 22932
rect 19852 22838 19908 22876
rect 20188 22820 20244 23100
rect 20188 22754 20244 22764
rect 19180 22318 19182 22370
rect 19234 22318 19236 22370
rect 19180 22306 19236 22318
rect 19404 22428 19684 22484
rect 19740 22596 19796 22606
rect 19404 22146 19460 22428
rect 19404 22094 19406 22146
rect 19458 22094 19460 22146
rect 19068 21634 19124 21644
rect 19180 21812 19236 21822
rect 18732 21588 18788 21598
rect 18732 20244 18788 21532
rect 19180 20802 19236 21756
rect 19404 21700 19460 22094
rect 19516 22148 19572 22158
rect 19516 22146 19684 22148
rect 19516 22094 19518 22146
rect 19570 22094 19684 22146
rect 19516 22092 19684 22094
rect 19516 22082 19572 22092
rect 19404 21634 19460 21644
rect 19516 21476 19572 21486
rect 19292 21474 19572 21476
rect 19292 21422 19518 21474
rect 19570 21422 19572 21474
rect 19292 21420 19572 21422
rect 19292 20914 19348 21420
rect 19516 21410 19572 21420
rect 19292 20862 19294 20914
rect 19346 20862 19348 20914
rect 19292 20850 19348 20862
rect 19180 20750 19182 20802
rect 19234 20750 19236 20802
rect 19180 20738 19236 20750
rect 19516 20804 19572 20814
rect 19628 20804 19684 22092
rect 19516 20802 19684 20804
rect 19516 20750 19518 20802
rect 19570 20750 19684 20802
rect 19516 20748 19684 20750
rect 19516 20738 19572 20748
rect 18844 20692 18900 20702
rect 18844 20598 18900 20636
rect 19740 20690 19796 22540
rect 19740 20638 19742 20690
rect 19794 20638 19796 20690
rect 19740 20626 19796 20638
rect 19852 22484 19908 22494
rect 19628 20580 19684 20590
rect 19628 20486 19684 20524
rect 19852 20356 19908 22428
rect 20524 22372 20580 23772
rect 20636 23762 20692 23772
rect 20636 23380 20692 23390
rect 20636 23154 20692 23324
rect 20748 23268 20804 25564
rect 20860 23492 20916 26852
rect 21196 26852 21364 26908
rect 21084 26740 21140 26750
rect 20972 26628 21028 26638
rect 20972 23828 21028 26572
rect 20972 23762 21028 23772
rect 21084 23604 21140 26684
rect 21196 25732 21252 26852
rect 21644 26850 21700 26862
rect 21644 26798 21646 26850
rect 21698 26798 21700 26850
rect 21644 26740 21700 26798
rect 21644 26674 21700 26684
rect 21644 26292 21700 26302
rect 21756 26292 21812 27244
rect 21644 26290 21812 26292
rect 21644 26238 21646 26290
rect 21698 26238 21812 26290
rect 21644 26236 21812 26238
rect 21644 26226 21700 26236
rect 21372 25900 21636 25910
rect 21428 25844 21476 25900
rect 21532 25844 21580 25900
rect 21372 25834 21636 25844
rect 21196 25676 21364 25732
rect 21196 25284 21252 25294
rect 21196 24722 21252 25228
rect 21196 24670 21198 24722
rect 21250 24670 21252 24722
rect 21196 24658 21252 24670
rect 21196 24500 21252 24510
rect 21308 24500 21364 25676
rect 21756 25396 21812 26236
rect 21868 26180 21924 28252
rect 22092 26516 22148 30046
rect 22316 29764 22372 29774
rect 22316 29650 22372 29708
rect 22316 29598 22318 29650
rect 22370 29598 22372 29650
rect 22316 29586 22372 29598
rect 22540 29708 23156 29764
rect 22540 29650 22596 29708
rect 22540 29598 22542 29650
rect 22594 29598 22596 29650
rect 22540 29586 22596 29598
rect 22988 29538 23044 29550
rect 22988 29486 22990 29538
rect 23042 29486 23044 29538
rect 22204 29426 22260 29438
rect 22204 29374 22206 29426
rect 22258 29374 22260 29426
rect 22204 29316 22260 29374
rect 22652 29428 22708 29438
rect 22204 29260 22484 29316
rect 22204 28642 22260 28654
rect 22204 28590 22206 28642
rect 22258 28590 22260 28642
rect 22204 27300 22260 28590
rect 22204 27234 22260 27244
rect 22316 28420 22372 28430
rect 22316 27186 22372 28364
rect 22316 27134 22318 27186
rect 22370 27134 22372 27186
rect 22316 27122 22372 27134
rect 22428 28420 22484 29260
rect 22652 28642 22708 29372
rect 22652 28590 22654 28642
rect 22706 28590 22708 28642
rect 22652 28578 22708 28590
rect 22764 29426 22820 29438
rect 22764 29374 22766 29426
rect 22818 29374 22820 29426
rect 22764 28420 22820 29374
rect 22876 29428 22932 29438
rect 22876 29334 22932 29372
rect 22988 29316 23044 29486
rect 23100 29538 23156 29708
rect 23100 29486 23102 29538
rect 23154 29486 23156 29538
rect 23100 29474 23156 29486
rect 23436 29426 23492 30156
rect 23436 29374 23438 29426
rect 23490 29374 23492 29426
rect 23436 29362 23492 29374
rect 23884 29316 23940 29326
rect 22988 29250 23044 29260
rect 23548 29314 23940 29316
rect 23548 29262 23886 29314
rect 23938 29262 23940 29314
rect 23548 29260 23940 29262
rect 23436 29204 23492 29214
rect 23436 28754 23492 29148
rect 23436 28702 23438 28754
rect 23490 28702 23492 28754
rect 23436 28690 23492 28702
rect 22428 28364 22820 28420
rect 22428 27188 22484 28364
rect 22428 27122 22484 27132
rect 23436 27188 23492 27198
rect 22092 26450 22148 26460
rect 23100 26404 23156 26414
rect 21868 26114 21924 26124
rect 22204 26180 22260 26190
rect 22204 25844 22260 26124
rect 22316 26178 22372 26190
rect 22316 26126 22318 26178
rect 22370 26126 22372 26178
rect 22316 26068 22372 26126
rect 22316 26002 22372 26012
rect 22204 25788 22372 25844
rect 22092 25732 22148 25742
rect 22148 25676 22260 25732
rect 22092 25666 22148 25676
rect 21980 25396 22036 25406
rect 21756 25394 22036 25396
rect 21756 25342 21982 25394
rect 22034 25342 22036 25394
rect 21756 25340 22036 25342
rect 21980 25284 22036 25340
rect 21252 24444 21364 24500
rect 21868 24610 21924 24622
rect 21868 24558 21870 24610
rect 21922 24558 21924 24610
rect 21196 24434 21252 24444
rect 21372 24332 21636 24342
rect 21196 24276 21252 24286
rect 21428 24276 21476 24332
rect 21532 24276 21580 24332
rect 21372 24266 21636 24276
rect 21196 23828 21252 24220
rect 21308 23828 21364 23838
rect 21196 23826 21364 23828
rect 21196 23774 21310 23826
rect 21362 23774 21364 23826
rect 21196 23772 21364 23774
rect 21308 23762 21364 23772
rect 21644 23714 21700 23726
rect 21644 23662 21646 23714
rect 21698 23662 21700 23714
rect 21084 23548 21252 23604
rect 20860 23426 20916 23436
rect 20748 23212 21028 23268
rect 20636 23102 20638 23154
rect 20690 23102 20692 23154
rect 20636 22484 20692 23102
rect 20860 23044 20916 23054
rect 20748 22596 20804 22606
rect 20748 22502 20804 22540
rect 20636 22418 20692 22428
rect 20524 22306 20580 22316
rect 20636 22260 20692 22270
rect 19964 22148 20020 22158
rect 20412 22148 20468 22158
rect 20636 22148 20692 22204
rect 19964 22146 20692 22148
rect 19964 22094 19966 22146
rect 20018 22094 20414 22146
rect 20466 22094 20692 22146
rect 19964 22092 20692 22094
rect 19964 22082 20020 22092
rect 20412 22082 20468 22092
rect 19964 21924 20020 21934
rect 19964 20804 20020 21868
rect 20524 21476 20580 21486
rect 20300 20804 20356 20814
rect 19964 20802 20132 20804
rect 19964 20750 19966 20802
rect 20018 20750 20132 20802
rect 19964 20748 20132 20750
rect 19964 20738 20020 20748
rect 18732 20178 18788 20188
rect 19740 20300 19908 20356
rect 20076 20356 20132 20748
rect 20300 20802 20468 20804
rect 20300 20750 20302 20802
rect 20354 20750 20468 20802
rect 20300 20748 20468 20750
rect 20300 20738 20356 20748
rect 20076 20300 20244 20356
rect 18620 19964 18900 20020
rect 18844 19458 18900 19964
rect 18844 19406 18846 19458
rect 18898 19406 18900 19458
rect 18844 19394 18900 19406
rect 19404 19908 19460 19918
rect 19068 19348 19124 19358
rect 19068 19254 19124 19292
rect 19404 19346 19460 19852
rect 19404 19294 19406 19346
rect 19458 19294 19460 19346
rect 18620 18676 18676 18686
rect 18620 18582 18676 18620
rect 19404 18676 19460 19294
rect 19460 18620 19684 18676
rect 19404 18610 19460 18620
rect 19068 18564 19124 18574
rect 18956 18340 19012 18350
rect 18732 18338 19012 18340
rect 18732 18286 18958 18338
rect 19010 18286 19012 18338
rect 18732 18284 19012 18286
rect 18620 17892 18676 17902
rect 18508 17836 18620 17892
rect 17612 17778 17668 17836
rect 18620 17826 18676 17836
rect 17836 17780 17892 17790
rect 17612 17726 17614 17778
rect 17666 17726 17668 17778
rect 17612 17714 17668 17726
rect 17724 17778 17892 17780
rect 17724 17726 17838 17778
rect 17890 17726 17892 17778
rect 17724 17724 17892 17726
rect 16716 17490 16772 17500
rect 17340 17276 17604 17286
rect 17396 17220 17444 17276
rect 17500 17220 17548 17276
rect 17340 17210 17604 17220
rect 16828 16884 16884 16894
rect 16828 16790 16884 16828
rect 15036 16258 15092 16268
rect 16940 16210 16996 16222
rect 16940 16158 16942 16210
rect 16994 16158 16996 16210
rect 16380 16100 16436 16110
rect 16380 16098 16772 16100
rect 16380 16046 16382 16098
rect 16434 16046 16772 16098
rect 16380 16044 16772 16046
rect 16380 16034 16436 16044
rect 16716 15988 16772 16044
rect 16828 15988 16884 15998
rect 16716 15986 16884 15988
rect 16716 15934 16830 15986
rect 16882 15934 16884 15986
rect 16716 15932 16884 15934
rect 16604 15874 16660 15886
rect 16604 15822 16606 15874
rect 16658 15822 16660 15874
rect 16604 15652 16660 15822
rect 16380 15596 16660 15652
rect 14084 15372 14196 15428
rect 14700 15428 14756 15438
rect 14028 15362 14084 15372
rect 12012 15202 12292 15204
rect 12012 15150 12014 15202
rect 12066 15150 12238 15202
rect 12290 15150 12292 15202
rect 12012 15148 12292 15150
rect 12460 15148 12628 15204
rect 12684 15314 13188 15316
rect 12684 15262 13134 15314
rect 13186 15262 13188 15314
rect 12684 15260 13188 15262
rect 12012 15138 12068 15148
rect 12236 15092 12404 15148
rect 11900 14532 11956 14542
rect 11900 14530 12180 14532
rect 11900 14478 11902 14530
rect 11954 14478 12180 14530
rect 11900 14476 12180 14478
rect 11900 14466 11956 14476
rect 11564 14308 11620 14318
rect 11564 13858 11620 14252
rect 11564 13806 11566 13858
rect 11618 13806 11620 13858
rect 11564 13794 11620 13806
rect 12012 13972 12068 13982
rect 11900 13748 11956 13758
rect 12012 13748 12068 13916
rect 11900 13746 12068 13748
rect 11900 13694 11902 13746
rect 11954 13694 12068 13746
rect 11900 13692 12068 13694
rect 11900 13682 11956 13692
rect 11676 13634 11732 13646
rect 11676 13582 11678 13634
rect 11730 13582 11732 13634
rect 11676 13524 11732 13582
rect 11676 13458 11732 13468
rect 12124 12852 12180 14476
rect 12236 14308 12292 14318
rect 12236 14214 12292 14252
rect 10892 11732 10948 11742
rect 10444 11396 10500 11406
rect 10220 11394 10500 11396
rect 10220 11342 10446 11394
rect 10498 11342 10500 11394
rect 10220 11340 10500 11342
rect 9884 11172 9940 11182
rect 9276 11004 9540 11014
rect 9332 10948 9380 11004
rect 9436 10948 9484 11004
rect 9276 10938 9540 10948
rect 9660 10724 9716 10734
rect 9212 9828 9268 9838
rect 8764 9762 8820 9772
rect 8876 9826 9268 9828
rect 8876 9774 9214 9826
rect 9266 9774 9268 9826
rect 8876 9772 9268 9774
rect 8652 9716 8708 9726
rect 8652 9622 8708 9660
rect 8764 9602 8820 9614
rect 8764 9550 8766 9602
rect 8818 9550 8820 9602
rect 8764 9492 8820 9550
rect 8540 9436 8820 9492
rect 8428 9324 8820 9380
rect 8540 7588 8596 7598
rect 8204 7422 8206 7474
rect 8258 7422 8260 7474
rect 8204 7410 8260 7422
rect 8316 7586 8596 7588
rect 8316 7534 8542 7586
rect 8594 7534 8596 7586
rect 8316 7532 8596 7534
rect 8316 7476 8372 7532
rect 8540 7522 8596 7532
rect 7420 6804 7476 6972
rect 8316 6804 8372 7420
rect 8764 7474 8820 9324
rect 8876 9042 8932 9772
rect 9212 9762 9268 9772
rect 8876 8990 8878 9042
rect 8930 8990 8932 9042
rect 8876 8372 8932 8990
rect 9100 9604 9156 9614
rect 8876 8370 9044 8372
rect 8876 8318 8878 8370
rect 8930 8318 9044 8370
rect 8876 8316 9044 8318
rect 8876 8306 8932 8316
rect 8764 7422 8766 7474
rect 8818 7422 8820 7474
rect 8764 7410 8820 7422
rect 7420 6738 7476 6748
rect 8204 6748 8372 6804
rect 8428 7252 8484 7262
rect 6860 6466 6916 6478
rect 6860 6414 6862 6466
rect 6914 6414 6916 6466
rect 6860 5124 6916 6414
rect 8092 6244 8148 6254
rect 8092 6018 8148 6188
rect 8092 5966 8094 6018
rect 8146 5966 8148 6018
rect 8092 5954 8148 5966
rect 6860 5058 6916 5068
rect 5740 3390 5742 3442
rect 5794 3390 5796 3442
rect 5740 3378 5796 3390
rect 5852 3388 5908 3398
rect 6524 3388 6580 4956
rect 5852 3386 6132 3388
rect 5852 3334 5854 3386
rect 5906 3334 6132 3386
rect 5852 3332 6132 3334
rect 6188 3332 6580 3388
rect 7084 5010 7140 5022
rect 7084 4958 7086 5010
rect 7138 4958 7140 5010
rect 7084 3388 7140 4958
rect 8204 4562 8260 6748
rect 8428 5348 8484 7196
rect 8204 4510 8206 4562
rect 8258 4510 8260 4562
rect 8204 4498 8260 4510
rect 8316 5292 8484 5348
rect 8764 6804 8820 6814
rect 8764 6466 8820 6748
rect 8764 6414 8766 6466
rect 8818 6414 8820 6466
rect 8316 4562 8372 5292
rect 8316 4510 8318 4562
rect 8370 4510 8372 4562
rect 8316 4498 8372 4510
rect 8428 5122 8484 5134
rect 8428 5070 8430 5122
rect 8482 5070 8484 5122
rect 7868 4340 7924 4350
rect 7868 4226 7924 4284
rect 8428 4340 8484 5070
rect 8428 4246 8484 4284
rect 8764 4338 8820 6414
rect 8876 5908 8932 5918
rect 8988 5908 9044 8316
rect 9100 6692 9156 9548
rect 9660 9604 9716 10668
rect 9884 9716 9940 11116
rect 10444 11060 10500 11340
rect 10892 11172 10948 11676
rect 11452 11508 11508 12348
rect 11900 12796 12180 12852
rect 10892 11078 10948 11116
rect 11004 11506 11508 11508
rect 11004 11454 11454 11506
rect 11506 11454 11508 11506
rect 11004 11452 11508 11454
rect 10444 11004 10724 11060
rect 10668 10836 10724 11004
rect 10556 10610 10612 10622
rect 10556 10558 10558 10610
rect 10610 10558 10612 10610
rect 9996 10500 10052 10510
rect 9996 9938 10052 10444
rect 9996 9886 9998 9938
rect 10050 9886 10052 9938
rect 9996 9874 10052 9886
rect 10444 10498 10500 10510
rect 10444 10446 10446 10498
rect 10498 10446 10500 10498
rect 9884 9660 10052 9716
rect 9660 9538 9716 9548
rect 9276 9436 9540 9446
rect 9332 9380 9380 9436
rect 9436 9380 9484 9436
rect 9276 9370 9540 9380
rect 9660 9268 9716 9278
rect 9660 9266 9940 9268
rect 9660 9214 9662 9266
rect 9714 9214 9940 9266
rect 9660 9212 9940 9214
rect 9660 9202 9716 9212
rect 9772 9042 9828 9054
rect 9772 8990 9774 9042
rect 9826 8990 9828 9042
rect 9772 8932 9828 8990
rect 9772 8866 9828 8876
rect 9660 8818 9716 8830
rect 9660 8766 9662 8818
rect 9714 8766 9716 8818
rect 9276 7868 9540 7878
rect 9332 7812 9380 7868
rect 9436 7812 9484 7868
rect 9276 7802 9540 7812
rect 9100 6626 9156 6636
rect 9212 7700 9268 7710
rect 9100 6468 9156 6478
rect 9212 6468 9268 7644
rect 9548 7362 9604 7374
rect 9548 7310 9550 7362
rect 9602 7310 9604 7362
rect 9436 6916 9492 6926
rect 9436 6578 9492 6860
rect 9436 6526 9438 6578
rect 9490 6526 9492 6578
rect 9436 6514 9492 6526
rect 9548 6580 9604 7310
rect 9660 6916 9716 8766
rect 9660 6850 9716 6860
rect 9660 6692 9716 6702
rect 9660 6598 9716 6636
rect 9548 6514 9604 6524
rect 9100 6466 9268 6468
rect 9100 6414 9102 6466
rect 9154 6414 9268 6466
rect 9100 6412 9268 6414
rect 9884 6468 9940 9212
rect 9996 7700 10052 9660
rect 10444 9492 10500 10446
rect 10444 9426 10500 9436
rect 10556 9268 10612 10558
rect 10668 10276 10724 10780
rect 11004 10722 11060 11452
rect 11452 11442 11508 11452
rect 11564 11620 11620 11630
rect 11564 10834 11620 11564
rect 11900 10948 11956 12796
rect 12124 12516 12180 12526
rect 12180 12460 12292 12516
rect 12124 12450 12180 12460
rect 12236 12402 12292 12460
rect 12236 12350 12238 12402
rect 12290 12350 12292 12402
rect 12012 12292 12068 12302
rect 12012 12178 12068 12236
rect 12012 12126 12014 12178
rect 12066 12126 12068 12178
rect 12012 12114 12068 12126
rect 12236 11620 12292 12350
rect 12348 12292 12404 15092
rect 12460 13972 12516 15148
rect 12572 14532 12628 14542
rect 12684 14532 12740 15260
rect 13132 15250 13188 15260
rect 13692 15314 13748 15326
rect 13692 15262 13694 15314
rect 13746 15262 13748 15314
rect 13308 14924 13572 14934
rect 13364 14868 13412 14924
rect 13468 14868 13516 14924
rect 13308 14858 13572 14868
rect 12572 14530 12740 14532
rect 12572 14478 12574 14530
rect 12626 14478 12740 14530
rect 12572 14476 12740 14478
rect 13580 14532 13636 14542
rect 13692 14532 13748 15262
rect 14476 15202 14532 15214
rect 14476 15150 14478 15202
rect 14530 15150 14532 15202
rect 14476 14644 14532 15150
rect 14476 14578 14532 14588
rect 13580 14530 13748 14532
rect 13580 14478 13582 14530
rect 13634 14478 13748 14530
rect 13580 14476 13748 14478
rect 12572 14466 12628 14476
rect 13580 14466 13636 14476
rect 12460 13878 12516 13916
rect 12572 14308 12628 14318
rect 12572 12516 12628 14252
rect 12908 13748 12964 13758
rect 12908 13074 12964 13692
rect 13308 13356 13572 13366
rect 13364 13300 13412 13356
rect 13468 13300 13516 13356
rect 13308 13290 13572 13300
rect 12908 13022 12910 13074
rect 12962 13022 12964 13074
rect 12908 13010 12964 13022
rect 13356 13076 13412 13086
rect 12348 12226 12404 12236
rect 12460 12460 12628 12516
rect 12236 11396 12292 11564
rect 12236 11330 12292 11340
rect 11900 10892 12292 10948
rect 11564 10782 11566 10834
rect 11618 10782 11620 10834
rect 11564 10770 11620 10782
rect 11004 10670 11006 10722
rect 11058 10670 11060 10722
rect 11004 10658 11060 10670
rect 11900 10722 11956 10734
rect 11900 10670 11902 10722
rect 11954 10670 11956 10722
rect 11228 10612 11284 10622
rect 11228 10610 11508 10612
rect 11228 10558 11230 10610
rect 11282 10558 11508 10610
rect 11228 10556 11508 10558
rect 11228 10546 11284 10556
rect 10780 10500 10836 10510
rect 10780 10406 10836 10444
rect 10668 10220 10836 10276
rect 10668 9268 10724 9278
rect 10332 9266 10724 9268
rect 10332 9214 10670 9266
rect 10722 9214 10724 9266
rect 10332 9212 10724 9214
rect 10220 9156 10276 9166
rect 10220 9062 10276 9100
rect 9996 7634 10052 7644
rect 10108 9042 10164 9054
rect 10108 8990 10110 9042
rect 10162 8990 10164 9042
rect 10108 8932 10164 8990
rect 10332 8932 10388 9212
rect 10668 9202 10724 9212
rect 10444 9044 10500 9054
rect 10444 9042 10612 9044
rect 10444 8990 10446 9042
rect 10498 8990 10612 9042
rect 10444 8988 10612 8990
rect 10444 8978 10500 8988
rect 10108 8876 10388 8932
rect 10108 6580 10164 8876
rect 10556 6692 10612 8988
rect 10780 8820 10836 10220
rect 10892 9492 10948 9502
rect 10892 9044 10948 9436
rect 11452 9266 11508 10556
rect 11452 9214 11454 9266
rect 11506 9214 11508 9266
rect 11452 9202 11508 9214
rect 11900 9604 11956 10670
rect 12236 10610 12292 10892
rect 12236 10558 12238 10610
rect 12290 10558 12292 10610
rect 12124 9940 12180 9950
rect 11564 9156 11620 9166
rect 10892 8950 10948 8988
rect 11340 9044 11396 9054
rect 11340 8950 11396 8988
rect 11564 9042 11620 9100
rect 11564 8990 11566 9042
rect 11618 8990 11620 9042
rect 10780 8754 10836 8764
rect 11564 8484 11620 8990
rect 11900 9042 11956 9548
rect 11900 8990 11902 9042
rect 11954 8990 11956 9042
rect 11900 8978 11956 8990
rect 12012 9938 12180 9940
rect 12012 9886 12126 9938
rect 12178 9886 12180 9938
rect 12012 9884 12180 9886
rect 11564 8418 11620 8428
rect 11788 8932 11844 8942
rect 11676 8260 11732 8270
rect 11676 8166 11732 8204
rect 10780 7364 10836 7374
rect 11676 7364 11732 7374
rect 10668 6692 10724 6702
rect 10556 6690 10724 6692
rect 10556 6638 10670 6690
rect 10722 6638 10724 6690
rect 10556 6636 10724 6638
rect 10668 6626 10724 6636
rect 10220 6580 10276 6590
rect 10108 6578 10276 6580
rect 10108 6526 10222 6578
rect 10274 6526 10276 6578
rect 10108 6524 10276 6526
rect 9100 6402 9156 6412
rect 9660 6356 9716 6366
rect 9276 6300 9540 6310
rect 9332 6244 9380 6300
rect 9436 6244 9484 6300
rect 9276 6234 9540 6244
rect 9660 6018 9716 6300
rect 9660 5966 9662 6018
rect 9714 5966 9716 6018
rect 9660 5954 9716 5966
rect 9772 6020 9828 6030
rect 9772 5926 9828 5964
rect 8876 5906 9044 5908
rect 8876 5854 8878 5906
rect 8930 5854 9044 5906
rect 8876 5852 9044 5854
rect 8876 5842 8932 5852
rect 8988 5122 9044 5852
rect 9772 5684 9828 5694
rect 9772 5590 9828 5628
rect 9772 5236 9828 5246
rect 9772 5142 9828 5180
rect 8988 5070 8990 5122
rect 9042 5070 9044 5122
rect 8988 5058 9044 5070
rect 9276 4732 9540 4742
rect 9332 4676 9380 4732
rect 9436 4676 9484 4732
rect 9276 4666 9540 4676
rect 8764 4286 8766 4338
rect 8818 4286 8820 4338
rect 8764 4274 8820 4286
rect 7868 4174 7870 4226
rect 7922 4174 7924 4226
rect 7868 3444 7924 4174
rect 7084 3332 7252 3388
rect 7868 3378 7924 3388
rect 8540 3666 8596 3678
rect 8540 3614 8542 3666
rect 8594 3614 8596 3666
rect 8540 3388 8596 3614
rect 9548 3668 9604 3678
rect 9884 3668 9940 6412
rect 10220 6356 10276 6524
rect 10332 6580 10388 6590
rect 10332 6486 10388 6524
rect 10220 6290 10276 6300
rect 10556 6466 10612 6478
rect 10556 6414 10558 6466
rect 10610 6414 10612 6466
rect 10444 6020 10500 6030
rect 10556 6020 10612 6414
rect 10444 6018 10612 6020
rect 10444 5966 10446 6018
rect 10498 5966 10612 6018
rect 10444 5964 10612 5966
rect 10780 6018 10836 7308
rect 10892 7362 11732 7364
rect 10892 7310 11678 7362
rect 11730 7310 11732 7362
rect 10892 7308 11732 7310
rect 10892 6802 10948 7308
rect 11676 7298 11732 7308
rect 10892 6750 10894 6802
rect 10946 6750 10948 6802
rect 10892 6738 10948 6750
rect 11788 6804 11844 8876
rect 12012 8484 12068 9884
rect 12124 9874 12180 9884
rect 12236 9156 12292 10558
rect 12460 9268 12516 12460
rect 12572 12290 12628 12302
rect 12572 12238 12574 12290
rect 12626 12238 12628 12290
rect 12572 11732 12628 12238
rect 12796 12292 12852 12302
rect 12796 12180 12852 12236
rect 13356 12292 13412 13020
rect 13580 12964 13636 12974
rect 13692 12964 13748 14476
rect 13580 12962 13748 12964
rect 13580 12910 13582 12962
rect 13634 12910 13748 12962
rect 13580 12908 13748 12910
rect 14028 14420 14084 14430
rect 13580 12292 13636 12908
rect 13692 12292 13748 12302
rect 13580 12290 13748 12292
rect 13580 12238 13694 12290
rect 13746 12238 13748 12290
rect 13580 12236 13748 12238
rect 13356 12198 13412 12236
rect 12572 11666 12628 11676
rect 12684 12178 12852 12180
rect 12684 12126 12798 12178
rect 12850 12126 12852 12178
rect 12684 12124 12852 12126
rect 12572 11508 12628 11518
rect 12684 11508 12740 12124
rect 12796 12114 12852 12124
rect 13308 11788 13572 11798
rect 13132 11732 13188 11742
rect 13364 11732 13412 11788
rect 13468 11732 13516 11788
rect 13308 11722 13572 11732
rect 12572 11506 12740 11508
rect 12572 11454 12574 11506
rect 12626 11454 12740 11506
rect 12572 11452 12740 11454
rect 12796 11620 12852 11630
rect 12572 11442 12628 11452
rect 12572 9940 12628 9950
rect 12796 9940 12852 11564
rect 13020 10498 13076 10510
rect 13020 10446 13022 10498
rect 13074 10446 13076 10498
rect 13020 9940 13076 10446
rect 12572 9938 12964 9940
rect 12572 9886 12574 9938
rect 12626 9886 12964 9938
rect 12572 9884 12964 9886
rect 12572 9874 12628 9884
rect 12908 9492 12964 9884
rect 13020 9874 13076 9884
rect 13132 9828 13188 11676
rect 13468 11396 13524 11406
rect 13468 11302 13524 11340
rect 13692 11396 13748 12236
rect 14028 12290 14084 14364
rect 14252 14418 14308 14430
rect 14252 14366 14254 14418
rect 14306 14366 14308 14418
rect 14140 13972 14196 13982
rect 14252 13972 14308 14366
rect 14140 13970 14308 13972
rect 14140 13918 14142 13970
rect 14194 13918 14308 13970
rect 14140 13916 14308 13918
rect 14476 14308 14532 14318
rect 14140 13906 14196 13916
rect 14476 13858 14532 14252
rect 14476 13806 14478 13858
rect 14530 13806 14532 13858
rect 14476 13794 14532 13806
rect 14252 12852 14308 12862
rect 14252 12850 14644 12852
rect 14252 12798 14254 12850
rect 14306 12798 14644 12850
rect 14252 12796 14644 12798
rect 14252 12786 14308 12796
rect 14588 12402 14644 12796
rect 14588 12350 14590 12402
rect 14642 12350 14644 12402
rect 14588 12338 14644 12350
rect 14028 12238 14030 12290
rect 14082 12238 14084 12290
rect 14028 12226 14084 12238
rect 13692 11330 13748 11340
rect 13804 11170 13860 11182
rect 14252 11172 14308 11182
rect 13804 11118 13806 11170
rect 13858 11118 13860 11170
rect 13308 10220 13572 10230
rect 13364 10164 13412 10220
rect 13468 10164 13516 10220
rect 13308 10154 13572 10164
rect 13804 10052 13860 11118
rect 13804 9986 13860 9996
rect 14028 11170 14308 11172
rect 14028 11118 14254 11170
rect 14306 11118 14308 11170
rect 14028 11116 14308 11118
rect 14700 11172 14756 15372
rect 16380 14756 16436 15596
rect 16604 15428 16660 15438
rect 16604 15202 16660 15372
rect 16604 15150 16606 15202
rect 16658 15150 16660 15202
rect 16604 15138 16660 15150
rect 16828 14980 16884 15932
rect 16828 14914 16884 14924
rect 16380 14642 16436 14700
rect 16380 14590 16382 14642
rect 16434 14590 16436 14642
rect 16380 14578 16436 14590
rect 16940 14532 16996 16158
rect 16940 14466 16996 14476
rect 17052 15986 17108 15998
rect 17052 15934 17054 15986
rect 17106 15934 17108 15986
rect 15148 14420 15204 14430
rect 15148 13970 15204 14364
rect 16828 14308 16884 14318
rect 16828 14214 16884 14252
rect 15148 13918 15150 13970
rect 15202 13918 15204 13970
rect 15148 13906 15204 13918
rect 17052 13972 17108 15934
rect 17612 15988 17668 15998
rect 17612 15894 17668 15932
rect 17340 15708 17604 15718
rect 17396 15652 17444 15708
rect 17500 15652 17548 15708
rect 17340 15642 17604 15652
rect 17164 15316 17220 15326
rect 17164 14756 17220 15260
rect 17724 15148 17780 17724
rect 17836 17714 17892 17724
rect 18508 17668 18564 17678
rect 18732 17668 18788 18284
rect 18956 18274 19012 18284
rect 19068 18004 19124 18508
rect 18508 17666 18732 17668
rect 18508 17614 18510 17666
rect 18562 17614 18732 17666
rect 18508 17612 18732 17614
rect 18508 17602 18564 17612
rect 18732 17574 18788 17612
rect 18844 17948 19124 18004
rect 19180 18226 19236 18238
rect 19516 18228 19572 18238
rect 19180 18174 19182 18226
rect 19234 18174 19236 18226
rect 18172 17554 18228 17566
rect 18172 17502 18174 17554
rect 18226 17502 18228 17554
rect 17948 17444 18004 17454
rect 17948 17442 18116 17444
rect 17948 17390 17950 17442
rect 18002 17390 18116 17442
rect 17948 17388 18116 17390
rect 17948 17378 18004 17388
rect 17948 17220 18004 17230
rect 17948 16884 18004 17164
rect 17836 16100 17892 16110
rect 17836 15986 17892 16044
rect 17836 15934 17838 15986
rect 17890 15934 17892 15986
rect 17836 15922 17892 15934
rect 17948 15986 18004 16828
rect 18060 16324 18116 17388
rect 18172 16660 18228 17502
rect 18844 17554 18900 17948
rect 18844 17502 18846 17554
rect 18898 17502 18900 17554
rect 18172 16594 18228 16604
rect 18620 17444 18676 17454
rect 18508 16324 18564 16334
rect 18620 16324 18676 17388
rect 18844 16772 18900 17502
rect 18844 16706 18900 16716
rect 18956 17668 19012 17678
rect 19180 17668 19236 18174
rect 18956 17666 19236 17668
rect 18956 17614 18958 17666
rect 19010 17614 19236 17666
rect 18956 17612 19236 17614
rect 19292 18226 19572 18228
rect 19292 18174 19518 18226
rect 19570 18174 19572 18226
rect 19292 18172 19572 18174
rect 18060 16268 18452 16324
rect 17948 15934 17950 15986
rect 18002 15934 18004 15986
rect 17836 15540 17892 15550
rect 17836 15446 17892 15484
rect 17948 15428 18004 15934
rect 18060 15874 18116 15886
rect 18060 15822 18062 15874
rect 18114 15822 18116 15874
rect 18060 15540 18116 15822
rect 18172 15876 18228 15886
rect 18172 15782 18228 15820
rect 18060 15474 18116 15484
rect 17948 15362 18004 15372
rect 18396 15426 18452 16268
rect 18508 16322 18676 16324
rect 18508 16270 18510 16322
rect 18562 16270 18676 16322
rect 18508 16268 18676 16270
rect 18732 16660 18788 16670
rect 18508 16258 18564 16268
rect 18732 16210 18788 16604
rect 18956 16436 19012 17612
rect 18732 16158 18734 16210
rect 18786 16158 18788 16210
rect 18732 16146 18788 16158
rect 18844 16380 19012 16436
rect 18620 16098 18676 16110
rect 18620 16046 18622 16098
rect 18674 16046 18676 16098
rect 18620 15876 18676 16046
rect 18508 15540 18564 15578
rect 18508 15474 18564 15484
rect 18396 15374 18398 15426
rect 18450 15374 18452 15426
rect 18396 15362 18452 15374
rect 18172 15314 18228 15326
rect 18172 15262 18174 15314
rect 18226 15262 18228 15314
rect 17724 15092 18004 15148
rect 17164 14662 17220 14700
rect 17836 14980 17892 14990
rect 17836 14418 17892 14924
rect 17948 14756 18004 15092
rect 18172 14980 18228 15262
rect 18284 15316 18340 15326
rect 18284 15222 18340 15260
rect 18508 15316 18564 15326
rect 18508 15148 18564 15260
rect 18620 15204 18676 15820
rect 18844 15764 18900 16380
rect 19292 16322 19348 18172
rect 19516 18162 19572 18172
rect 19628 17554 19684 18620
rect 19740 18228 19796 20300
rect 20076 20132 20132 20142
rect 19964 19458 20020 19470
rect 19964 19406 19966 19458
rect 20018 19406 20020 19458
rect 19964 19346 20020 19406
rect 19964 19294 19966 19346
rect 20018 19294 20020 19346
rect 19964 19282 20020 19294
rect 19964 18564 20020 18574
rect 19964 18470 20020 18508
rect 19852 18452 19908 18462
rect 19852 18358 19908 18396
rect 19964 18228 20020 18238
rect 19740 18226 20020 18228
rect 19740 18174 19966 18226
rect 20018 18174 20020 18226
rect 19740 18172 20020 18174
rect 19964 18162 20020 18172
rect 19964 18004 20020 18014
rect 19628 17502 19630 17554
rect 19682 17502 19684 17554
rect 19404 17444 19460 17454
rect 19404 17350 19460 17388
rect 19516 17442 19572 17454
rect 19516 17390 19518 17442
rect 19570 17390 19572 17442
rect 19292 16270 19294 16322
rect 19346 16270 19348 16322
rect 19292 16258 19348 16270
rect 19404 16548 19460 16558
rect 19068 16100 19124 16110
rect 19068 16006 19124 16044
rect 19292 15876 19348 15886
rect 18844 15698 18900 15708
rect 19068 15820 19292 15876
rect 18844 15540 18900 15550
rect 18732 15428 18788 15438
rect 18732 15334 18788 15372
rect 18620 15148 18788 15204
rect 18172 14914 18228 14924
rect 18396 15092 18564 15148
rect 17948 14700 18340 14756
rect 17836 14366 17838 14418
rect 17890 14366 17892 14418
rect 17836 14196 17892 14366
rect 17340 14140 17604 14150
rect 17396 14084 17444 14140
rect 17500 14084 17548 14140
rect 17836 14130 17892 14140
rect 17948 14530 18004 14542
rect 17948 14478 17950 14530
rect 18002 14478 18004 14530
rect 17340 14074 17604 14084
rect 17052 13906 17108 13916
rect 17836 13970 17892 13982
rect 17836 13918 17838 13970
rect 17890 13918 17892 13970
rect 16604 13858 16660 13870
rect 16604 13806 16606 13858
rect 16658 13806 16660 13858
rect 14812 13748 14868 13758
rect 14812 13654 14868 13692
rect 15932 13636 15988 13646
rect 15932 13542 15988 13580
rect 16380 13636 16436 13646
rect 14924 13524 14980 13534
rect 14924 12290 14980 13468
rect 15596 13524 15652 13534
rect 15596 13430 15652 13468
rect 16380 13074 16436 13580
rect 16380 13022 16382 13074
rect 16434 13022 16436 13074
rect 16380 13010 16436 13022
rect 16604 12964 16660 13806
rect 16716 13860 16772 13870
rect 16716 13746 16772 13804
rect 16716 13694 16718 13746
rect 16770 13694 16772 13746
rect 16716 13682 16772 13694
rect 17612 13748 17668 13758
rect 17612 13654 17668 13692
rect 17724 13746 17780 13758
rect 17724 13694 17726 13746
rect 17778 13694 17780 13746
rect 17724 13524 17780 13694
rect 17724 13458 17780 13468
rect 16604 12898 16660 12908
rect 17164 12964 17220 12974
rect 17164 12870 17220 12908
rect 17340 12572 17604 12582
rect 17396 12516 17444 12572
rect 17500 12516 17548 12572
rect 17340 12506 17604 12516
rect 14924 12238 14926 12290
rect 14978 12238 14980 12290
rect 14924 12226 14980 12238
rect 16716 11956 16772 11966
rect 16716 11508 16772 11900
rect 16716 11442 16772 11452
rect 17836 11506 17892 13918
rect 17948 13186 18004 14478
rect 18284 14530 18340 14700
rect 18284 14478 18286 14530
rect 18338 14478 18340 14530
rect 18284 14466 18340 14478
rect 18396 14308 18452 15092
rect 18508 14644 18564 14654
rect 18508 14550 18564 14588
rect 18620 14532 18676 14542
rect 18620 14438 18676 14476
rect 18172 14252 18452 14308
rect 18732 14308 18788 15148
rect 18172 13746 18228 14252
rect 18732 14242 18788 14252
rect 18508 13972 18564 13982
rect 18508 13878 18564 13916
rect 18172 13694 18174 13746
rect 18226 13694 18228 13746
rect 18172 13682 18228 13694
rect 18396 13746 18452 13758
rect 18396 13694 18398 13746
rect 18450 13694 18452 13746
rect 18396 13300 18452 13694
rect 18732 13748 18788 13758
rect 18844 13748 18900 15484
rect 19068 15538 19124 15820
rect 19292 15810 19348 15820
rect 19068 15486 19070 15538
rect 19122 15486 19124 15538
rect 19068 15474 19124 15486
rect 19292 15540 19348 15550
rect 19292 15446 19348 15484
rect 19404 15426 19460 16492
rect 19404 15374 19406 15426
rect 19458 15374 19460 15426
rect 19404 15204 19460 15374
rect 19404 15138 19460 15148
rect 19516 14980 19572 17390
rect 19628 17220 19684 17502
rect 19852 17666 19908 17678
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19852 17444 19908 17614
rect 19964 17554 20020 17948
rect 19964 17502 19966 17554
rect 20018 17502 20020 17554
rect 19964 17490 20020 17502
rect 19852 17378 19908 17388
rect 19628 17154 19684 17164
rect 20076 16996 20132 20076
rect 20188 19908 20244 20300
rect 20300 19908 20356 19918
rect 20188 19906 20356 19908
rect 20188 19854 20302 19906
rect 20354 19854 20356 19906
rect 20188 19852 20356 19854
rect 20300 19842 20356 19852
rect 20300 19458 20356 19470
rect 20300 19406 20302 19458
rect 20354 19406 20356 19458
rect 20300 19348 20356 19406
rect 20300 19254 20356 19292
rect 20412 19124 20468 20748
rect 20524 20188 20580 21420
rect 20636 20692 20692 22092
rect 20860 20914 20916 22988
rect 20972 21028 21028 23212
rect 20972 20962 21028 20972
rect 20860 20862 20862 20914
rect 20914 20862 20916 20914
rect 20860 20850 20916 20862
rect 20636 20636 20916 20692
rect 20524 20132 20692 20188
rect 20524 20020 20580 20030
rect 20524 19458 20580 19964
rect 20524 19406 20526 19458
rect 20578 19406 20580 19458
rect 20524 19394 20580 19406
rect 20412 19058 20468 19068
rect 18956 14924 19572 14980
rect 19628 16994 20132 16996
rect 19628 16942 20078 16994
rect 20130 16942 20132 16994
rect 19628 16940 20132 16942
rect 18956 14530 19012 14924
rect 18956 14478 18958 14530
rect 19010 14478 19012 14530
rect 18956 14466 19012 14478
rect 19068 14532 19124 14542
rect 18732 13746 18900 13748
rect 18732 13694 18734 13746
rect 18786 13694 18900 13746
rect 18732 13692 18900 13694
rect 18956 13748 19012 13758
rect 19068 13748 19124 14476
rect 19292 14420 19348 14430
rect 19180 14306 19236 14318
rect 19180 14254 19182 14306
rect 19234 14254 19236 14306
rect 19180 13860 19236 14254
rect 19292 13972 19348 14364
rect 19516 14420 19572 14430
rect 19404 14308 19460 14318
rect 19404 14214 19460 14252
rect 19516 14084 19572 14364
rect 19292 13878 19348 13916
rect 19404 14028 19572 14084
rect 19180 13794 19236 13804
rect 18956 13746 19124 13748
rect 18956 13694 18958 13746
rect 19010 13694 19124 13746
rect 18956 13692 19124 13694
rect 18732 13524 18788 13692
rect 18732 13458 18788 13468
rect 18956 13300 19012 13692
rect 17948 13134 17950 13186
rect 18002 13134 18004 13186
rect 17948 13122 18004 13134
rect 18060 13244 18396 13300
rect 18060 12850 18116 13244
rect 18396 13234 18452 13244
rect 18508 13244 19012 13300
rect 18284 12964 18340 12974
rect 18508 12964 18564 13244
rect 19068 13188 19124 13198
rect 19404 13188 19460 14028
rect 19628 13748 19684 16940
rect 20076 16930 20132 16940
rect 20188 18452 20244 18462
rect 20188 16548 20244 18396
rect 20524 18452 20580 18462
rect 20636 18452 20692 20132
rect 20524 18450 20692 18452
rect 20524 18398 20526 18450
rect 20578 18398 20692 18450
rect 20524 18396 20692 18398
rect 20748 19010 20804 19022
rect 20748 18958 20750 19010
rect 20802 18958 20804 19010
rect 20748 18900 20804 18958
rect 20524 18004 20580 18396
rect 20748 18340 20804 18844
rect 20860 18564 20916 20636
rect 20972 20132 21028 20142
rect 20972 20038 21028 20076
rect 21196 19236 21252 23548
rect 21308 23492 21364 23502
rect 21308 23378 21364 23436
rect 21308 23326 21310 23378
rect 21362 23326 21364 23378
rect 21308 23314 21364 23326
rect 21644 23380 21700 23662
rect 21868 23716 21924 24558
rect 21868 23650 21924 23660
rect 21980 23940 22036 25228
rect 21644 23314 21700 23324
rect 21532 23266 21588 23278
rect 21532 23214 21534 23266
rect 21586 23214 21588 23266
rect 21532 23156 21588 23214
rect 21532 23090 21588 23100
rect 21644 23156 21700 23166
rect 21644 23154 21812 23156
rect 21644 23102 21646 23154
rect 21698 23102 21812 23154
rect 21644 23100 21812 23102
rect 21644 23090 21700 23100
rect 21372 22764 21636 22774
rect 21428 22708 21476 22764
rect 21532 22708 21580 22764
rect 21372 22698 21636 22708
rect 21420 22260 21476 22270
rect 21644 22260 21700 22270
rect 21476 22204 21588 22260
rect 21420 22194 21476 22204
rect 21308 22148 21364 22158
rect 21308 22054 21364 22092
rect 21532 22146 21588 22204
rect 21644 22166 21700 22204
rect 21532 22094 21534 22146
rect 21586 22094 21588 22146
rect 21532 22082 21588 22094
rect 21644 21700 21700 21710
rect 21644 21474 21700 21644
rect 21644 21422 21646 21474
rect 21698 21422 21700 21474
rect 21644 21410 21700 21422
rect 21372 21196 21636 21206
rect 21428 21140 21476 21196
rect 21532 21140 21580 21196
rect 21372 21130 21636 21140
rect 21756 21140 21812 23100
rect 21868 22820 21924 22830
rect 21868 21476 21924 22764
rect 21980 22370 22036 23884
rect 22092 23716 22148 23726
rect 22092 23622 22148 23660
rect 21980 22318 21982 22370
rect 22034 22318 22036 22370
rect 21980 21588 22036 22318
rect 21980 21522 22036 21532
rect 21868 21410 21924 21420
rect 21756 21074 21812 21084
rect 21868 21252 21924 21262
rect 21420 20802 21476 20814
rect 21420 20750 21422 20802
rect 21474 20750 21476 20802
rect 21420 20244 21476 20750
rect 21420 20178 21476 20188
rect 21756 20020 21812 20030
rect 21868 20020 21924 21196
rect 22092 20690 22148 20702
rect 22092 20638 22094 20690
rect 22146 20638 22148 20690
rect 21812 19964 21924 20020
rect 21980 20020 22036 20030
rect 21756 19954 21812 19964
rect 21532 19906 21588 19918
rect 21532 19854 21534 19906
rect 21586 19854 21588 19906
rect 21532 19796 21588 19854
rect 21532 19730 21588 19740
rect 21980 19906 22036 19964
rect 21980 19854 21982 19906
rect 22034 19854 22036 19906
rect 21980 19796 22036 19854
rect 21980 19730 22036 19740
rect 21372 19628 21636 19638
rect 21428 19572 21476 19628
rect 21532 19572 21580 19628
rect 21372 19562 21636 19572
rect 21868 19460 21924 19470
rect 21868 19346 21924 19404
rect 22092 19458 22148 20638
rect 22204 20132 22260 25676
rect 22316 23378 22372 25788
rect 22652 24612 22708 24622
rect 22428 24052 22484 24062
rect 22428 23826 22484 23996
rect 22428 23774 22430 23826
rect 22482 23774 22484 23826
rect 22428 23762 22484 23774
rect 22316 23326 22318 23378
rect 22370 23326 22372 23378
rect 22316 21700 22372 23326
rect 22652 23266 22708 24556
rect 23100 24162 23156 26348
rect 23436 26180 23492 27132
rect 23436 26114 23492 26124
rect 23100 24110 23102 24162
rect 23154 24110 23156 24162
rect 23100 24098 23156 24110
rect 23436 23940 23492 23950
rect 23436 23846 23492 23884
rect 22876 23828 22932 23838
rect 22876 23734 22932 23772
rect 22988 23714 23044 23726
rect 22988 23662 22990 23714
rect 23042 23662 23044 23714
rect 22988 23492 23044 23662
rect 23548 23604 23604 29260
rect 23884 29250 23940 29260
rect 23996 28868 24052 34200
rect 24556 31332 24612 31342
rect 24556 31218 24612 31276
rect 24556 31166 24558 31218
rect 24610 31166 24612 31218
rect 24556 31154 24612 31166
rect 24892 31108 24948 31118
rect 24892 31014 24948 31052
rect 24332 30212 24388 30222
rect 24332 29988 24388 30156
rect 24332 29894 24388 29932
rect 24892 30210 24948 30222
rect 24892 30158 24894 30210
rect 24946 30158 24948 30210
rect 24108 29652 24164 29662
rect 24108 29426 24164 29596
rect 24668 29652 24724 29662
rect 24108 29374 24110 29426
rect 24162 29374 24164 29426
rect 24108 29362 24164 29374
rect 24444 29428 24500 29438
rect 24444 29426 24612 29428
rect 24444 29374 24446 29426
rect 24498 29374 24612 29426
rect 24444 29372 24612 29374
rect 24444 29362 24500 29372
rect 23996 28802 24052 28812
rect 24556 28644 24612 29372
rect 24332 28308 24388 28318
rect 24332 28082 24388 28252
rect 24332 28030 24334 28082
rect 24386 28030 24388 28082
rect 24332 28018 24388 28030
rect 24556 28082 24612 28588
rect 24556 28030 24558 28082
rect 24610 28030 24612 28082
rect 24556 28018 24612 28030
rect 24668 28756 24724 29596
rect 24668 27970 24724 28700
rect 24668 27918 24670 27970
rect 24722 27918 24724 27970
rect 24668 27906 24724 27918
rect 24780 29316 24836 29326
rect 23996 27860 24052 27870
rect 23996 27746 24052 27804
rect 23996 27694 23998 27746
rect 24050 27694 24052 27746
rect 23996 27682 24052 27694
rect 24108 27074 24164 27086
rect 24108 27022 24110 27074
rect 24162 27022 24164 27074
rect 24108 26964 24164 27022
rect 24780 26908 24836 29260
rect 24892 29204 24948 30158
rect 24892 29138 24948 29148
rect 25116 27524 25172 34200
rect 26236 31444 26292 34200
rect 25404 31388 25668 31398
rect 26236 31388 26852 31444
rect 25460 31332 25508 31388
rect 25564 31332 25612 31388
rect 25404 31322 25668 31332
rect 26236 31220 26292 31230
rect 26236 31126 26292 31164
rect 25228 31108 25284 31118
rect 25228 30772 25284 31052
rect 25228 29428 25284 30716
rect 25340 30994 25396 31006
rect 25340 30942 25342 30994
rect 25394 30942 25396 30994
rect 25340 30212 25396 30942
rect 25340 30146 25396 30156
rect 26572 30212 26628 30222
rect 25564 30100 25620 30110
rect 25564 30006 25620 30044
rect 25404 29820 25668 29830
rect 25460 29764 25508 29820
rect 25564 29764 25612 29820
rect 25404 29754 25668 29764
rect 25452 29428 25508 29438
rect 26124 29428 26180 29438
rect 25228 29426 25844 29428
rect 25228 29374 25454 29426
rect 25506 29374 25844 29426
rect 25228 29372 25844 29374
rect 25452 29362 25508 29372
rect 25228 29204 25284 29214
rect 25228 28084 25284 29148
rect 25676 29202 25732 29214
rect 25676 29150 25678 29202
rect 25730 29150 25732 29202
rect 25564 28756 25620 28766
rect 25564 28662 25620 28700
rect 25676 28420 25732 29150
rect 25676 28354 25732 28364
rect 25788 28308 25844 29372
rect 26124 29426 26404 29428
rect 26124 29374 26126 29426
rect 26178 29374 26404 29426
rect 26124 29372 26404 29374
rect 26124 29362 26180 29372
rect 26124 29202 26180 29214
rect 26124 29150 26126 29202
rect 26178 29150 26180 29202
rect 26124 28756 26180 29150
rect 26012 28700 26180 28756
rect 26236 29202 26292 29214
rect 26236 29150 26238 29202
rect 26290 29150 26292 29202
rect 25404 28252 25668 28262
rect 25460 28196 25508 28252
rect 25564 28196 25612 28252
rect 25788 28242 25844 28252
rect 25900 28642 25956 28654
rect 25900 28590 25902 28642
rect 25954 28590 25956 28642
rect 25404 28186 25668 28196
rect 25788 28084 25844 28094
rect 25228 28028 25396 28084
rect 25116 27458 25172 27468
rect 25228 27746 25284 27758
rect 25228 27694 25230 27746
rect 25282 27694 25284 27746
rect 24108 26898 24164 26908
rect 24556 26852 24836 26908
rect 25004 27412 25060 27422
rect 23996 26292 24052 26302
rect 23996 25396 24052 26236
rect 24444 26178 24500 26190
rect 24444 26126 24446 26178
rect 24498 26126 24500 26178
rect 24444 25620 24500 26126
rect 24444 25554 24500 25564
rect 23996 24610 24052 25340
rect 24332 24724 24388 24734
rect 23996 24558 23998 24610
rect 24050 24558 24052 24610
rect 23996 24546 24052 24558
rect 24108 24722 24388 24724
rect 24108 24670 24334 24722
rect 24386 24670 24388 24722
rect 24108 24668 24388 24670
rect 22652 23214 22654 23266
rect 22706 23214 22708 23266
rect 22652 23202 22708 23214
rect 22764 23436 23044 23492
rect 23100 23548 23604 23604
rect 22540 23156 22596 23194
rect 22540 23090 22596 23100
rect 22764 22484 22820 23436
rect 22988 23266 23044 23278
rect 22988 23214 22990 23266
rect 23042 23214 23044 23266
rect 22988 22820 23044 23214
rect 22988 22754 23044 22764
rect 22316 21634 22372 21644
rect 22428 22428 22820 22484
rect 22316 21474 22372 21486
rect 22316 21422 22318 21474
rect 22370 21422 22372 21474
rect 22316 21252 22372 21422
rect 22316 21186 22372 21196
rect 22428 20356 22484 22428
rect 22764 22258 22820 22270
rect 22764 22206 22766 22258
rect 22818 22206 22820 22258
rect 22764 21812 22820 22206
rect 22764 21746 22820 21756
rect 22876 21698 22932 21710
rect 22876 21646 22878 21698
rect 22930 21646 22932 21698
rect 22764 21588 22820 21598
rect 22204 20066 22260 20076
rect 22316 20300 22484 20356
rect 22540 21476 22596 21486
rect 22092 19406 22094 19458
rect 22146 19406 22148 19458
rect 22092 19394 22148 19406
rect 21868 19294 21870 19346
rect 21922 19294 21924 19346
rect 21196 19180 21812 19236
rect 21532 19010 21588 19022
rect 21532 18958 21534 19010
rect 21586 18958 21588 19010
rect 21532 18676 21588 18958
rect 20860 18498 20916 18508
rect 20972 18620 21588 18676
rect 20748 18274 20804 18284
rect 20972 18338 21028 18620
rect 21308 18452 21364 18462
rect 20972 18286 20974 18338
rect 21026 18286 21028 18338
rect 20972 18116 21028 18286
rect 20524 17938 20580 17948
rect 20636 18060 21028 18116
rect 21084 18450 21364 18452
rect 21084 18398 21310 18450
rect 21362 18398 21364 18450
rect 21084 18396 21364 18398
rect 20636 17780 20692 18060
rect 21084 18004 21140 18396
rect 21308 18386 21364 18396
rect 21532 18450 21588 18462
rect 21532 18398 21534 18450
rect 21586 18398 21588 18450
rect 21532 18228 21588 18398
rect 21644 18452 21700 18462
rect 21644 18358 21700 18396
rect 21756 18340 21812 19180
rect 21868 18788 21924 19294
rect 22316 19236 22372 20300
rect 22428 20130 22484 20142
rect 22428 20078 22430 20130
rect 22482 20078 22484 20130
rect 22428 20020 22484 20078
rect 22540 20130 22596 21420
rect 22652 21362 22708 21374
rect 22652 21310 22654 21362
rect 22706 21310 22708 21362
rect 22652 20916 22708 21310
rect 22652 20580 22708 20860
rect 22652 20514 22708 20524
rect 22540 20078 22542 20130
rect 22594 20078 22596 20130
rect 22540 20066 22596 20078
rect 22428 19954 22484 19964
rect 22428 19796 22484 19806
rect 22764 19796 22820 21532
rect 22876 21252 22932 21646
rect 22876 21186 22932 21196
rect 22988 21362 23044 21374
rect 22988 21310 22990 21362
rect 23042 21310 23044 21362
rect 22988 21028 23044 21310
rect 22988 20962 23044 20972
rect 23100 20188 23156 23548
rect 23884 23492 23940 23502
rect 23324 23156 23380 23166
rect 23324 23154 23604 23156
rect 23324 23102 23326 23154
rect 23378 23102 23604 23154
rect 23324 23100 23604 23102
rect 23324 23090 23380 23100
rect 23436 22932 23492 22942
rect 23212 22148 23268 22158
rect 23212 21586 23268 22092
rect 23212 21534 23214 21586
rect 23266 21534 23268 21586
rect 23212 21522 23268 21534
rect 22876 20132 22932 20142
rect 23100 20132 23268 20188
rect 22876 20038 22932 20076
rect 23100 20018 23156 20030
rect 23100 19966 23102 20018
rect 23154 19966 23156 20018
rect 22428 19794 22820 19796
rect 22428 19742 22430 19794
rect 22482 19742 22820 19794
rect 22428 19740 22820 19742
rect 22988 19906 23044 19918
rect 22988 19854 22990 19906
rect 23042 19854 23044 19906
rect 22428 19730 22484 19740
rect 22876 19460 22932 19470
rect 22988 19460 23044 19854
rect 22876 19458 23044 19460
rect 22876 19406 22878 19458
rect 22930 19406 23044 19458
rect 22876 19404 23044 19406
rect 23100 19460 23156 19966
rect 22876 19394 22932 19404
rect 23100 19394 23156 19404
rect 22988 19236 23044 19246
rect 23212 19236 23268 20132
rect 23436 19348 23492 22876
rect 23548 21364 23604 23100
rect 23884 23154 23940 23436
rect 23884 23102 23886 23154
rect 23938 23102 23940 23154
rect 23884 22596 23940 23102
rect 23884 22530 23940 22540
rect 23884 22148 23940 22158
rect 23772 21812 23828 21822
rect 23772 21718 23828 21756
rect 23884 21810 23940 22092
rect 23884 21758 23886 21810
rect 23938 21758 23940 21810
rect 23884 21746 23940 21758
rect 23660 21588 23716 21598
rect 23660 21494 23716 21532
rect 23548 21308 23828 21364
rect 23548 20020 23604 20030
rect 23548 20018 23716 20020
rect 23548 19966 23550 20018
rect 23602 19966 23716 20018
rect 23548 19964 23716 19966
rect 23548 19954 23604 19964
rect 23660 19460 23716 19964
rect 23772 20018 23828 21308
rect 23772 19966 23774 20018
rect 23826 19966 23828 20018
rect 23772 19908 23828 19966
rect 23772 19842 23828 19852
rect 23884 20132 23940 20142
rect 23772 19460 23828 19470
rect 23660 19458 23828 19460
rect 23660 19406 23774 19458
rect 23826 19406 23828 19458
rect 23660 19404 23828 19406
rect 23772 19394 23828 19404
rect 23436 19292 23716 19348
rect 22316 19180 22484 19236
rect 21868 18722 21924 18732
rect 22316 19010 22372 19022
rect 22316 18958 22318 19010
rect 22370 18958 22372 19010
rect 22316 18900 22372 18958
rect 22316 18564 22372 18844
rect 22316 18498 22372 18508
rect 22092 18452 22148 18462
rect 22092 18358 22148 18396
rect 21756 18284 21924 18340
rect 20748 17948 21140 18004
rect 21196 18172 21588 18228
rect 21868 18228 21924 18284
rect 20748 17890 20804 17948
rect 20748 17838 20750 17890
rect 20802 17838 20804 17890
rect 20748 17826 20804 17838
rect 20188 16482 20244 16492
rect 20300 17668 20356 17678
rect 20188 16098 20244 16110
rect 20188 16046 20190 16098
rect 20242 16046 20244 16098
rect 19740 15876 19796 15886
rect 19740 15782 19796 15820
rect 19852 15874 19908 15886
rect 19852 15822 19854 15874
rect 19906 15822 19908 15874
rect 19740 15090 19796 15102
rect 19740 15038 19742 15090
rect 19794 15038 19796 15090
rect 19740 14980 19796 15038
rect 19852 15092 19908 15822
rect 19964 15874 20020 15886
rect 19964 15822 19966 15874
rect 20018 15822 20020 15874
rect 19964 15428 20020 15822
rect 19964 15362 20020 15372
rect 20076 15764 20132 15774
rect 20076 15314 20132 15708
rect 20188 15652 20244 16046
rect 20188 15586 20244 15596
rect 20076 15262 20078 15314
rect 20130 15262 20132 15314
rect 20076 15250 20132 15262
rect 20300 15314 20356 17612
rect 20636 17554 20692 17724
rect 21196 17668 21252 18172
rect 21868 18162 21924 18172
rect 21372 18060 21636 18070
rect 21428 18004 21476 18060
rect 21532 18004 21580 18060
rect 21372 17994 21636 18004
rect 21980 18004 22036 18014
rect 21980 17780 22036 17948
rect 20636 17502 20638 17554
rect 20690 17502 20692 17554
rect 20524 17444 20580 17454
rect 20300 15262 20302 15314
rect 20354 15262 20356 15314
rect 20300 15250 20356 15262
rect 20412 16772 20468 16782
rect 20412 15316 20468 16716
rect 20524 16098 20580 17388
rect 20636 16996 20692 17502
rect 20636 16930 20692 16940
rect 20748 17612 21252 17668
rect 21308 17668 21364 17678
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 20524 16034 20580 16046
rect 20748 15764 20804 17612
rect 21308 17556 21364 17612
rect 21196 17554 21364 17556
rect 21196 17502 21310 17554
rect 21362 17502 21364 17554
rect 21196 17500 21364 17502
rect 21084 17220 21140 17230
rect 21084 15876 21140 17164
rect 21196 16100 21252 17500
rect 21308 17490 21364 17500
rect 21644 17554 21700 17566
rect 21644 17502 21646 17554
rect 21698 17502 21700 17554
rect 21644 16996 21700 17502
rect 21980 17332 22036 17724
rect 22204 17780 22260 17790
rect 22204 17444 22260 17724
rect 22204 17378 22260 17388
rect 21980 17266 22036 17276
rect 21644 16930 21700 16940
rect 21372 16492 21636 16502
rect 21428 16436 21476 16492
rect 21532 16436 21580 16492
rect 21372 16426 21636 16436
rect 22204 16212 22260 16222
rect 22204 16210 22372 16212
rect 22204 16158 22206 16210
rect 22258 16158 22372 16210
rect 22204 16156 22372 16158
rect 22204 16146 22260 16156
rect 21308 16100 21364 16110
rect 21196 16098 21364 16100
rect 21196 16046 21310 16098
rect 21362 16046 21364 16098
rect 21196 16044 21364 16046
rect 21308 16034 21364 16044
rect 21532 15988 21588 15998
rect 21532 15894 21588 15932
rect 21644 15986 21700 15998
rect 21644 15934 21646 15986
rect 21698 15934 21700 15986
rect 21644 15876 21700 15934
rect 21084 15820 21364 15876
rect 20636 15708 20804 15764
rect 20524 15428 20580 15438
rect 20524 15334 20580 15372
rect 20412 15250 20468 15260
rect 19852 15036 20020 15092
rect 19740 14924 19908 14980
rect 19068 13186 19460 13188
rect 19068 13134 19070 13186
rect 19122 13134 19460 13186
rect 19068 13132 19460 13134
rect 19516 13692 19684 13748
rect 19740 14756 19796 14766
rect 19068 13122 19124 13132
rect 18732 13074 18788 13086
rect 18732 13022 18734 13074
rect 18786 13022 18788 13074
rect 18284 12962 18564 12964
rect 18284 12910 18286 12962
rect 18338 12910 18564 12962
rect 18284 12908 18564 12910
rect 18620 12964 18676 12974
rect 18732 12964 18788 13022
rect 18620 12962 18788 12964
rect 18620 12910 18622 12962
rect 18674 12910 18788 12962
rect 18620 12908 18788 12910
rect 19068 12964 19124 12974
rect 18284 12898 18340 12908
rect 18620 12898 18676 12908
rect 19068 12870 19124 12908
rect 19516 12852 19572 13692
rect 19628 13524 19684 13534
rect 19740 13524 19796 14700
rect 19852 14420 19908 14924
rect 19852 14354 19908 14364
rect 19628 13522 19796 13524
rect 19628 13470 19630 13522
rect 19682 13470 19796 13522
rect 19628 13468 19796 13470
rect 19852 13634 19908 13646
rect 19852 13582 19854 13634
rect 19906 13582 19908 13634
rect 19852 13524 19908 13582
rect 19964 13636 20020 15036
rect 20076 14532 20132 14542
rect 20076 14438 20132 14476
rect 20524 14532 20580 14542
rect 20524 14438 20580 14476
rect 20636 14308 20692 15708
rect 21196 15540 21252 15550
rect 21196 15446 21252 15484
rect 20636 14214 20692 14252
rect 20748 15426 20804 15438
rect 20748 15374 20750 15426
rect 20802 15374 20804 15426
rect 20188 13972 20244 13982
rect 20188 13914 20244 13916
rect 20188 13862 20190 13914
rect 20242 13862 20244 13914
rect 20412 13972 20468 13982
rect 20188 13850 20244 13862
rect 20300 13860 20356 13870
rect 20412 13860 20468 13916
rect 20300 13858 20468 13860
rect 20300 13806 20302 13858
rect 20354 13806 20468 13858
rect 20300 13804 20468 13806
rect 20300 13636 20356 13804
rect 20524 13748 20580 13758
rect 20524 13654 20580 13692
rect 19964 13580 20132 13636
rect 20076 13524 20132 13580
rect 20300 13570 20356 13580
rect 20636 13636 20692 13646
rect 20748 13636 20804 15374
rect 21308 15426 21364 15820
rect 21644 15810 21700 15820
rect 22316 15540 22372 16156
rect 22092 15484 22372 15540
rect 21308 15374 21310 15426
rect 21362 15374 21364 15426
rect 20860 15314 20916 15326
rect 20860 15262 20862 15314
rect 20914 15262 20916 15314
rect 20860 14420 20916 15262
rect 21308 15092 21364 15374
rect 21644 15428 21700 15438
rect 21644 15334 21700 15372
rect 21980 15316 22036 15326
rect 21980 15222 22036 15260
rect 21308 15026 21364 15036
rect 21980 15092 22036 15102
rect 21372 14924 21636 14934
rect 21428 14868 21476 14924
rect 21532 14868 21580 14924
rect 21372 14858 21636 14868
rect 21196 14532 21252 14542
rect 21084 14420 21140 14430
rect 20860 14364 21084 14420
rect 21084 13858 21140 14364
rect 21084 13806 21086 13858
rect 21138 13806 21140 13858
rect 21084 13794 21140 13806
rect 20748 13580 21140 13636
rect 20076 13468 20244 13524
rect 19628 13458 19684 13468
rect 19852 13458 19908 13468
rect 18060 12798 18062 12850
rect 18114 12798 18116 12850
rect 18060 12786 18116 12798
rect 19180 12796 19572 12852
rect 19628 13188 19684 13198
rect 20076 13188 20132 13198
rect 17836 11454 17838 11506
rect 17890 11454 17892 11506
rect 17836 11442 17892 11454
rect 17052 11396 17108 11406
rect 17052 11302 17108 11340
rect 14812 11172 14868 11182
rect 14700 11170 14868 11172
rect 14700 11118 14814 11170
rect 14866 11118 14868 11170
rect 14700 11116 14868 11118
rect 13916 9940 13972 9950
rect 13916 9846 13972 9884
rect 13132 9762 13188 9772
rect 13804 9716 13860 9726
rect 13804 9622 13860 9660
rect 12908 9436 13188 9492
rect 12460 9212 12740 9268
rect 11788 6748 11956 6804
rect 10780 5966 10782 6018
rect 10834 5966 10836 6018
rect 10444 5954 10500 5964
rect 10780 5954 10836 5966
rect 11004 6692 11060 6702
rect 11004 6018 11060 6636
rect 11340 6692 11396 6702
rect 11340 6598 11396 6636
rect 11900 6690 11956 6748
rect 11900 6638 11902 6690
rect 11954 6638 11956 6690
rect 11116 6578 11172 6590
rect 11116 6526 11118 6578
rect 11170 6526 11172 6578
rect 11116 6356 11172 6526
rect 11788 6580 11844 6590
rect 11564 6466 11620 6478
rect 11564 6414 11566 6466
rect 11618 6414 11620 6466
rect 11564 6356 11620 6414
rect 11116 6300 11620 6356
rect 11004 5966 11006 6018
rect 11058 5966 11060 6018
rect 11004 5954 11060 5966
rect 11788 5906 11844 6524
rect 11900 6356 11956 6638
rect 11900 6290 11956 6300
rect 11788 5854 11790 5906
rect 11842 5854 11844 5906
rect 11788 5842 11844 5854
rect 11900 6020 11956 6030
rect 10556 5794 10612 5806
rect 10556 5742 10558 5794
rect 10610 5742 10612 5794
rect 10556 5236 10612 5742
rect 10556 5170 10612 5180
rect 11900 5234 11956 5964
rect 11900 5182 11902 5234
rect 11954 5182 11956 5234
rect 11900 5170 11956 5182
rect 11676 5124 11732 5134
rect 9548 3666 9940 3668
rect 9548 3614 9550 3666
rect 9602 3614 9940 3666
rect 9548 3612 9940 3614
rect 10332 4226 10388 4238
rect 10332 4174 10334 4226
rect 10386 4174 10388 4226
rect 9548 3602 9604 3612
rect 8540 3332 8820 3388
rect 5852 3322 5908 3332
rect 6076 3276 6244 3332
rect 7196 800 7252 3332
rect 8764 800 8820 3332
rect 9276 3164 9540 3174
rect 9332 3108 9380 3164
rect 9436 3108 9484 3164
rect 9276 3098 9540 3108
rect 10332 800 10388 4174
rect 11676 3666 11732 5068
rect 12012 4338 12068 8428
rect 12124 9042 12180 9054
rect 12124 8990 12126 9042
rect 12178 8990 12180 9042
rect 12124 7364 12180 8990
rect 12236 7476 12292 9100
rect 12348 9154 12404 9166
rect 12348 9102 12350 9154
rect 12402 9102 12404 9154
rect 12348 7700 12404 9102
rect 12460 9042 12516 9054
rect 12460 8990 12462 9042
rect 12514 8990 12516 9042
rect 12460 8932 12516 8990
rect 12460 8866 12516 8876
rect 12572 9044 12628 9054
rect 12348 7634 12404 7644
rect 12460 8260 12516 8270
rect 12348 7476 12404 7486
rect 12236 7474 12404 7476
rect 12236 7422 12350 7474
rect 12402 7422 12404 7474
rect 12236 7420 12404 7422
rect 12124 7298 12180 7308
rect 12124 6916 12180 6926
rect 12180 6860 12292 6916
rect 12124 6850 12180 6860
rect 12236 6244 12292 6860
rect 12348 6692 12404 7420
rect 12348 6626 12404 6636
rect 12460 6690 12516 8204
rect 12572 8258 12628 8988
rect 12572 8206 12574 8258
rect 12626 8206 12628 8258
rect 12572 8194 12628 8206
rect 12684 7812 12740 9212
rect 12908 9044 12964 9436
rect 13132 9266 13188 9436
rect 13132 9214 13134 9266
rect 13186 9214 13188 9266
rect 13132 9202 13188 9214
rect 12908 8978 12964 8988
rect 13692 9156 13748 9166
rect 13692 9042 13748 9100
rect 13692 8990 13694 9042
rect 13746 8990 13748 9042
rect 13692 8978 13748 8990
rect 13308 8652 13572 8662
rect 13364 8596 13412 8652
rect 13468 8596 13516 8652
rect 13308 8586 13572 8596
rect 12908 8036 12964 8046
rect 12908 8034 13412 8036
rect 12908 7982 12910 8034
rect 12962 7982 13412 8034
rect 12908 7980 13412 7982
rect 12908 7970 12964 7980
rect 12572 7756 12740 7812
rect 12572 6804 12628 7756
rect 13244 7700 13300 7710
rect 12572 6738 12628 6748
rect 12684 7698 13300 7700
rect 12684 7646 13246 7698
rect 13298 7646 13300 7698
rect 12684 7644 13300 7646
rect 12460 6638 12462 6690
rect 12514 6638 12516 6690
rect 12460 6626 12516 6638
rect 12572 6468 12628 6478
rect 12572 6374 12628 6412
rect 12236 6188 12628 6244
rect 12124 5684 12180 5694
rect 12348 5684 12404 5694
rect 12124 5122 12180 5628
rect 12124 5070 12126 5122
rect 12178 5070 12180 5122
rect 12124 5058 12180 5070
rect 12236 5682 12404 5684
rect 12236 5630 12350 5682
rect 12402 5630 12404 5682
rect 12236 5628 12404 5630
rect 12012 4286 12014 4338
rect 12066 4286 12068 4338
rect 12012 4274 12068 4286
rect 11676 3614 11678 3666
rect 11730 3614 11732 3666
rect 11676 3602 11732 3614
rect 12236 3388 12292 5628
rect 12348 5618 12404 5628
rect 12460 5684 12516 5694
rect 12348 5124 12404 5134
rect 12348 5030 12404 5068
rect 12460 3554 12516 5628
rect 12572 5122 12628 6188
rect 12572 5070 12574 5122
rect 12626 5070 12628 5122
rect 12572 5058 12628 5070
rect 12460 3502 12462 3554
rect 12514 3502 12516 3554
rect 12460 3490 12516 3502
rect 12684 4226 12740 7644
rect 13244 7634 13300 7644
rect 13132 7476 13188 7486
rect 13356 7476 13412 7980
rect 12908 7474 13412 7476
rect 12908 7422 13134 7474
rect 13186 7422 13412 7474
rect 12908 7420 13412 7422
rect 12908 6690 12964 7420
rect 13132 7410 13188 7420
rect 13356 7364 13412 7420
rect 13356 7298 13412 7308
rect 13692 7700 13748 7710
rect 13692 7474 13748 7644
rect 13692 7422 13694 7474
rect 13746 7422 13748 7474
rect 13244 7252 13300 7262
rect 13132 7250 13300 7252
rect 13132 7198 13246 7250
rect 13298 7198 13300 7250
rect 13132 7196 13300 7198
rect 12908 6638 12910 6690
rect 12962 6638 12964 6690
rect 12908 6626 12964 6638
rect 13020 6804 13076 6814
rect 12796 6580 12852 6590
rect 12796 6244 12852 6524
rect 12796 6178 12852 6188
rect 12796 5124 12852 5134
rect 13020 5124 13076 6748
rect 13132 6020 13188 7196
rect 13244 7186 13300 7196
rect 13308 7084 13572 7094
rect 13364 7028 13412 7084
rect 13468 7028 13516 7084
rect 13308 7018 13572 7028
rect 13692 6916 13748 7422
rect 13356 6860 13748 6916
rect 13244 6132 13300 6142
rect 13356 6132 13412 6860
rect 13300 6076 13412 6132
rect 13580 6692 13636 6702
rect 13244 6066 13300 6076
rect 13132 5954 13188 5964
rect 13580 5684 13636 6636
rect 14028 6580 14084 11116
rect 14252 11106 14308 11116
rect 14140 10612 14196 10622
rect 14140 9826 14196 10556
rect 14140 9774 14142 9826
rect 14194 9774 14196 9826
rect 14140 9762 14196 9774
rect 14252 10500 14308 10510
rect 14812 10500 14868 11116
rect 17340 11004 17604 11014
rect 17396 10948 17444 11004
rect 17500 10948 17548 11004
rect 17340 10938 17604 10948
rect 15596 10610 15652 10622
rect 15596 10558 15598 10610
rect 15650 10558 15652 10610
rect 15148 10500 15204 10510
rect 14252 9156 14308 10444
rect 14588 10444 14868 10500
rect 15036 10498 15204 10500
rect 15036 10446 15150 10498
rect 15202 10446 15204 10498
rect 15036 10444 15204 10446
rect 14364 10164 14420 10174
rect 14364 9826 14420 10108
rect 14364 9774 14366 9826
rect 14418 9774 14420 9826
rect 14364 9762 14420 9774
rect 14476 9156 14532 9166
rect 14252 9154 14532 9156
rect 14252 9102 14478 9154
rect 14530 9102 14532 9154
rect 14252 9100 14532 9102
rect 14476 9090 14532 9100
rect 13580 5618 13636 5628
rect 13692 6356 13748 6366
rect 13308 5516 13572 5526
rect 13364 5460 13412 5516
rect 13468 5460 13516 5516
rect 13308 5450 13572 5460
rect 13692 5348 13748 6300
rect 13580 5292 13748 5348
rect 13580 5124 13636 5292
rect 12796 5122 13076 5124
rect 12796 5070 12798 5122
rect 12850 5070 13076 5122
rect 12796 5068 13076 5070
rect 13132 5068 13636 5124
rect 12796 5058 12852 5068
rect 12684 4174 12686 4226
rect 12738 4174 12740 4226
rect 11900 3332 12292 3388
rect 12684 3444 12740 4174
rect 13132 3556 13188 5068
rect 13580 5010 13636 5068
rect 13916 5124 13972 5134
rect 14028 5124 14084 6524
rect 14364 6578 14420 6590
rect 14364 6526 14366 6578
rect 14418 6526 14420 6578
rect 13916 5122 14084 5124
rect 13916 5070 13918 5122
rect 13970 5070 14084 5122
rect 13916 5068 14084 5070
rect 14140 6468 14196 6478
rect 14140 5122 14196 6412
rect 14252 6244 14308 6254
rect 14252 5906 14308 6188
rect 14252 5854 14254 5906
rect 14306 5854 14308 5906
rect 14252 5842 14308 5854
rect 14364 5908 14420 6526
rect 14364 5842 14420 5852
rect 14476 5124 14532 5134
rect 14140 5070 14142 5122
rect 14194 5070 14196 5122
rect 13916 5058 13972 5068
rect 14140 5058 14196 5070
rect 14252 5122 14532 5124
rect 14252 5070 14478 5122
rect 14530 5070 14532 5122
rect 14252 5068 14532 5070
rect 13580 4958 13582 5010
rect 13634 4958 13636 5010
rect 13580 4946 13636 4958
rect 14252 4004 14308 5068
rect 14476 5058 14532 5068
rect 14588 5124 14644 10444
rect 14812 9604 14868 9614
rect 14812 9510 14868 9548
rect 15036 9602 15092 10444
rect 15148 10434 15204 10444
rect 15148 10164 15204 10174
rect 15148 9938 15204 10108
rect 15148 9886 15150 9938
rect 15202 9886 15204 9938
rect 15148 9874 15204 9886
rect 15596 9940 15652 10558
rect 15708 10612 15764 10622
rect 15708 10518 15764 10556
rect 16156 10610 16212 10622
rect 17276 10612 17332 10622
rect 16156 10558 16158 10610
rect 16210 10558 16212 10610
rect 15932 10500 15988 10510
rect 15932 10406 15988 10444
rect 15708 9940 15764 9950
rect 15596 9938 15764 9940
rect 15596 9886 15710 9938
rect 15762 9886 15764 9938
rect 15596 9884 15764 9886
rect 15708 9874 15764 9884
rect 15036 9550 15038 9602
rect 15090 9550 15092 9602
rect 14924 8260 14980 8270
rect 14924 8166 14980 8204
rect 14924 7362 14980 7374
rect 14924 7310 14926 7362
rect 14978 7310 14980 7362
rect 14588 5058 14644 5068
rect 14812 5236 14868 5246
rect 14812 5122 14868 5180
rect 14812 5070 14814 5122
rect 14866 5070 14868 5122
rect 14812 5058 14868 5070
rect 14476 4898 14532 4910
rect 14476 4846 14478 4898
rect 14530 4846 14532 4898
rect 14476 4564 14532 4846
rect 14476 4508 14868 4564
rect 14812 4450 14868 4508
rect 14812 4398 14814 4450
rect 14866 4398 14868 4450
rect 14812 4386 14868 4398
rect 13308 3948 13572 3958
rect 13364 3892 13412 3948
rect 13468 3892 13516 3948
rect 13308 3882 13572 3892
rect 13692 3948 14308 4004
rect 13244 3556 13300 3566
rect 13132 3554 13300 3556
rect 13132 3502 13246 3554
rect 13298 3502 13300 3554
rect 13132 3500 13300 3502
rect 13244 3490 13300 3500
rect 13580 3556 13636 3566
rect 13692 3556 13748 3948
rect 13580 3554 13748 3556
rect 13580 3502 13582 3554
rect 13634 3502 13748 3554
rect 13580 3500 13748 3502
rect 13804 3554 13860 3566
rect 13804 3502 13806 3554
rect 13858 3502 13860 3554
rect 13580 3490 13636 3500
rect 12684 3378 12740 3388
rect 13356 3444 13412 3482
rect 13356 3378 13412 3388
rect 13804 3444 13860 3502
rect 14924 3388 14980 7310
rect 15036 6692 15092 9550
rect 15260 9604 15316 9614
rect 15596 9604 15652 9614
rect 15260 9602 15596 9604
rect 15260 9550 15262 9602
rect 15314 9550 15596 9602
rect 15260 9548 15596 9550
rect 15260 9538 15316 9548
rect 15596 9510 15652 9548
rect 15820 9602 15876 9614
rect 15820 9550 15822 9602
rect 15874 9550 15876 9602
rect 15820 8932 15876 9550
rect 16156 9156 16212 10558
rect 17164 10610 17332 10612
rect 17164 10558 17278 10610
rect 17330 10558 17332 10610
rect 17164 10556 17332 10558
rect 16268 9826 16324 9838
rect 16268 9774 16270 9826
rect 16322 9774 16324 9826
rect 16268 9268 16324 9774
rect 16604 9828 16660 9838
rect 16604 9826 16772 9828
rect 16604 9774 16606 9826
rect 16658 9774 16772 9826
rect 16604 9772 16772 9774
rect 16604 9762 16660 9772
rect 16268 9202 16324 9212
rect 16156 9090 16212 9100
rect 16716 9044 16772 9772
rect 15820 8866 15876 8876
rect 16604 8932 16660 8942
rect 16604 7700 16660 8876
rect 16716 8484 16772 8988
rect 16716 8418 16772 8428
rect 16828 9156 16884 9166
rect 16604 7634 16660 7644
rect 16492 7588 16548 7598
rect 16492 6802 16548 7532
rect 16716 7588 16772 7598
rect 16716 7494 16772 7532
rect 16492 6750 16494 6802
rect 16546 6750 16548 6802
rect 16492 6738 16548 6750
rect 16604 7474 16660 7486
rect 16604 7422 16606 7474
rect 16658 7422 16660 7474
rect 15036 6626 15092 6636
rect 16604 6580 16660 7422
rect 16828 6804 16884 9100
rect 17164 7700 17220 10556
rect 17276 10546 17332 10556
rect 17612 10612 17668 10622
rect 17612 10518 17668 10556
rect 17836 10610 17892 10622
rect 17836 10558 17838 10610
rect 17890 10558 17892 10610
rect 17500 10498 17556 10510
rect 17500 10446 17502 10498
rect 17554 10446 17556 10498
rect 17500 10052 17556 10446
rect 17276 9996 17556 10052
rect 17276 9938 17332 9996
rect 17276 9886 17278 9938
rect 17330 9886 17332 9938
rect 17276 9874 17332 9886
rect 17340 9436 17604 9446
rect 17396 9380 17444 9436
rect 17500 9380 17548 9436
rect 17340 9370 17604 9380
rect 17500 9268 17556 9278
rect 17500 9174 17556 9212
rect 17836 9266 17892 10558
rect 17836 9214 17838 9266
rect 17890 9214 17892 9266
rect 17836 9202 17892 9214
rect 17948 9828 18004 9838
rect 17948 9604 18004 9772
rect 17948 9266 18004 9548
rect 17948 9214 17950 9266
rect 18002 9214 18004 9266
rect 17948 9202 18004 9214
rect 18172 9716 18228 9726
rect 18172 9266 18228 9660
rect 18172 9214 18174 9266
rect 18226 9214 18228 9266
rect 18172 9202 18228 9214
rect 19068 9268 19124 9278
rect 18396 9154 18452 9166
rect 18396 9102 18398 9154
rect 18450 9102 18452 9154
rect 17724 9044 17780 9054
rect 17724 8950 17780 8988
rect 17836 8484 17892 8494
rect 17836 8146 17892 8428
rect 17836 8094 17838 8146
rect 17890 8094 17892 8146
rect 17340 7868 17604 7878
rect 17396 7812 17444 7868
rect 17500 7812 17548 7868
rect 17340 7802 17604 7812
rect 17500 7700 17556 7710
rect 17164 7698 17556 7700
rect 17164 7646 17502 7698
rect 17554 7646 17556 7698
rect 17164 7644 17556 7646
rect 17500 7634 17556 7644
rect 17612 7700 17668 7710
rect 17612 7606 17668 7644
rect 16940 7474 16996 7486
rect 16940 7422 16942 7474
rect 16994 7422 16996 7474
rect 16940 7252 16996 7422
rect 17388 7476 17444 7486
rect 17388 7364 17444 7420
rect 16940 7186 16996 7196
rect 17164 7308 17444 7364
rect 16940 6804 16996 6814
rect 16828 6802 16996 6804
rect 16828 6750 16942 6802
rect 16994 6750 16996 6802
rect 16828 6748 16996 6750
rect 16940 6738 16996 6748
rect 17052 6692 17108 6702
rect 17052 6598 17108 6636
rect 15260 5684 15316 5694
rect 13804 3378 13860 3388
rect 14252 3332 14980 3388
rect 15036 5682 15316 5684
rect 15036 5630 15262 5682
rect 15314 5630 15316 5682
rect 15036 5628 15316 5630
rect 11900 800 11956 3332
rect 13468 924 13860 980
rect 13468 800 13524 924
rect 896 0 1008 800
rect 2464 0 2576 800
rect 4032 0 4144 800
rect 5600 0 5712 800
rect 7168 0 7280 800
rect 8736 0 8848 800
rect 10304 0 10416 800
rect 11872 0 11984 800
rect 13440 0 13552 800
rect 13804 756 13860 924
rect 14252 756 14308 3332
rect 15036 800 15092 5628
rect 15260 5618 15316 5628
rect 15820 5684 15876 5694
rect 15148 5236 15204 5246
rect 15148 5010 15204 5180
rect 15372 5124 15428 5134
rect 15820 5124 15876 5628
rect 16604 5684 16660 6524
rect 16828 6468 16884 6478
rect 17164 6468 17220 7308
rect 17612 7252 17668 7262
rect 17668 7196 17780 7252
rect 17612 7186 17668 7196
rect 16828 6466 17220 6468
rect 16828 6414 16830 6466
rect 16882 6414 17220 6466
rect 16828 6412 17220 6414
rect 17276 6468 17332 6506
rect 16828 6402 16884 6412
rect 17276 6402 17332 6412
rect 17340 6300 17604 6310
rect 17396 6244 17444 6300
rect 17500 6244 17548 6300
rect 17340 6234 17604 6244
rect 17276 6020 17332 6030
rect 17276 5906 17332 5964
rect 17724 6018 17780 7196
rect 17836 6690 17892 8094
rect 18060 8484 18116 8494
rect 18060 7474 18116 8428
rect 18396 7812 18452 9102
rect 18396 7746 18452 7756
rect 18508 9042 18564 9054
rect 18508 8990 18510 9042
rect 18562 8990 18564 9042
rect 18060 7422 18062 7474
rect 18114 7422 18116 7474
rect 18060 7410 18116 7422
rect 18284 7474 18340 7486
rect 18284 7422 18286 7474
rect 18338 7422 18340 7474
rect 17836 6638 17838 6690
rect 17890 6638 17892 6690
rect 17836 6626 17892 6638
rect 18284 6132 18340 7422
rect 18508 7476 18564 8990
rect 19068 9042 19124 9212
rect 19068 8990 19070 9042
rect 19122 8990 19124 9042
rect 18508 7410 18564 7420
rect 18620 7644 19012 7700
rect 18620 7474 18676 7644
rect 18620 7422 18622 7474
rect 18674 7422 18676 7474
rect 18620 7410 18676 7422
rect 18844 7474 18900 7486
rect 18844 7422 18846 7474
rect 18898 7422 18900 7474
rect 18732 7362 18788 7374
rect 18732 7310 18734 7362
rect 18786 7310 18788 7362
rect 18620 6578 18676 6590
rect 18620 6526 18622 6578
rect 18674 6526 18676 6578
rect 18620 6468 18676 6526
rect 18620 6402 18676 6412
rect 17724 5966 17726 6018
rect 17778 5966 17780 6018
rect 17724 5954 17780 5966
rect 17948 6076 18340 6132
rect 17948 6018 18004 6076
rect 18732 6020 18788 7310
rect 17948 5966 17950 6018
rect 18002 5966 18004 6018
rect 17276 5854 17278 5906
rect 17330 5854 17332 5906
rect 17276 5842 17332 5854
rect 17500 5908 17556 5918
rect 17500 5814 17556 5852
rect 16604 5618 16660 5628
rect 16940 5796 16996 5806
rect 15372 5030 15428 5068
rect 15596 5122 15876 5124
rect 15596 5070 15822 5122
rect 15874 5070 15876 5122
rect 15596 5068 15876 5070
rect 15148 4958 15150 5010
rect 15202 4958 15204 5010
rect 15148 4946 15204 4958
rect 15596 4340 15652 5068
rect 15820 5058 15876 5068
rect 16380 5572 16436 5582
rect 16380 5236 16436 5516
rect 15596 4246 15652 4284
rect 16380 4338 16436 5180
rect 16604 5010 16660 5022
rect 16604 4958 16606 5010
rect 16658 4958 16660 5010
rect 16604 4562 16660 4958
rect 16604 4510 16606 4562
rect 16658 4510 16660 4562
rect 16604 4498 16660 4510
rect 16380 4286 16382 4338
rect 16434 4286 16436 4338
rect 16380 4274 16436 4286
rect 16604 4340 16660 4350
rect 16604 4338 16772 4340
rect 16604 4286 16606 4338
rect 16658 4286 16772 4338
rect 16604 4284 16772 4286
rect 16604 4274 16660 4284
rect 16716 3892 16772 4284
rect 16940 4338 16996 5740
rect 17724 5684 17780 5694
rect 16940 4286 16942 4338
rect 16994 4286 16996 4338
rect 16940 4274 16996 4286
rect 17164 4900 17220 4910
rect 16716 3836 16996 3892
rect 16156 3666 16212 3678
rect 16156 3614 16158 3666
rect 16210 3614 16212 3666
rect 16156 3388 16212 3614
rect 16940 3554 16996 3836
rect 16940 3502 16942 3554
rect 16994 3502 16996 3554
rect 16940 3490 16996 3502
rect 17164 3442 17220 4844
rect 17340 4732 17604 4742
rect 17396 4676 17444 4732
rect 17500 4676 17548 4732
rect 17340 4666 17604 4676
rect 17724 4564 17780 5628
rect 17948 5572 18004 5966
rect 17948 5506 18004 5516
rect 18172 5964 18788 6020
rect 17276 4508 17780 4564
rect 17276 3554 17332 4508
rect 18172 4450 18228 5964
rect 18396 5794 18452 5806
rect 18396 5742 18398 5794
rect 18450 5742 18452 5794
rect 18396 5684 18452 5742
rect 18396 5124 18452 5628
rect 18844 5460 18900 7422
rect 18844 5394 18900 5404
rect 18396 5058 18452 5068
rect 18732 5234 18788 5246
rect 18732 5182 18734 5234
rect 18786 5182 18788 5234
rect 18732 4900 18788 5182
rect 18956 5122 19012 7644
rect 19068 5908 19124 8990
rect 19180 8260 19236 12796
rect 19628 12178 19684 13132
rect 19628 12126 19630 12178
rect 19682 12126 19684 12178
rect 19628 12114 19684 12126
rect 19964 13132 20076 13188
rect 19964 12068 20020 13132
rect 20076 13122 20132 13132
rect 20188 12178 20244 13468
rect 20188 12126 20190 12178
rect 20242 12126 20244 12178
rect 20188 12114 20244 12126
rect 19964 11506 20020 12012
rect 19964 11454 19966 11506
rect 20018 11454 20020 11506
rect 19964 11442 20020 11454
rect 19740 10836 19796 10846
rect 20188 10836 20244 10846
rect 19740 10742 19796 10780
rect 19852 10834 20244 10836
rect 19852 10782 20190 10834
rect 20242 10782 20244 10834
rect 19852 10780 20244 10782
rect 19404 10724 19460 10734
rect 19292 10722 19460 10724
rect 19292 10670 19406 10722
rect 19458 10670 19460 10722
rect 19292 10668 19460 10670
rect 19292 9828 19348 10668
rect 19404 10658 19460 10668
rect 19852 10276 19908 10780
rect 20188 10770 20244 10780
rect 19740 10220 19908 10276
rect 19964 10610 20020 10622
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19404 9940 19460 9950
rect 19404 9938 19684 9940
rect 19404 9886 19406 9938
rect 19458 9886 19684 9938
rect 19404 9884 19684 9886
rect 19404 9874 19460 9884
rect 19292 9762 19348 9772
rect 19180 8194 19236 8204
rect 19628 9044 19684 9884
rect 19740 9154 19796 10220
rect 19964 10052 20020 10558
rect 20300 10612 20356 10622
rect 20300 10518 20356 10556
rect 20524 10610 20580 10622
rect 20524 10558 20526 10610
rect 20578 10558 20580 10610
rect 20524 10052 20580 10558
rect 20636 10276 20692 13580
rect 20860 13412 20916 13422
rect 20860 13074 20916 13356
rect 20860 13022 20862 13074
rect 20914 13022 20916 13074
rect 20860 13010 20916 13022
rect 21084 13300 21140 13580
rect 21084 12964 21140 13244
rect 21196 13188 21252 14476
rect 21308 14420 21364 14430
rect 21308 13636 21364 14364
rect 21420 14308 21476 14318
rect 21420 14214 21476 14252
rect 21868 14084 21924 14094
rect 21644 13858 21700 13870
rect 21644 13806 21646 13858
rect 21698 13806 21700 13858
rect 21644 13748 21700 13806
rect 21644 13682 21700 13692
rect 21756 13860 21812 13870
rect 21756 13746 21812 13804
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 21756 13682 21812 13694
rect 21308 13570 21364 13580
rect 21372 13356 21636 13366
rect 21428 13300 21476 13356
rect 21532 13300 21580 13356
rect 21372 13290 21636 13300
rect 21196 13132 21476 13188
rect 21420 13074 21476 13132
rect 21420 13022 21422 13074
rect 21474 13022 21476 13074
rect 21420 13010 21476 13022
rect 21308 12964 21364 12974
rect 21084 12962 21364 12964
rect 21084 12910 21310 12962
rect 21362 12910 21364 12962
rect 21084 12908 21364 12910
rect 21308 12898 21364 12908
rect 21868 11956 21924 14028
rect 21980 13074 22036 15036
rect 22092 14308 22148 15484
rect 22428 15428 22484 19180
rect 22988 19142 23044 19180
rect 23100 19180 23268 19236
rect 22876 19010 22932 19022
rect 22876 18958 22878 19010
rect 22930 18958 22932 19010
rect 22764 18564 22820 18574
rect 22764 18470 22820 18508
rect 22876 17892 22932 18958
rect 22764 17836 22932 17892
rect 22988 18788 23044 18798
rect 23100 18788 23156 19180
rect 23324 19124 23380 19134
rect 23548 19124 23604 19134
rect 23324 19122 23548 19124
rect 23324 19070 23326 19122
rect 23378 19070 23548 19122
rect 23324 19068 23548 19070
rect 23324 19058 23380 19068
rect 23548 19058 23604 19068
rect 23212 19010 23268 19022
rect 23212 18958 23214 19010
rect 23266 18958 23268 19010
rect 23212 18900 23268 18958
rect 23660 18900 23716 19292
rect 23884 19234 23940 20076
rect 24108 19684 24164 24668
rect 24332 24658 24388 24668
rect 24220 23828 24276 23838
rect 24220 23734 24276 23772
rect 24444 23044 24500 23054
rect 24556 23044 24612 26852
rect 24668 25396 24724 25406
rect 24668 24946 24724 25340
rect 24668 24894 24670 24946
rect 24722 24894 24724 24946
rect 24668 24882 24724 24894
rect 24444 23042 24612 23044
rect 24444 22990 24446 23042
rect 24498 22990 24612 23042
rect 24444 22988 24612 22990
rect 24444 22978 24500 22988
rect 24444 22372 24500 22382
rect 24332 22316 24444 22372
rect 24220 21700 24276 21710
rect 24220 21606 24276 21644
rect 24220 20916 24276 20926
rect 24332 20916 24388 22316
rect 24444 22306 24500 22316
rect 24444 21700 24500 21710
rect 24444 21606 24500 21644
rect 24220 20914 24500 20916
rect 24220 20862 24222 20914
rect 24274 20862 24500 20914
rect 24220 20860 24500 20862
rect 24220 20850 24276 20860
rect 24108 19348 24164 19628
rect 24108 19282 24164 19292
rect 24220 20020 24276 20030
rect 24220 19906 24276 19964
rect 24220 19854 24222 19906
rect 24274 19854 24276 19906
rect 23884 19182 23886 19234
rect 23938 19182 23940 19234
rect 23884 19170 23940 19182
rect 24220 19124 24276 19854
rect 24332 19460 24388 19470
rect 24332 19366 24388 19404
rect 24444 19234 24500 20860
rect 24444 19182 24446 19234
rect 24498 19182 24500 19234
rect 24444 19170 24500 19182
rect 24332 19124 24388 19134
rect 24220 19122 24388 19124
rect 24220 19070 24334 19122
rect 24386 19070 24388 19122
rect 24220 19068 24388 19070
rect 24332 19058 24388 19068
rect 23212 18844 23380 18900
rect 23324 18788 23380 18844
rect 23100 18732 23268 18788
rect 22540 17556 22596 17566
rect 22540 17462 22596 17500
rect 22764 16882 22820 17836
rect 22988 17780 23044 18732
rect 22764 16830 22766 16882
rect 22818 16830 22820 16882
rect 22652 16100 22708 16110
rect 22652 16006 22708 16044
rect 22540 15988 22596 15998
rect 22540 15894 22596 15932
rect 22204 15372 22484 15428
rect 22204 15092 22260 15372
rect 22428 15204 22484 15242
rect 22428 15092 22708 15148
rect 22204 15026 22260 15036
rect 22652 14418 22708 15092
rect 22652 14366 22654 14418
rect 22706 14366 22708 14418
rect 22652 14354 22708 14366
rect 22092 14252 22260 14308
rect 22204 14084 22260 14252
rect 22204 14018 22260 14028
rect 22092 13972 22148 13982
rect 22092 13858 22148 13916
rect 22092 13806 22094 13858
rect 22146 13806 22148 13858
rect 22092 13794 22148 13806
rect 21980 13022 21982 13074
rect 22034 13022 22036 13074
rect 21980 13010 22036 13022
rect 22092 13636 22148 13646
rect 22092 13076 22148 13580
rect 22204 13524 22260 13534
rect 22204 13522 22708 13524
rect 22204 13470 22206 13522
rect 22258 13470 22708 13522
rect 22204 13468 22708 13470
rect 22204 13458 22260 13468
rect 22428 13188 22484 13198
rect 22428 13094 22484 13132
rect 22652 13186 22708 13468
rect 22652 13134 22654 13186
rect 22706 13134 22708 13186
rect 22652 13122 22708 13134
rect 22316 13076 22372 13086
rect 22092 13074 22372 13076
rect 22092 13022 22318 13074
rect 22370 13022 22372 13074
rect 22092 13020 22372 13022
rect 22316 12964 22372 13020
rect 22316 12908 22596 12964
rect 22540 12402 22596 12908
rect 22540 12350 22542 12402
rect 22594 12350 22596 12402
rect 22540 12338 22596 12350
rect 21868 11890 21924 11900
rect 21372 11788 21636 11798
rect 21428 11732 21476 11788
rect 21532 11732 21580 11788
rect 21372 11722 21636 11732
rect 21532 11396 21588 11406
rect 21532 11302 21588 11340
rect 21868 11170 21924 11182
rect 21868 11118 21870 11170
rect 21922 11118 21924 11170
rect 21308 10836 21364 10846
rect 21308 10742 21364 10780
rect 20972 10722 21028 10734
rect 20972 10670 20974 10722
rect 21026 10670 21028 10722
rect 20972 10612 21028 10670
rect 20972 10546 21028 10556
rect 21868 10610 21924 11118
rect 22316 11170 22372 11182
rect 22316 11118 22318 11170
rect 22370 11118 22372 11170
rect 22316 10612 22372 11118
rect 21868 10558 21870 10610
rect 21922 10558 21924 10610
rect 21868 10276 21924 10558
rect 20636 10220 20804 10276
rect 19740 9102 19742 9154
rect 19794 9102 19796 9154
rect 19740 9090 19796 9102
rect 19852 9996 20020 10052
rect 20188 9996 20580 10052
rect 20636 10052 20692 10062
rect 19628 8258 19684 8988
rect 19628 8206 19630 8258
rect 19682 8206 19684 8258
rect 19628 8194 19684 8206
rect 19740 8260 19796 8270
rect 19852 8260 19908 9996
rect 20076 9940 20132 9950
rect 20188 9940 20244 9996
rect 20076 9938 20244 9940
rect 20076 9886 20078 9938
rect 20130 9886 20244 9938
rect 20076 9884 20244 9886
rect 20076 9874 20132 9884
rect 19964 9828 20020 9838
rect 20300 9828 20356 9838
rect 19964 9734 20020 9772
rect 20188 9772 20300 9828
rect 20188 9714 20244 9772
rect 20300 9762 20356 9772
rect 20636 9826 20692 9996
rect 20636 9774 20638 9826
rect 20690 9774 20692 9826
rect 20188 9662 20190 9714
rect 20242 9662 20244 9714
rect 20188 9650 20244 9662
rect 20636 9604 20692 9774
rect 20636 9538 20692 9548
rect 20748 8260 20804 10220
rect 21372 10220 21636 10230
rect 21428 10164 21476 10220
rect 21532 10164 21580 10220
rect 21868 10210 21924 10220
rect 22092 10556 22372 10612
rect 21372 10154 21636 10164
rect 21868 9828 21924 9838
rect 21868 8930 21924 9772
rect 21868 8878 21870 8930
rect 21922 8878 21924 8930
rect 21868 8866 21924 8878
rect 21372 8652 21636 8662
rect 21428 8596 21476 8652
rect 21532 8596 21580 8652
rect 21372 8586 21636 8596
rect 19852 8204 20020 8260
rect 19292 8148 19348 8158
rect 19292 8036 19348 8092
rect 19404 8036 19460 8046
rect 19180 8034 19460 8036
rect 19180 7982 19406 8034
rect 19458 7982 19460 8034
rect 19180 7980 19460 7982
rect 19180 7476 19236 7980
rect 19404 7970 19460 7980
rect 19516 8034 19572 8046
rect 19516 7982 19518 8034
rect 19570 7982 19572 8034
rect 19516 7924 19572 7982
rect 19516 7858 19572 7868
rect 19740 7700 19796 8204
rect 19852 8036 19908 8046
rect 19852 7942 19908 7980
rect 19964 7924 20020 8204
rect 20412 8204 20804 8260
rect 21980 8482 22036 8494
rect 21980 8430 21982 8482
rect 22034 8430 22036 8482
rect 20300 8148 20356 8158
rect 20300 8054 20356 8092
rect 19964 7858 20020 7868
rect 19852 7700 19908 7710
rect 19740 7698 19908 7700
rect 19740 7646 19854 7698
rect 19906 7646 19908 7698
rect 19740 7644 19908 7646
rect 19852 7634 19908 7644
rect 20300 7700 20356 7710
rect 20412 7700 20468 8204
rect 21868 8148 21924 8158
rect 21868 8054 21924 8092
rect 20300 7698 20468 7700
rect 20300 7646 20302 7698
rect 20354 7646 20468 7698
rect 20300 7644 20468 7646
rect 20636 8034 20692 8046
rect 20636 7982 20638 8034
rect 20690 7982 20692 8034
rect 20636 7700 20692 7982
rect 19292 7588 19348 7598
rect 19292 7494 19348 7532
rect 20076 7588 20132 7598
rect 19180 7410 19236 7420
rect 19404 7474 19460 7486
rect 19404 7422 19406 7474
rect 19458 7422 19460 7474
rect 19404 7364 19460 7422
rect 19460 7308 19572 7364
rect 19404 7298 19460 7308
rect 19068 5814 19124 5852
rect 19292 7250 19348 7262
rect 19292 7198 19294 7250
rect 19346 7198 19348 7250
rect 19292 5796 19348 7198
rect 19292 5730 19348 5740
rect 18956 5070 18958 5122
rect 19010 5070 19012 5122
rect 18956 5058 19012 5070
rect 19292 5012 19348 5022
rect 19516 5012 19572 7308
rect 19740 6020 19796 6030
rect 19740 5926 19796 5964
rect 19740 5460 19796 5470
rect 19796 5404 19908 5460
rect 19740 5394 19796 5404
rect 19852 5124 19908 5404
rect 19964 5124 20020 5134
rect 19852 5122 20020 5124
rect 19852 5070 19966 5122
rect 20018 5070 20020 5122
rect 19852 5068 20020 5070
rect 19964 5058 20020 5068
rect 19628 5012 19684 5022
rect 19516 5010 19684 5012
rect 19516 4958 19630 5010
rect 19682 4958 19684 5010
rect 19516 4956 19684 4958
rect 19292 4918 19348 4956
rect 19628 4946 19684 4956
rect 18732 4834 18788 4844
rect 19180 4898 19236 4910
rect 19180 4846 19182 4898
rect 19234 4846 19236 4898
rect 18172 4398 18174 4450
rect 18226 4398 18228 4450
rect 18172 4386 18228 4398
rect 17388 4340 17444 4350
rect 17388 4246 17444 4284
rect 19180 4228 19236 4846
rect 19180 4162 19236 4172
rect 19740 4900 19796 4910
rect 19740 4116 19796 4844
rect 19740 4050 19796 4060
rect 17276 3502 17278 3554
rect 17330 3502 17332 3554
rect 17276 3490 17332 3502
rect 18172 3666 18228 3678
rect 18172 3614 18174 3666
rect 18226 3614 18228 3666
rect 17164 3390 17166 3442
rect 17218 3390 17220 3442
rect 16156 3332 16660 3388
rect 17164 3378 17220 3390
rect 16604 800 16660 3332
rect 17340 3164 17604 3174
rect 17396 3108 17444 3164
rect 17500 3108 17548 3164
rect 17340 3098 17604 3108
rect 18172 800 18228 3614
rect 19852 3668 19908 3678
rect 19852 3388 19908 3612
rect 20076 3554 20132 7532
rect 20300 5234 20356 7644
rect 20636 7634 20692 7644
rect 21644 7812 21700 7822
rect 21644 7698 21700 7756
rect 21644 7646 21646 7698
rect 21698 7646 21700 7698
rect 21644 7634 21700 7646
rect 21756 7588 21812 7598
rect 21756 7494 21812 7532
rect 21308 7364 21364 7374
rect 21084 7362 21364 7364
rect 21084 7310 21310 7362
rect 21362 7310 21364 7362
rect 21084 7308 21364 7310
rect 20748 6804 20804 6814
rect 20748 6710 20804 6748
rect 20300 5182 20302 5234
rect 20354 5182 20356 5234
rect 20300 5124 20356 5182
rect 20300 5058 20356 5068
rect 20748 5908 20804 5918
rect 20748 5234 20804 5852
rect 20748 5182 20750 5234
rect 20802 5182 20804 5234
rect 20748 4340 20804 5182
rect 20860 4340 20916 4350
rect 20748 4284 20860 4340
rect 20860 4246 20916 4284
rect 20300 4228 20356 4238
rect 20300 4134 20356 4172
rect 20076 3502 20078 3554
rect 20130 3502 20132 3554
rect 20076 3490 20132 3502
rect 20748 4116 20804 4126
rect 20748 3554 20804 4060
rect 21084 3780 21140 7308
rect 21308 7298 21364 7308
rect 21644 7252 21700 7262
rect 21644 7250 21812 7252
rect 21644 7198 21646 7250
rect 21698 7198 21812 7250
rect 21644 7196 21812 7198
rect 21644 7186 21700 7196
rect 21372 7084 21636 7094
rect 21428 7028 21476 7084
rect 21532 7028 21580 7084
rect 21372 7018 21636 7028
rect 21644 6692 21700 6702
rect 21756 6692 21812 7196
rect 21980 6804 22036 8430
rect 22092 8260 22148 10556
rect 22540 10500 22596 10510
rect 22540 10406 22596 10444
rect 22316 10276 22372 10286
rect 22204 9940 22260 9950
rect 22204 9846 22260 9884
rect 22316 9268 22372 10220
rect 22764 10164 22820 16830
rect 22876 17724 23044 17780
rect 23100 18450 23156 18462
rect 23100 18398 23102 18450
rect 23154 18398 23156 18450
rect 22876 15764 22932 17724
rect 22988 17554 23044 17566
rect 22988 17502 22990 17554
rect 23042 17502 23044 17554
rect 22988 17332 23044 17502
rect 22988 17266 23044 17276
rect 23100 16884 23156 18398
rect 23212 17780 23268 18732
rect 23324 18722 23380 18732
rect 23436 18844 23716 18900
rect 23772 19010 23828 19022
rect 23772 18958 23774 19010
rect 23826 18958 23828 19010
rect 23772 18900 23828 18958
rect 23436 18564 23492 18844
rect 23772 18834 23828 18844
rect 24556 18788 24612 22988
rect 24892 24500 24948 24510
rect 24892 22482 24948 24444
rect 24892 22430 24894 22482
rect 24946 22430 24948 22482
rect 24668 21698 24724 21710
rect 24668 21646 24670 21698
rect 24722 21646 24724 21698
rect 24668 20804 24724 21646
rect 24892 21476 24948 22430
rect 24892 21410 24948 21420
rect 24780 21364 24836 21374
rect 24780 21270 24836 21308
rect 24668 20748 24836 20804
rect 24668 20580 24724 20590
rect 24668 20486 24724 20524
rect 24780 19796 24836 20748
rect 24892 20578 24948 20590
rect 24892 20526 24894 20578
rect 24946 20526 24948 20578
rect 24892 20132 24948 20526
rect 24892 20066 24948 20076
rect 24780 19730 24836 19740
rect 25004 19460 25060 27356
rect 25228 26964 25284 27694
rect 25340 27074 25396 28028
rect 25788 27990 25844 28028
rect 25452 27972 25508 27982
rect 25452 27858 25508 27916
rect 25452 27806 25454 27858
rect 25506 27806 25508 27858
rect 25452 27794 25508 27806
rect 25900 27860 25956 28590
rect 25900 27794 25956 27804
rect 26012 27186 26068 28700
rect 26012 27134 26014 27186
rect 26066 27134 26068 27186
rect 26012 27122 26068 27134
rect 26124 28308 26180 28318
rect 26124 28082 26180 28252
rect 26124 28030 26126 28082
rect 26178 28030 26180 28082
rect 25340 27022 25342 27074
rect 25394 27022 25396 27074
rect 25340 27010 25396 27022
rect 25228 26898 25284 26908
rect 25788 26740 25844 26750
rect 25404 26684 25668 26694
rect 25460 26628 25508 26684
rect 25564 26628 25612 26684
rect 25404 26618 25668 26628
rect 25340 26292 25396 26302
rect 25340 26198 25396 26236
rect 25228 25284 25284 25294
rect 25228 24722 25284 25228
rect 25404 25116 25668 25126
rect 25460 25060 25508 25116
rect 25564 25060 25612 25116
rect 25404 25050 25668 25060
rect 25564 24948 25620 24958
rect 25564 24854 25620 24892
rect 25228 24670 25230 24722
rect 25282 24670 25284 24722
rect 25228 23492 25284 24670
rect 25404 23548 25668 23558
rect 25460 23492 25508 23548
rect 25564 23492 25612 23548
rect 25404 23482 25668 23492
rect 25228 23268 25284 23436
rect 25228 23202 25284 23212
rect 25452 23156 25508 23166
rect 25452 22484 25508 23100
rect 25564 23156 25620 23166
rect 25788 23156 25844 26684
rect 26124 25508 26180 28030
rect 26236 28082 26292 29150
rect 26348 29204 26404 29372
rect 26348 29138 26404 29148
rect 26572 29426 26628 30156
rect 26572 29374 26574 29426
rect 26626 29374 26628 29426
rect 26572 29092 26628 29374
rect 26572 29026 26628 29036
rect 26796 28644 26852 31388
rect 27356 29764 27412 34200
rect 28364 30994 28420 31006
rect 28364 30942 28366 30994
rect 28418 30942 28420 30994
rect 27692 30322 27748 30334
rect 27692 30270 27694 30322
rect 27746 30270 27748 30322
rect 27356 29708 27636 29764
rect 27356 29316 27412 29326
rect 27356 29314 27524 29316
rect 27356 29262 27358 29314
rect 27410 29262 27524 29314
rect 27356 29260 27524 29262
rect 27356 29250 27412 29260
rect 26908 28868 26964 28878
rect 26908 28774 26964 28812
rect 26796 28588 26964 28644
rect 26460 28532 26516 28542
rect 26236 28030 26238 28082
rect 26290 28030 26292 28082
rect 26236 28018 26292 28030
rect 26348 28420 26404 28430
rect 26348 28082 26404 28364
rect 26348 28030 26350 28082
rect 26402 28030 26404 28082
rect 26348 28018 26404 28030
rect 26460 27972 26516 28476
rect 26460 27878 26516 27916
rect 26796 28420 26852 28430
rect 26124 25442 26180 25452
rect 26572 25732 26628 25742
rect 26572 25506 26628 25676
rect 26572 25454 26574 25506
rect 26626 25454 26628 25506
rect 26572 25442 26628 25454
rect 26124 25172 26180 25182
rect 25900 23940 25956 23950
rect 25900 23604 25956 23884
rect 25900 23538 25956 23548
rect 25564 23154 25844 23156
rect 25564 23102 25566 23154
rect 25618 23102 25844 23154
rect 25564 23100 25844 23102
rect 25564 23090 25620 23100
rect 25452 22370 25508 22428
rect 25452 22318 25454 22370
rect 25506 22318 25508 22370
rect 25452 22306 25508 22318
rect 25564 22596 25620 22606
rect 25564 22482 25620 22540
rect 25564 22430 25566 22482
rect 25618 22430 25620 22482
rect 25228 22260 25284 22270
rect 25116 22148 25172 22158
rect 25116 22054 25172 22092
rect 25228 21924 25284 22204
rect 25564 22148 25620 22430
rect 25564 22082 25620 22092
rect 25788 22484 25844 22494
rect 24892 19404 25060 19460
rect 25116 21868 25284 21924
rect 25404 21980 25668 21990
rect 25460 21924 25508 21980
rect 25564 21924 25612 21980
rect 25404 21914 25668 21924
rect 24892 18900 24948 19404
rect 25116 19346 25172 21868
rect 25788 21812 25844 22428
rect 25452 21756 25844 21812
rect 25900 22370 25956 22382
rect 25900 22318 25902 22370
rect 25954 22318 25956 22370
rect 25340 21700 25396 21710
rect 25340 21606 25396 21644
rect 25228 21586 25284 21598
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 25228 21476 25284 21534
rect 25340 21476 25396 21486
rect 25228 21420 25340 21476
rect 25340 21410 25396 21420
rect 25340 20804 25396 20814
rect 25452 20804 25508 21756
rect 25788 21588 25844 21598
rect 25788 21494 25844 21532
rect 25900 21476 25956 22318
rect 26124 22148 26180 25116
rect 26124 22082 26180 22092
rect 26236 24388 26292 24398
rect 26124 21476 26180 21486
rect 25900 21474 26180 21476
rect 25900 21422 26126 21474
rect 26178 21422 26180 21474
rect 25900 21420 26180 21422
rect 25340 20802 25508 20804
rect 25340 20750 25342 20802
rect 25394 20750 25508 20802
rect 25340 20748 25508 20750
rect 25676 20804 25732 20814
rect 26012 20804 26068 21420
rect 26124 21410 26180 21420
rect 26124 20916 26180 20926
rect 26124 20822 26180 20860
rect 25676 20802 26068 20804
rect 25676 20750 25678 20802
rect 25730 20750 26068 20802
rect 25676 20748 26068 20750
rect 25340 20738 25396 20748
rect 25676 20738 25732 20748
rect 25404 20412 25668 20422
rect 25460 20356 25508 20412
rect 25564 20356 25612 20412
rect 25404 20346 25668 20356
rect 25340 20244 25396 20254
rect 25340 20150 25396 20188
rect 25676 20244 25732 20254
rect 25676 20150 25732 20188
rect 25116 19294 25118 19346
rect 25170 19294 25172 19346
rect 25116 19282 25172 19294
rect 25452 19348 25508 19358
rect 25004 19234 25060 19246
rect 25004 19182 25006 19234
rect 25058 19182 25060 19234
rect 25004 19124 25060 19182
rect 25004 19058 25060 19068
rect 25452 19122 25508 19292
rect 25788 19348 25844 20748
rect 26236 20132 26292 24332
rect 26796 24162 26852 28364
rect 26908 28196 26964 28588
rect 26908 28130 26964 28140
rect 26908 27860 26964 27870
rect 26908 27766 26964 27804
rect 27244 27858 27300 27870
rect 27244 27806 27246 27858
rect 27298 27806 27300 27858
rect 26908 27524 26964 27534
rect 26908 26402 26964 27468
rect 27244 26908 27300 27806
rect 26908 26350 26910 26402
rect 26962 26350 26964 26402
rect 26908 26338 26964 26350
rect 27132 26852 27300 26908
rect 27356 27076 27412 27086
rect 27132 25956 27188 26852
rect 27356 25956 27412 27020
rect 27132 25890 27188 25900
rect 27244 25900 27412 25956
rect 27244 25732 27300 25900
rect 27132 25676 27300 25732
rect 27356 25732 27412 25742
rect 27020 25506 27076 25518
rect 27020 25454 27022 25506
rect 27074 25454 27076 25506
rect 27020 25396 27076 25454
rect 27020 25330 27076 25340
rect 26796 24110 26798 24162
rect 26850 24110 26852 24162
rect 26348 24052 26404 24062
rect 26348 24050 26516 24052
rect 26348 23998 26350 24050
rect 26402 23998 26516 24050
rect 26348 23996 26516 23998
rect 26348 23986 26404 23996
rect 26348 21812 26404 21822
rect 26460 21812 26516 23996
rect 26404 21756 26516 21812
rect 26572 23604 26628 23614
rect 26348 21746 26404 21756
rect 26572 21476 26628 23548
rect 26796 22260 26852 24110
rect 27020 24052 27076 24062
rect 27020 23958 27076 23996
rect 26796 22166 26852 22204
rect 26908 23940 26964 23950
rect 26572 20356 26628 21420
rect 26796 22036 26852 22046
rect 26796 20916 26852 21980
rect 26908 21586 26964 23884
rect 26908 21534 26910 21586
rect 26962 21534 26964 21586
rect 26908 21140 26964 21534
rect 26908 21074 26964 21084
rect 27020 23716 27076 23726
rect 27020 22146 27076 23660
rect 27020 22094 27022 22146
rect 27074 22094 27076 22146
rect 27020 21474 27076 22094
rect 27132 22820 27188 25676
rect 27244 25508 27300 25518
rect 27244 25414 27300 25452
rect 27244 24948 27300 24958
rect 27244 24388 27300 24892
rect 27356 24610 27412 25676
rect 27468 25618 27524 29260
rect 27580 28420 27636 29708
rect 27692 28644 27748 30270
rect 28364 30212 28420 30942
rect 28364 30146 28420 30156
rect 28476 30100 28532 34200
rect 28476 30034 28532 30044
rect 28700 31220 28756 31230
rect 27692 28578 27748 28588
rect 28028 29986 28084 29998
rect 28028 29934 28030 29986
rect 28082 29934 28084 29986
rect 27580 28354 27636 28364
rect 27804 26964 27860 26974
rect 27804 25730 27860 26908
rect 27804 25678 27806 25730
rect 27858 25678 27860 25730
rect 27804 25666 27860 25678
rect 27468 25566 27470 25618
rect 27522 25566 27524 25618
rect 27468 25554 27524 25566
rect 27580 25394 27636 25406
rect 27580 25342 27582 25394
rect 27634 25342 27636 25394
rect 27580 25284 27636 25342
rect 27580 25218 27636 25228
rect 27356 24558 27358 24610
rect 27410 24558 27412 24610
rect 27356 24546 27412 24558
rect 27468 25060 27524 25070
rect 27244 24332 27412 24388
rect 27356 23938 27412 24332
rect 27356 23886 27358 23938
rect 27410 23886 27412 23938
rect 27356 23874 27412 23886
rect 27244 23828 27300 23838
rect 27244 23734 27300 23772
rect 27356 23380 27412 23390
rect 27132 22258 27188 22764
rect 27244 22932 27300 22942
rect 27244 22484 27300 22876
rect 27356 22820 27412 23324
rect 27468 23042 27524 25004
rect 27692 24724 27748 24734
rect 28028 24724 28084 29934
rect 28364 29986 28420 29998
rect 28364 29934 28366 29986
rect 28418 29934 28420 29986
rect 28140 27860 28196 27870
rect 28140 27186 28196 27804
rect 28140 27134 28142 27186
rect 28194 27134 28196 27186
rect 28140 25506 28196 27134
rect 28252 27636 28308 27646
rect 28252 26740 28308 27580
rect 28364 27412 28420 29934
rect 28588 28644 28644 28654
rect 28364 27346 28420 27356
rect 28476 27748 28532 27758
rect 28476 27298 28532 27692
rect 28476 27246 28478 27298
rect 28530 27246 28532 27298
rect 28476 27234 28532 27246
rect 28588 27186 28644 28588
rect 28588 27134 28590 27186
rect 28642 27134 28644 27186
rect 28588 27122 28644 27134
rect 28252 25956 28308 26684
rect 28476 26180 28532 26190
rect 28476 26178 28644 26180
rect 28476 26126 28478 26178
rect 28530 26126 28644 26178
rect 28476 26124 28644 26126
rect 28476 26114 28532 26124
rect 28252 25900 28532 25956
rect 28140 25454 28142 25506
rect 28194 25454 28196 25506
rect 28140 25442 28196 25454
rect 28252 25618 28308 25630
rect 28252 25566 28254 25618
rect 28306 25566 28308 25618
rect 28140 24724 28196 24734
rect 28028 24722 28196 24724
rect 28028 24670 28142 24722
rect 28194 24670 28196 24722
rect 28028 24668 28196 24670
rect 27580 23826 27636 23838
rect 27580 23774 27582 23826
rect 27634 23774 27636 23826
rect 27580 23156 27636 23774
rect 27692 23380 27748 24668
rect 28140 24658 28196 24668
rect 27692 23314 27748 23324
rect 28028 23938 28084 23950
rect 28028 23886 28030 23938
rect 28082 23886 28084 23938
rect 27580 23100 27860 23156
rect 27468 22990 27470 23042
rect 27522 22990 27524 23042
rect 27468 22978 27524 22990
rect 27804 22932 27860 23100
rect 27580 22876 27860 22932
rect 27356 22764 27524 22820
rect 27244 22428 27412 22484
rect 27132 22206 27134 22258
rect 27186 22206 27188 22258
rect 27132 22036 27188 22206
rect 27132 21970 27188 21980
rect 27244 22258 27300 22270
rect 27244 22206 27246 22258
rect 27298 22206 27300 22258
rect 27244 21924 27300 22206
rect 27244 21858 27300 21868
rect 27020 21422 27022 21474
rect 27074 21422 27076 21474
rect 27020 20916 27076 21422
rect 27132 21698 27188 21710
rect 27356 21700 27412 22428
rect 27132 21646 27134 21698
rect 27186 21646 27188 21698
rect 27132 21476 27188 21646
rect 27132 21410 27188 21420
rect 27244 21644 27412 21700
rect 26796 20860 26964 20916
rect 26908 20802 26964 20860
rect 26908 20750 26910 20802
rect 26962 20750 26964 20802
rect 26796 20690 26852 20702
rect 26796 20638 26798 20690
rect 26850 20638 26852 20690
rect 26796 20580 26852 20638
rect 26796 20514 26852 20524
rect 26572 20290 26628 20300
rect 26908 20188 26964 20750
rect 27020 20692 27076 20860
rect 27244 20914 27300 21644
rect 27468 21588 27524 22764
rect 27580 22482 27636 22876
rect 27916 22820 27972 22830
rect 27916 22596 27972 22764
rect 28028 22708 28084 23886
rect 28252 23380 28308 25566
rect 28364 25284 28420 25294
rect 28364 25190 28420 25228
rect 28476 25172 28532 25900
rect 28588 25396 28644 26124
rect 28700 25732 28756 31164
rect 29148 31108 29204 31118
rect 29148 31014 29204 31052
rect 29260 30996 29316 31006
rect 29260 30210 29316 30940
rect 29596 30772 29652 34200
rect 30492 31108 30548 31118
rect 29596 30716 30212 30772
rect 29436 30604 29700 30614
rect 29492 30548 29540 30604
rect 29596 30548 29644 30604
rect 29436 30538 29700 30548
rect 29260 30158 29262 30210
rect 29314 30158 29316 30210
rect 29260 28868 29316 30158
rect 29596 30212 29652 30222
rect 29596 30118 29652 30156
rect 29484 29316 29540 29326
rect 29484 29314 30100 29316
rect 29484 29262 29486 29314
rect 29538 29262 30100 29314
rect 29484 29260 30100 29262
rect 29484 29250 29540 29260
rect 29436 29036 29700 29046
rect 29492 28980 29540 29036
rect 29596 28980 29644 29036
rect 29436 28970 29700 28980
rect 29596 28868 29652 28878
rect 29260 28812 29428 28868
rect 29148 28756 29204 28766
rect 29204 28700 29316 28756
rect 29148 28690 29204 28700
rect 29148 28420 29204 28430
rect 28700 25666 28756 25676
rect 28812 28418 29204 28420
rect 28812 28366 29150 28418
rect 29202 28366 29204 28418
rect 28812 28364 29204 28366
rect 28812 26290 28868 28364
rect 29148 28354 29204 28364
rect 29260 27972 29316 28700
rect 29372 28532 29428 28812
rect 29372 28438 29428 28476
rect 29484 28812 29596 28868
rect 29484 28530 29540 28812
rect 29596 28802 29652 28812
rect 29932 28756 29988 28766
rect 29820 28754 29988 28756
rect 29820 28702 29934 28754
rect 29986 28702 29988 28754
rect 29820 28700 29988 28702
rect 29484 28478 29486 28530
rect 29538 28478 29540 28530
rect 28812 26238 28814 26290
rect 28866 26238 28868 26290
rect 28588 25302 28644 25340
rect 28700 25508 28756 25518
rect 28700 25172 28756 25452
rect 28476 25106 28532 25116
rect 28588 25116 28756 25172
rect 28476 23938 28532 23950
rect 28476 23886 28478 23938
rect 28530 23886 28532 23938
rect 28476 23604 28532 23886
rect 28476 23538 28532 23548
rect 28476 23380 28532 23390
rect 28252 23324 28420 23380
rect 28252 23156 28308 23166
rect 28252 23062 28308 23100
rect 28140 22932 28196 22942
rect 28140 22838 28196 22876
rect 28364 22820 28420 23324
rect 28476 23266 28532 23324
rect 28476 23214 28478 23266
rect 28530 23214 28532 23266
rect 28476 23202 28532 23214
rect 28588 22932 28644 25116
rect 28812 24052 28868 26238
rect 28924 27916 29316 27972
rect 29484 28308 29540 28478
rect 29484 27972 29540 28252
rect 28924 24724 28980 27916
rect 29484 27906 29540 27916
rect 29596 28530 29652 28542
rect 29596 28478 29598 28530
rect 29650 28478 29652 28530
rect 29596 27748 29652 28478
rect 29036 27692 29652 27748
rect 29036 26516 29092 27692
rect 29436 27468 29700 27478
rect 29492 27412 29540 27468
rect 29596 27412 29644 27468
rect 29436 27402 29700 27412
rect 29596 27076 29652 27114
rect 29596 27010 29652 27020
rect 29260 26964 29316 27002
rect 29260 26898 29316 26908
rect 29372 26962 29428 26974
rect 29372 26910 29374 26962
rect 29426 26910 29428 26962
rect 29148 26850 29204 26862
rect 29148 26798 29150 26850
rect 29202 26798 29204 26850
rect 29148 26628 29204 26798
rect 29372 26740 29428 26910
rect 29820 26908 29876 28700
rect 29932 28690 29988 28700
rect 29372 26674 29428 26684
rect 29596 26852 29876 26908
rect 29932 27076 29988 27086
rect 30044 27076 30100 29260
rect 30156 28532 30212 30716
rect 30156 28466 30212 28476
rect 30268 30212 30324 30222
rect 30268 28642 30324 30156
rect 30380 30098 30436 30110
rect 30380 30046 30382 30098
rect 30434 30046 30436 30098
rect 30380 29540 30436 30046
rect 30380 29474 30436 29484
rect 30268 28590 30270 28642
rect 30322 28590 30324 28642
rect 29932 27074 30100 27076
rect 29932 27022 29934 27074
rect 29986 27022 30100 27074
rect 29932 27020 30100 27022
rect 30156 28308 30212 28318
rect 29484 26628 29540 26638
rect 29148 26572 29316 26628
rect 29036 26460 29204 26516
rect 29148 26404 29204 26460
rect 29036 26292 29092 26302
rect 29036 26068 29092 26236
rect 29036 26002 29092 26012
rect 29036 25844 29092 25854
rect 29036 25508 29092 25788
rect 29148 25620 29204 26348
rect 29260 25844 29316 26572
rect 29484 26290 29540 26572
rect 29596 26402 29652 26852
rect 29596 26350 29598 26402
rect 29650 26350 29652 26402
rect 29596 26338 29652 26350
rect 29820 26628 29876 26638
rect 29484 26238 29486 26290
rect 29538 26238 29540 26290
rect 29484 26226 29540 26238
rect 29484 26068 29540 26106
rect 29484 26002 29540 26012
rect 29436 25900 29700 25910
rect 29492 25844 29540 25900
rect 29596 25844 29644 25900
rect 29436 25834 29700 25844
rect 29260 25778 29316 25788
rect 29820 25732 29876 26572
rect 29596 25676 29876 25732
rect 29260 25620 29316 25630
rect 29148 25564 29260 25620
rect 29260 25554 29316 25564
rect 29036 25442 29092 25452
rect 29372 25506 29428 25518
rect 29372 25454 29374 25506
rect 29426 25454 29428 25506
rect 29372 25284 29428 25454
rect 29372 25218 29428 25228
rect 29596 24948 29652 25676
rect 29596 24882 29652 24892
rect 29708 25506 29764 25518
rect 29708 25454 29710 25506
rect 29762 25454 29764 25506
rect 29708 24724 29764 25454
rect 28924 24722 29316 24724
rect 28924 24670 28926 24722
rect 28978 24670 29316 24722
rect 28924 24668 29316 24670
rect 28924 24658 28980 24668
rect 28700 23156 28756 23166
rect 28812 23156 28868 23996
rect 29148 23940 29204 23950
rect 29148 23846 29204 23884
rect 29260 23604 29316 24668
rect 29708 24658 29764 24668
rect 29820 25282 29876 25294
rect 29820 25230 29822 25282
rect 29874 25230 29876 25282
rect 29436 24332 29700 24342
rect 29492 24276 29540 24332
rect 29596 24276 29644 24332
rect 29436 24266 29700 24276
rect 29708 24164 29764 24174
rect 29484 24108 29708 24164
rect 29484 23826 29540 24108
rect 29708 24098 29764 24108
rect 29820 23828 29876 25230
rect 29484 23774 29486 23826
rect 29538 23774 29540 23826
rect 29484 23762 29540 23774
rect 29708 23772 29876 23828
rect 29260 23548 29540 23604
rect 29484 23378 29540 23548
rect 29484 23326 29486 23378
rect 29538 23326 29540 23378
rect 29484 23314 29540 23326
rect 29372 23268 29428 23278
rect 29372 23174 29428 23212
rect 28700 23154 28868 23156
rect 28700 23102 28702 23154
rect 28754 23102 28868 23154
rect 28700 23100 28868 23102
rect 29484 23156 29540 23166
rect 28700 23090 28756 23100
rect 28924 22932 28980 22942
rect 28588 22930 28980 22932
rect 28588 22878 28926 22930
rect 28978 22878 28980 22930
rect 28588 22876 28980 22878
rect 28364 22754 28420 22764
rect 28028 22652 28308 22708
rect 28252 22596 28308 22652
rect 27916 22540 28084 22596
rect 28252 22540 28644 22596
rect 27580 22430 27582 22482
rect 27634 22430 27636 22482
rect 27580 22418 27636 22430
rect 27804 22484 27860 22494
rect 27860 22428 27972 22484
rect 27804 22418 27860 22428
rect 27244 20862 27246 20914
rect 27298 20862 27300 20914
rect 27244 20850 27300 20862
rect 27356 21252 27412 21262
rect 27356 20802 27412 21196
rect 27356 20750 27358 20802
rect 27410 20750 27412 20802
rect 27356 20738 27412 20750
rect 27132 20692 27188 20702
rect 27020 20690 27188 20692
rect 27020 20638 27134 20690
rect 27186 20638 27188 20690
rect 27020 20636 27188 20638
rect 27132 20626 27188 20636
rect 26124 20076 26292 20132
rect 26572 20132 26964 20188
rect 27244 20356 27300 20366
rect 27244 20132 27300 20300
rect 26012 19796 26068 19806
rect 26012 19702 26068 19740
rect 25788 19282 25844 19292
rect 25452 19070 25454 19122
rect 25506 19070 25508 19122
rect 25452 19058 25508 19070
rect 26012 19236 26068 19246
rect 26124 19236 26180 20076
rect 26236 19908 26292 19918
rect 26236 19906 26516 19908
rect 26236 19854 26238 19906
rect 26290 19854 26516 19906
rect 26236 19852 26516 19854
rect 26236 19842 26292 19852
rect 26460 19572 26516 19852
rect 26012 19234 26180 19236
rect 26012 19182 26014 19234
rect 26066 19182 26180 19234
rect 26012 19180 26180 19182
rect 26236 19348 26292 19358
rect 25788 18900 25844 18910
rect 24892 18844 25060 18900
rect 24556 18732 24948 18788
rect 24108 18676 24164 18686
rect 23436 18450 23492 18508
rect 23436 18398 23438 18450
rect 23490 18398 23492 18450
rect 23436 18386 23492 18398
rect 23772 18564 23828 18574
rect 23772 18450 23828 18508
rect 24108 18562 24164 18620
rect 24108 18510 24110 18562
rect 24162 18510 24164 18562
rect 24108 18498 24164 18510
rect 23772 18398 23774 18450
rect 23826 18398 23828 18450
rect 23772 18386 23828 18398
rect 24668 18450 24724 18462
rect 24668 18398 24670 18450
rect 24722 18398 24724 18450
rect 23436 18228 23492 18238
rect 23212 17666 23268 17724
rect 23212 17614 23214 17666
rect 23266 17614 23268 17666
rect 23212 17602 23268 17614
rect 23324 18226 23492 18228
rect 23324 18174 23438 18226
rect 23490 18174 23492 18226
rect 23324 18172 23492 18174
rect 23212 16884 23268 16894
rect 23100 16828 23212 16884
rect 23212 16098 23268 16828
rect 23324 16436 23380 18172
rect 23436 18162 23492 18172
rect 24668 17668 24724 18398
rect 24780 17780 24836 17790
rect 24780 17686 24836 17724
rect 23884 17556 23940 17566
rect 23436 17442 23492 17454
rect 23436 17390 23438 17442
rect 23490 17390 23492 17442
rect 23436 16884 23492 17390
rect 23436 16818 23492 16828
rect 23548 16996 23604 17006
rect 23548 16772 23604 16940
rect 23548 16678 23604 16716
rect 23660 16994 23716 17006
rect 23660 16942 23662 16994
rect 23714 16942 23716 16994
rect 23324 16380 23492 16436
rect 23212 16046 23214 16098
rect 23266 16046 23268 16098
rect 23212 16034 23268 16046
rect 23212 15876 23268 15886
rect 22876 15708 23044 15764
rect 22876 15540 22932 15550
rect 22876 15446 22932 15484
rect 22988 14980 23044 15708
rect 23212 15538 23268 15820
rect 23212 15486 23214 15538
rect 23266 15486 23268 15538
rect 23212 15474 23268 15486
rect 23436 15148 23492 16380
rect 23548 16324 23604 16334
rect 23548 16230 23604 16268
rect 23548 15428 23604 15438
rect 23660 15428 23716 16942
rect 23884 16994 23940 17500
rect 23996 17556 24052 17566
rect 23996 17554 24164 17556
rect 23996 17502 23998 17554
rect 24050 17502 24164 17554
rect 23996 17500 24164 17502
rect 23996 17490 24052 17500
rect 23884 16942 23886 16994
rect 23938 16942 23940 16994
rect 23884 16930 23940 16942
rect 24108 16882 24164 17500
rect 24108 16830 24110 16882
rect 24162 16830 24164 16882
rect 24108 16436 24164 16830
rect 23604 15372 23716 15428
rect 23772 16380 24164 16436
rect 24220 17442 24276 17454
rect 24220 17390 24222 17442
rect 24274 17390 24276 17442
rect 23548 15334 23604 15372
rect 23772 15148 23828 16380
rect 23884 16098 23940 16110
rect 24108 16100 24164 16110
rect 23884 16046 23886 16098
rect 23938 16046 23940 16098
rect 23884 15540 23940 16046
rect 23884 15474 23940 15484
rect 23996 16098 24164 16100
rect 23996 16046 24110 16098
rect 24162 16046 24164 16098
rect 23996 16044 24164 16046
rect 22988 14914 23044 14924
rect 23212 15092 23492 15148
rect 23548 15092 23828 15148
rect 23884 15316 23940 15326
rect 23884 15148 23940 15260
rect 23996 15148 24052 16044
rect 24108 16034 24164 16044
rect 24220 15876 24276 17390
rect 24444 17442 24500 17454
rect 24444 17390 24446 17442
rect 24498 17390 24500 17442
rect 24444 16772 24500 17390
rect 24556 17444 24612 17454
rect 24556 17350 24612 17388
rect 24556 17108 24612 17118
rect 24668 17108 24724 17612
rect 24556 17106 24724 17108
rect 24556 17054 24558 17106
rect 24610 17054 24724 17106
rect 24556 17052 24724 17054
rect 24556 17042 24612 17052
rect 24444 16706 24500 16716
rect 24780 16098 24836 16110
rect 24780 16046 24782 16098
rect 24834 16046 24836 16098
rect 24556 15988 24612 15998
rect 24444 15876 24500 15886
rect 24220 15874 24500 15876
rect 24220 15822 24446 15874
rect 24498 15822 24500 15874
rect 24220 15820 24500 15822
rect 24108 15764 24164 15774
rect 24108 15426 24164 15708
rect 24108 15374 24110 15426
rect 24162 15374 24164 15426
rect 24108 15362 24164 15374
rect 24444 15428 24500 15820
rect 24444 15362 24500 15372
rect 23884 15092 24052 15148
rect 24220 15314 24276 15326
rect 24220 15262 24222 15314
rect 24274 15262 24276 15314
rect 22876 14532 22932 14542
rect 22876 13970 22932 14476
rect 23212 14084 23268 15092
rect 22876 13918 22878 13970
rect 22930 13918 22932 13970
rect 22876 13906 22932 13918
rect 22988 14028 23268 14084
rect 23436 14530 23492 14542
rect 23436 14478 23438 14530
rect 23490 14478 23492 14530
rect 22988 13412 23044 14028
rect 23324 13972 23380 13982
rect 23100 13858 23156 13870
rect 23100 13806 23102 13858
rect 23154 13806 23156 13858
rect 23100 13748 23156 13806
rect 23156 13692 23268 13748
rect 23100 13682 23156 13692
rect 22876 13356 23044 13412
rect 22876 12516 22932 13356
rect 22988 13186 23044 13198
rect 22988 13134 22990 13186
rect 23042 13134 23044 13186
rect 22988 12964 23044 13134
rect 23100 12964 23156 12974
rect 22988 12962 23156 12964
rect 22988 12910 23102 12962
rect 23154 12910 23156 12962
rect 22988 12908 23156 12910
rect 23212 12964 23268 13692
rect 23324 13746 23380 13916
rect 23436 13860 23492 14478
rect 23436 13794 23492 13804
rect 23324 13694 23326 13746
rect 23378 13694 23380 13746
rect 23324 13682 23380 13694
rect 23548 13074 23604 15092
rect 23772 14532 23828 14542
rect 23772 14438 23828 14476
rect 23660 14418 23716 14430
rect 23660 14366 23662 14418
rect 23714 14366 23716 14418
rect 23660 13748 23716 14366
rect 23884 13970 23940 15092
rect 23884 13918 23886 13970
rect 23938 13918 23940 13970
rect 23884 13906 23940 13918
rect 23996 13972 24052 13982
rect 23772 13860 23828 13870
rect 23772 13766 23828 13804
rect 23660 13682 23716 13692
rect 23996 13746 24052 13916
rect 24220 13972 24276 15262
rect 24556 15148 24612 15932
rect 24668 15876 24724 15886
rect 24668 15538 24724 15820
rect 24668 15486 24670 15538
rect 24722 15486 24724 15538
rect 24668 15474 24724 15486
rect 24780 15316 24836 16046
rect 24780 15250 24836 15260
rect 24892 15148 24948 18732
rect 25004 18452 25060 18844
rect 25404 18844 25668 18854
rect 25460 18788 25508 18844
rect 25564 18788 25612 18844
rect 25404 18778 25668 18788
rect 25004 18386 25060 18396
rect 25452 18452 25508 18462
rect 25788 18452 25844 18844
rect 25452 18450 25844 18452
rect 25452 18398 25454 18450
rect 25506 18398 25844 18450
rect 25452 18396 25844 18398
rect 25900 18452 25956 18462
rect 25452 18340 25508 18396
rect 25900 18358 25956 18396
rect 25452 18274 25508 18284
rect 25900 17668 25956 17678
rect 25340 17556 25396 17566
rect 25340 17462 25396 17500
rect 25900 17554 25956 17612
rect 25900 17502 25902 17554
rect 25954 17502 25956 17554
rect 25900 17490 25956 17502
rect 25788 17442 25844 17454
rect 25788 17390 25790 17442
rect 25842 17390 25844 17442
rect 25404 17276 25668 17286
rect 25460 17220 25508 17276
rect 25564 17220 25612 17276
rect 25404 17210 25668 17220
rect 25116 16772 25172 16782
rect 25116 16212 25172 16716
rect 25564 16660 25620 16670
rect 25564 16566 25620 16604
rect 24556 15092 24724 15148
rect 24220 13906 24276 13916
rect 24668 14642 24724 15092
rect 24668 14590 24670 14642
rect 24722 14590 24724 14642
rect 23996 13694 23998 13746
rect 24050 13694 24052 13746
rect 23548 13022 23550 13074
rect 23602 13022 23604 13074
rect 23548 13010 23604 13022
rect 23772 13300 23828 13310
rect 23996 13300 24052 13694
rect 23828 13244 24052 13300
rect 24332 13746 24388 13758
rect 24332 13694 24334 13746
rect 24386 13694 24388 13746
rect 23324 12964 23380 12974
rect 23212 12908 23324 12964
rect 23100 12898 23156 12908
rect 23324 12870 23380 12908
rect 23772 12962 23828 13244
rect 24220 13188 24276 13198
rect 24332 13188 24388 13694
rect 24276 13132 24388 13188
rect 24220 13122 24276 13132
rect 23772 12910 23774 12962
rect 23826 12910 23828 12962
rect 23772 12898 23828 12910
rect 23996 12964 24052 12974
rect 23996 12870 24052 12908
rect 24556 12964 24612 12974
rect 24556 12870 24612 12908
rect 22876 12460 23268 12516
rect 22876 10836 22932 12460
rect 23212 12404 23268 12460
rect 23212 12310 23268 12348
rect 23884 12404 23940 12414
rect 23884 12310 23940 12348
rect 22876 10770 22932 10780
rect 23548 12290 23604 12302
rect 23548 12238 23550 12290
rect 23602 12238 23604 12290
rect 23324 10500 23380 10510
rect 23380 10444 23492 10500
rect 23324 10434 23380 10444
rect 22764 10098 22820 10108
rect 22988 10388 23044 10398
rect 22316 9174 22372 9212
rect 22540 9940 22596 9950
rect 22540 9826 22596 9884
rect 22540 9774 22542 9826
rect 22594 9774 22596 9826
rect 22540 8932 22596 9774
rect 22876 9604 22932 9614
rect 22988 9604 23044 10332
rect 23436 9938 23492 10444
rect 23436 9886 23438 9938
rect 23490 9886 23492 9938
rect 23436 9874 23492 9886
rect 23548 9940 23604 12238
rect 24220 12292 24276 12302
rect 24220 12198 24276 12236
rect 24668 12068 24724 14590
rect 24780 15092 24948 15148
rect 25004 16098 25060 16110
rect 25004 16046 25006 16098
rect 25058 16046 25060 16098
rect 25004 15988 25060 16046
rect 24780 12516 24836 15092
rect 25004 13412 25060 15932
rect 25116 15764 25172 16156
rect 25788 16100 25844 17390
rect 26012 17220 26068 19180
rect 26236 19122 26292 19292
rect 26236 19070 26238 19122
rect 26290 19070 26292 19122
rect 26236 19058 26292 19070
rect 26348 19122 26404 19134
rect 26348 19070 26350 19122
rect 26402 19070 26404 19122
rect 26124 19010 26180 19022
rect 26124 18958 26126 19010
rect 26178 18958 26180 19010
rect 26124 18564 26180 18958
rect 26124 18498 26180 18508
rect 26348 18450 26404 19070
rect 26460 18676 26516 19516
rect 26460 18562 26516 18620
rect 26460 18510 26462 18562
rect 26514 18510 26516 18562
rect 26460 18498 26516 18510
rect 26348 18398 26350 18450
rect 26402 18398 26404 18450
rect 26348 17780 26404 18398
rect 26236 17668 26292 17678
rect 25900 17164 26068 17220
rect 26124 17556 26180 17566
rect 26124 17220 26180 17500
rect 25900 16212 25956 17164
rect 26012 16996 26068 17006
rect 26012 16902 26068 16940
rect 26124 16994 26180 17164
rect 26124 16942 26126 16994
rect 26178 16942 26180 16994
rect 26124 16930 26180 16942
rect 26236 16994 26292 17612
rect 26236 16942 26238 16994
rect 26290 16942 26292 16994
rect 26236 16930 26292 16942
rect 26348 17556 26404 17724
rect 26460 17556 26516 17566
rect 26348 17554 26516 17556
rect 26348 17502 26462 17554
rect 26514 17502 26516 17554
rect 26348 17500 26516 17502
rect 26124 16660 26180 16670
rect 26180 16604 26292 16660
rect 26124 16594 26180 16604
rect 26012 16212 26068 16222
rect 25900 16210 26068 16212
rect 25900 16158 26014 16210
rect 26066 16158 26068 16210
rect 25900 16156 26068 16158
rect 25788 16044 25956 16100
rect 25564 15876 25620 15914
rect 25564 15810 25620 15820
rect 25116 15698 25172 15708
rect 25404 15708 25668 15718
rect 25460 15652 25508 15708
rect 25564 15652 25612 15708
rect 25404 15642 25668 15652
rect 25116 15540 25172 15550
rect 25116 15148 25172 15484
rect 25564 15540 25620 15550
rect 25564 15316 25620 15484
rect 25788 15428 25844 15438
rect 25788 15334 25844 15372
rect 25676 15316 25732 15326
rect 25620 15314 25732 15316
rect 25620 15262 25678 15314
rect 25730 15262 25732 15314
rect 25620 15260 25732 15262
rect 25564 15148 25620 15260
rect 25676 15250 25732 15260
rect 25116 15092 25284 15148
rect 25564 15092 25844 15148
rect 25228 15090 25284 15092
rect 25228 15038 25230 15090
rect 25282 15038 25284 15090
rect 25228 15026 25284 15038
rect 25676 14644 25732 14654
rect 25676 14550 25732 14588
rect 25404 14140 25668 14150
rect 25460 14084 25508 14140
rect 25564 14084 25612 14140
rect 25404 14074 25668 14084
rect 25452 13972 25508 13982
rect 25788 13972 25844 15092
rect 25900 14420 25956 16044
rect 26012 15988 26068 16156
rect 26012 15922 26068 15932
rect 26012 15652 26068 15662
rect 26012 15314 26068 15596
rect 26012 15262 26014 15314
rect 26066 15262 26068 15314
rect 26012 15250 26068 15262
rect 26124 15428 26180 15438
rect 25900 14354 25956 14364
rect 25452 13878 25508 13916
rect 25564 13916 25844 13972
rect 25564 13858 25620 13916
rect 25564 13806 25566 13858
rect 25618 13806 25620 13858
rect 25564 13794 25620 13806
rect 25228 13746 25284 13758
rect 25228 13694 25230 13746
rect 25282 13694 25284 13746
rect 25228 13636 25284 13694
rect 25228 13570 25284 13580
rect 26124 13634 26180 15372
rect 26124 13582 26126 13634
rect 26178 13582 26180 13634
rect 25004 13356 25284 13412
rect 24892 13188 24948 13198
rect 24892 12962 24948 13132
rect 24892 12910 24894 12962
rect 24946 12910 24948 12962
rect 24892 12898 24948 12910
rect 25228 12964 25284 13356
rect 26124 13076 26180 13582
rect 26124 13010 26180 13020
rect 25228 12850 25284 12908
rect 25676 12964 25732 12974
rect 25676 12962 25844 12964
rect 25676 12910 25678 12962
rect 25730 12910 25844 12962
rect 25676 12908 25844 12910
rect 25676 12898 25732 12908
rect 25228 12798 25230 12850
rect 25282 12798 25284 12850
rect 25228 12786 25284 12798
rect 25404 12572 25668 12582
rect 25460 12516 25508 12572
rect 25564 12516 25612 12572
rect 25404 12506 25668 12516
rect 24780 12450 24836 12460
rect 24556 12066 24724 12068
rect 24556 12014 24670 12066
rect 24722 12014 24724 12066
rect 24556 12012 24724 12014
rect 24556 10724 24612 12012
rect 24668 12002 24724 12012
rect 25228 12292 25284 12302
rect 24556 10658 24612 10668
rect 25004 11284 25060 11294
rect 24668 10612 24724 10622
rect 23548 9826 23604 9884
rect 23548 9774 23550 9826
rect 23602 9774 23604 9826
rect 23548 9762 23604 9774
rect 23884 10500 23940 10510
rect 23884 9826 23940 10444
rect 24668 10498 24724 10556
rect 24668 10446 24670 10498
rect 24722 10446 24724 10498
rect 24668 10434 24724 10446
rect 25004 10276 25060 11228
rect 24892 10164 24948 10174
rect 23884 9774 23886 9826
rect 23938 9774 23940 9826
rect 23884 9762 23940 9774
rect 24444 9828 24500 9838
rect 24444 9734 24500 9772
rect 24780 9826 24836 9838
rect 24780 9774 24782 9826
rect 24834 9774 24836 9826
rect 23324 9716 23380 9726
rect 23324 9622 23380 9660
rect 24332 9716 24388 9726
rect 24332 9622 24388 9660
rect 22876 9602 23044 9604
rect 22876 9550 22878 9602
rect 22930 9550 23044 9602
rect 22876 9548 23044 9550
rect 22876 9538 22932 9548
rect 22876 8932 22932 8942
rect 22540 8866 22596 8876
rect 22764 8930 22932 8932
rect 22764 8878 22878 8930
rect 22930 8878 22932 8930
rect 22764 8876 22932 8878
rect 22764 8482 22820 8876
rect 22876 8866 22932 8876
rect 22764 8430 22766 8482
rect 22818 8430 22820 8482
rect 22764 8418 22820 8430
rect 22316 8372 22372 8382
rect 22316 8278 22372 8316
rect 22092 8194 22148 8204
rect 22764 8036 22820 8046
rect 22652 8034 22820 8036
rect 22652 7982 22766 8034
rect 22818 7982 22820 8034
rect 22652 7980 22820 7982
rect 22092 7588 22148 7598
rect 22092 7494 22148 7532
rect 22316 7476 22372 7486
rect 22316 7474 22596 7476
rect 22316 7422 22318 7474
rect 22370 7422 22596 7474
rect 22316 7420 22596 7422
rect 22316 7410 22372 7420
rect 22204 7362 22260 7374
rect 22204 7310 22206 7362
rect 22258 7310 22260 7362
rect 22204 6916 22260 7310
rect 22204 6860 22484 6916
rect 21980 6748 22148 6804
rect 21644 6690 21812 6692
rect 21644 6638 21646 6690
rect 21698 6638 21812 6690
rect 21644 6636 21812 6638
rect 21644 6626 21700 6636
rect 21980 6578 22036 6590
rect 21980 6526 21982 6578
rect 22034 6526 22036 6578
rect 21756 6468 21812 6478
rect 21756 6374 21812 6412
rect 21980 6468 22036 6526
rect 21980 6402 22036 6412
rect 21868 5796 21924 5806
rect 21868 5702 21924 5740
rect 21372 5516 21636 5526
rect 21428 5460 21476 5516
rect 21532 5460 21580 5516
rect 21372 5450 21636 5460
rect 21308 5236 21364 5246
rect 21084 3714 21140 3724
rect 21196 5180 21308 5236
rect 20748 3502 20750 3554
rect 20802 3502 20804 3554
rect 20748 3490 20804 3502
rect 19740 3332 19908 3388
rect 21196 3388 21252 5180
rect 21308 5170 21364 5180
rect 21532 5122 21588 5134
rect 21532 5070 21534 5122
rect 21586 5070 21588 5122
rect 21532 4228 21588 5070
rect 21644 5124 21700 5134
rect 21644 4450 21700 5068
rect 21644 4398 21646 4450
rect 21698 4398 21700 4450
rect 21644 4386 21700 4398
rect 21532 4162 21588 4172
rect 21372 3948 21636 3958
rect 21428 3892 21476 3948
rect 21532 3892 21580 3948
rect 21372 3882 21636 3892
rect 22092 3892 22148 6748
rect 22428 6690 22484 6860
rect 22428 6638 22430 6690
rect 22482 6638 22484 6690
rect 22428 6626 22484 6638
rect 22540 6804 22596 7420
rect 22204 6580 22260 6590
rect 22204 6578 22372 6580
rect 22204 6526 22206 6578
rect 22258 6526 22372 6578
rect 22204 6524 22372 6526
rect 22204 6514 22260 6524
rect 22204 6132 22260 6142
rect 22204 6038 22260 6076
rect 22316 6130 22372 6524
rect 22316 6078 22318 6130
rect 22370 6078 22372 6130
rect 22316 6066 22372 6078
rect 22428 6132 22484 6142
rect 22540 6132 22596 6748
rect 22652 6692 22708 7980
rect 22764 7970 22820 7980
rect 22876 8034 22932 8046
rect 22876 7982 22878 8034
rect 22930 7982 22932 8034
rect 22764 7476 22820 7486
rect 22764 7382 22820 7420
rect 22652 6626 22708 6636
rect 22764 6690 22820 6702
rect 22764 6638 22766 6690
rect 22818 6638 22820 6690
rect 22428 6130 22596 6132
rect 22428 6078 22430 6130
rect 22482 6078 22596 6130
rect 22428 6076 22596 6078
rect 22652 6466 22708 6478
rect 22652 6414 22654 6466
rect 22706 6414 22708 6466
rect 22428 6066 22484 6076
rect 22652 6020 22708 6414
rect 22764 6468 22820 6638
rect 22764 6402 22820 6412
rect 22876 6356 22932 7982
rect 22988 7140 23044 9548
rect 24220 9602 24276 9614
rect 24220 9550 24222 9602
rect 24274 9550 24276 9602
rect 24220 9492 24276 9550
rect 24220 9436 24500 9492
rect 23772 9268 23828 9278
rect 23548 9156 23604 9166
rect 23548 9154 23716 9156
rect 23548 9102 23550 9154
rect 23602 9102 23716 9154
rect 23548 9100 23716 9102
rect 23548 9090 23604 9100
rect 23212 8930 23268 8942
rect 23212 8878 23214 8930
rect 23266 8878 23268 8930
rect 23212 8820 23268 8878
rect 23212 8754 23268 8764
rect 23660 8708 23716 9100
rect 23772 9042 23828 9212
rect 23772 8990 23774 9042
rect 23826 8990 23828 9042
rect 23772 8978 23828 8990
rect 24332 9268 24388 9278
rect 24332 9042 24388 9212
rect 24444 9156 24500 9436
rect 24556 9156 24612 9166
rect 24444 9100 24556 9156
rect 24556 9062 24612 9100
rect 24332 8990 24334 9042
rect 24386 8990 24388 9042
rect 24332 8978 24388 8990
rect 24444 8932 24500 8942
rect 24500 8876 24612 8932
rect 24444 8866 24500 8876
rect 23324 8652 23716 8708
rect 23212 8260 23268 8270
rect 23324 8260 23380 8652
rect 23212 8258 23380 8260
rect 23212 8206 23214 8258
rect 23266 8206 23380 8258
rect 23212 8204 23380 8206
rect 23436 8484 23492 8494
rect 23212 8194 23268 8204
rect 23100 8034 23156 8046
rect 23100 7982 23102 8034
rect 23154 7982 23156 8034
rect 23100 7812 23156 7982
rect 23436 8034 23492 8428
rect 23660 8260 23716 8652
rect 23772 8260 23828 8270
rect 24332 8260 24388 8270
rect 23660 8258 24388 8260
rect 23660 8206 23774 8258
rect 23826 8206 24334 8258
rect 24386 8206 24388 8258
rect 23660 8204 24388 8206
rect 23772 8194 23828 8204
rect 23436 7982 23438 8034
rect 23490 7982 23492 8034
rect 23436 7970 23492 7982
rect 23660 8034 23716 8046
rect 23660 7982 23662 8034
rect 23714 7982 23716 8034
rect 23324 7812 23380 7822
rect 23100 7756 23324 7812
rect 23324 7698 23380 7756
rect 23324 7646 23326 7698
rect 23378 7646 23380 7698
rect 23324 7634 23380 7646
rect 23100 7476 23156 7486
rect 23100 7382 23156 7420
rect 23436 7476 23492 7486
rect 23436 7382 23492 7420
rect 23660 7364 23716 7982
rect 23996 8036 24052 8046
rect 23996 7942 24052 7980
rect 24220 8034 24276 8046
rect 24220 7982 24222 8034
rect 24274 7982 24276 8034
rect 23660 7298 23716 7308
rect 22988 7084 24164 7140
rect 23548 6804 23604 6814
rect 23436 6802 23604 6804
rect 23436 6750 23550 6802
rect 23602 6750 23604 6802
rect 23436 6748 23604 6750
rect 23100 6692 23156 6702
rect 23436 6692 23492 6748
rect 23548 6738 23604 6748
rect 23100 6690 23492 6692
rect 23100 6638 23102 6690
rect 23154 6638 23492 6690
rect 23100 6636 23492 6638
rect 24108 6690 24164 7084
rect 24220 6916 24276 7982
rect 24332 8036 24388 8204
rect 24332 7970 24388 7980
rect 24556 7700 24612 8876
rect 24780 8482 24836 9774
rect 24780 8430 24782 8482
rect 24834 8430 24836 8482
rect 24780 8418 24836 8430
rect 24668 8146 24724 8158
rect 24668 8094 24670 8146
rect 24722 8094 24724 8146
rect 24668 8036 24724 8094
rect 24668 7970 24724 7980
rect 24780 8034 24836 8046
rect 24780 7982 24782 8034
rect 24834 7982 24836 8034
rect 24668 7700 24724 7710
rect 24556 7698 24724 7700
rect 24556 7646 24670 7698
rect 24722 7646 24724 7698
rect 24556 7644 24724 7646
rect 24556 7476 24612 7486
rect 24332 7362 24388 7374
rect 24332 7310 24334 7362
rect 24386 7310 24388 7362
rect 24332 7140 24388 7310
rect 24332 7074 24388 7084
rect 24444 7364 24500 7374
rect 24220 6850 24276 6860
rect 24108 6638 24110 6690
rect 24162 6638 24164 6690
rect 23100 6626 23156 6636
rect 22876 6290 22932 6300
rect 23436 6466 23492 6478
rect 23436 6414 23438 6466
rect 23490 6414 23492 6466
rect 22652 5954 22708 5964
rect 22764 6244 22820 6254
rect 22764 5906 22820 6188
rect 23436 6132 23492 6414
rect 23660 6466 23716 6478
rect 23660 6414 23662 6466
rect 23714 6414 23716 6466
rect 23436 6066 23492 6076
rect 23548 6356 23604 6366
rect 23548 6130 23604 6300
rect 23548 6078 23550 6130
rect 23602 6078 23604 6130
rect 23548 6066 23604 6078
rect 22764 5854 22766 5906
rect 22818 5854 22820 5906
rect 22764 5842 22820 5854
rect 23100 5908 23156 5918
rect 23100 5814 23156 5852
rect 23324 5908 23380 5918
rect 23660 5908 23716 6414
rect 24108 6244 24164 6638
rect 24444 6578 24500 7308
rect 24556 6804 24612 7420
rect 24668 7364 24724 7644
rect 24780 7476 24836 7982
rect 24780 7410 24836 7420
rect 24668 7298 24724 7308
rect 24556 6690 24612 6748
rect 24556 6638 24558 6690
rect 24610 6638 24612 6690
rect 24556 6626 24612 6638
rect 24444 6526 24446 6578
rect 24498 6526 24500 6578
rect 24220 6466 24276 6478
rect 24220 6414 24222 6466
rect 24274 6414 24276 6466
rect 24220 6356 24276 6414
rect 24220 6290 24276 6300
rect 24444 6356 24500 6526
rect 24444 6290 24500 6300
rect 24780 6468 24836 6478
rect 24108 6130 24164 6188
rect 24108 6078 24110 6130
rect 24162 6078 24164 6130
rect 24108 6066 24164 6078
rect 24332 6132 24388 6142
rect 24388 6076 24612 6132
rect 24332 6066 24388 6076
rect 24556 6018 24612 6076
rect 24556 5966 24558 6018
rect 24610 5966 24612 6018
rect 24556 5954 24612 5966
rect 24332 5908 24388 5918
rect 23324 5906 23716 5908
rect 23324 5854 23326 5906
rect 23378 5854 23716 5906
rect 23324 5852 23716 5854
rect 23996 5906 24388 5908
rect 23996 5854 24334 5906
rect 24386 5854 24388 5906
rect 23996 5852 24388 5854
rect 23212 5794 23268 5806
rect 23212 5742 23214 5794
rect 23266 5742 23268 5794
rect 22540 5236 22596 5246
rect 22540 5142 22596 5180
rect 23212 5124 23268 5742
rect 23324 5796 23380 5852
rect 23324 5730 23380 5740
rect 23212 5058 23268 5068
rect 23660 5684 23716 5694
rect 22092 3826 22148 3836
rect 21868 3668 21924 3678
rect 21868 3574 21924 3612
rect 22876 3444 22932 3454
rect 21196 3332 21364 3388
rect 19740 800 19796 3332
rect 21308 800 21364 3332
rect 22876 800 22932 3388
rect 23660 3442 23716 5628
rect 23996 5012 24052 5852
rect 24332 5842 24388 5852
rect 24444 5796 24500 5806
rect 24444 5794 24724 5796
rect 24444 5742 24446 5794
rect 24498 5742 24724 5794
rect 24444 5740 24724 5742
rect 24444 5730 24500 5740
rect 23772 4228 23828 4238
rect 23996 4228 24052 4956
rect 24108 5572 24164 5582
rect 24108 4562 24164 5516
rect 24556 5236 24612 5246
rect 24556 5142 24612 5180
rect 24332 5124 24388 5134
rect 24332 5030 24388 5068
rect 24668 4900 24724 5740
rect 24780 5122 24836 6412
rect 24892 6244 24948 10108
rect 25004 8708 25060 10220
rect 25228 10610 25284 12236
rect 25340 12180 25396 12190
rect 25396 12124 25508 12180
rect 25340 12086 25396 12124
rect 25452 11284 25508 12124
rect 25788 11844 25844 12908
rect 25900 12740 25956 12750
rect 25900 12646 25956 12684
rect 26236 12516 26292 16604
rect 26348 15316 26404 17500
rect 26460 17490 26516 17500
rect 26572 17332 26628 20132
rect 27132 20130 27300 20132
rect 27132 20078 27246 20130
rect 27298 20078 27300 20130
rect 27132 20076 27300 20078
rect 26908 20020 26964 20030
rect 26796 19234 26852 19246
rect 26796 19182 26798 19234
rect 26850 19182 26852 19234
rect 26684 19012 26740 19022
rect 26684 18674 26740 18956
rect 26684 18622 26686 18674
rect 26738 18622 26740 18674
rect 26684 18610 26740 18622
rect 26796 18676 26852 19182
rect 26796 18610 26852 18620
rect 26908 18564 26964 19964
rect 27020 19908 27076 19918
rect 27020 19814 27076 19852
rect 27132 19572 27188 20076
rect 27244 20066 27300 20076
rect 27132 19506 27188 19516
rect 27356 20018 27412 20030
rect 27356 19966 27358 20018
rect 27410 19966 27412 20018
rect 27356 18788 27412 19966
rect 27468 18900 27524 21532
rect 27804 22260 27860 22270
rect 27692 21364 27748 21374
rect 27692 20914 27748 21308
rect 27692 20862 27694 20914
rect 27746 20862 27748 20914
rect 27692 20850 27748 20862
rect 27804 20692 27860 22204
rect 27916 22258 27972 22428
rect 27916 22206 27918 22258
rect 27970 22206 27972 22258
rect 27916 21924 27972 22206
rect 27916 21858 27972 21868
rect 27916 20804 27972 20814
rect 28028 20804 28084 22540
rect 28140 22372 28196 22382
rect 28140 22278 28196 22316
rect 28476 22260 28532 22270
rect 28476 22166 28532 22204
rect 28364 22146 28420 22158
rect 28364 22094 28366 22146
rect 28418 22094 28420 22146
rect 28364 22036 28420 22094
rect 28364 21980 28532 22036
rect 28252 21700 28308 21710
rect 27916 20802 28084 20804
rect 27916 20750 27918 20802
rect 27970 20750 28084 20802
rect 27916 20748 28084 20750
rect 28140 21476 28196 21486
rect 27916 20738 27972 20748
rect 27692 20636 27860 20692
rect 28140 20690 28196 21420
rect 28140 20638 28142 20690
rect 28194 20638 28196 20690
rect 27580 20132 27636 20142
rect 27580 19572 27636 20076
rect 27580 19506 27636 19516
rect 27692 19124 27748 20636
rect 28140 20626 28196 20638
rect 28252 20356 28308 21644
rect 28364 20804 28420 20814
rect 28476 20804 28532 21980
rect 28364 20802 28532 20804
rect 28364 20750 28366 20802
rect 28418 20750 28532 20802
rect 28364 20748 28532 20750
rect 28364 20738 28420 20748
rect 28588 20692 28644 22540
rect 28924 21252 28980 22876
rect 29484 22930 29540 23100
rect 29708 23044 29764 23772
rect 29932 23268 29988 27020
rect 29932 23154 29988 23212
rect 29932 23102 29934 23154
rect 29986 23102 29988 23154
rect 29932 23090 29988 23102
rect 30044 25508 30100 25518
rect 29708 22978 29764 22988
rect 29484 22878 29486 22930
rect 29538 22878 29540 22930
rect 29484 22866 29540 22878
rect 29436 22764 29700 22774
rect 29492 22708 29540 22764
rect 29596 22708 29644 22764
rect 29436 22698 29700 22708
rect 29484 22370 29540 22382
rect 29484 22318 29486 22370
rect 29538 22318 29540 22370
rect 29484 22260 29540 22318
rect 29484 22194 29540 22204
rect 29932 22258 29988 22270
rect 29932 22206 29934 22258
rect 29986 22206 29988 22258
rect 28924 21186 28980 21196
rect 29260 22146 29316 22158
rect 29260 22094 29262 22146
rect 29314 22094 29316 22146
rect 29148 20804 29204 20814
rect 29148 20710 29204 20748
rect 28140 20300 28308 20356
rect 28476 20636 28588 20692
rect 27916 19908 27972 19918
rect 27468 18834 27524 18844
rect 27580 19122 27748 19124
rect 27580 19070 27694 19122
rect 27746 19070 27748 19122
rect 27580 19068 27748 19070
rect 26908 18498 26964 18508
rect 27132 18732 27412 18788
rect 26796 17668 26852 17678
rect 26460 17276 26628 17332
rect 26684 17612 26796 17668
rect 26460 16212 26516 17276
rect 26572 17108 26628 17118
rect 26572 17014 26628 17052
rect 26684 16996 26740 17612
rect 26796 17574 26852 17612
rect 27020 17442 27076 17454
rect 27020 17390 27022 17442
rect 27074 17390 27076 17442
rect 27020 17332 27076 17390
rect 27020 17266 27076 17276
rect 26684 16930 26740 16940
rect 26796 17108 26852 17118
rect 26684 16212 26740 16222
rect 26460 16210 26740 16212
rect 26460 16158 26686 16210
rect 26738 16158 26740 16210
rect 26460 16156 26740 16158
rect 26684 16146 26740 16156
rect 26796 15428 26852 17052
rect 27132 17108 27188 18732
rect 27244 18564 27300 18574
rect 27580 18564 27636 19068
rect 27692 19058 27748 19068
rect 27804 19346 27860 19358
rect 27804 19294 27806 19346
rect 27858 19294 27860 19346
rect 27244 18562 27636 18564
rect 27244 18510 27246 18562
rect 27298 18510 27636 18562
rect 27244 18508 27636 18510
rect 27692 18564 27748 18574
rect 27244 17668 27300 18508
rect 27692 18470 27748 18508
rect 27468 18228 27524 18238
rect 27468 17890 27524 18172
rect 27468 17838 27470 17890
rect 27522 17838 27524 17890
rect 27468 17826 27524 17838
rect 27580 18226 27636 18238
rect 27580 18174 27582 18226
rect 27634 18174 27636 18226
rect 27244 17602 27300 17612
rect 27356 17444 27412 17454
rect 27412 17388 27524 17444
rect 27356 17378 27412 17388
rect 27132 17042 27188 17052
rect 27244 17332 27300 17342
rect 27020 16884 27076 16894
rect 27076 16828 27188 16884
rect 27020 16818 27076 16828
rect 27132 16212 27188 16828
rect 27020 16156 27188 16212
rect 27020 16098 27076 16156
rect 27020 16046 27022 16098
rect 27074 16046 27076 16098
rect 27020 16034 27076 16046
rect 26796 15362 26852 15372
rect 26908 15426 26964 15438
rect 26908 15374 26910 15426
rect 26962 15374 26964 15426
rect 26460 15316 26516 15326
rect 26348 15260 26460 15316
rect 26460 15250 26516 15260
rect 26572 15314 26628 15326
rect 26572 15262 26574 15314
rect 26626 15262 26628 15314
rect 26572 14756 26628 15262
rect 26572 14690 26628 14700
rect 26908 14756 26964 15374
rect 27244 15148 27300 17276
rect 27356 16884 27412 16894
rect 27356 16790 27412 16828
rect 27468 16882 27524 17388
rect 27468 16830 27470 16882
rect 27522 16830 27524 16882
rect 27468 16818 27524 16830
rect 27580 16660 27636 18174
rect 27692 17666 27748 17678
rect 27692 17614 27694 17666
rect 27746 17614 27748 17666
rect 27692 17444 27748 17614
rect 27692 17378 27748 17388
rect 27804 16996 27860 19294
rect 27916 18676 27972 19852
rect 28028 19460 28084 19470
rect 28028 19234 28084 19404
rect 28028 19182 28030 19234
rect 28082 19182 28084 19234
rect 28028 19170 28084 19182
rect 27916 18582 27972 18620
rect 27916 17892 27972 17902
rect 28140 17892 28196 20300
rect 28364 20132 28420 20142
rect 28476 20132 28532 20636
rect 28588 20626 28644 20636
rect 28364 20130 28532 20132
rect 28364 20078 28366 20130
rect 28418 20078 28532 20130
rect 28364 20076 28532 20078
rect 28700 20578 28756 20590
rect 28700 20526 28702 20578
rect 28754 20526 28756 20578
rect 28364 19908 28420 20076
rect 28364 19842 28420 19852
rect 28476 19236 28532 19246
rect 28364 19180 28476 19236
rect 28364 19122 28420 19180
rect 28476 19170 28532 19180
rect 28700 19236 28756 20526
rect 29260 20356 29316 22094
rect 29820 21588 29876 21598
rect 29436 21196 29700 21206
rect 29492 21140 29540 21196
rect 29596 21140 29644 21196
rect 29436 21130 29700 21140
rect 29260 20290 29316 20300
rect 29372 21028 29428 21038
rect 29372 20020 29428 20972
rect 29372 19954 29428 19964
rect 29820 20018 29876 21532
rect 29820 19966 29822 20018
rect 29874 19966 29876 20018
rect 29436 19628 29700 19638
rect 29492 19572 29540 19628
rect 29596 19572 29644 19628
rect 29436 19562 29700 19572
rect 29148 19460 29204 19470
rect 29148 19366 29204 19404
rect 29484 19460 29540 19470
rect 29820 19460 29876 19966
rect 29484 19236 29540 19404
rect 28700 19170 28756 19180
rect 29148 19234 29540 19236
rect 29148 19182 29486 19234
rect 29538 19182 29540 19234
rect 29148 19180 29540 19182
rect 28364 19070 28366 19122
rect 28418 19070 28420 19122
rect 28364 19058 28420 19070
rect 28476 19010 28532 19022
rect 28476 18958 28478 19010
rect 28530 18958 28532 19010
rect 28476 18900 28532 18958
rect 28476 18834 28532 18844
rect 28700 19010 28756 19022
rect 28700 18958 28702 19010
rect 28754 18958 28756 19010
rect 28700 18676 28756 18958
rect 29148 19012 29204 19180
rect 29484 19170 29540 19180
rect 29708 19404 29876 19460
rect 29932 20132 29988 22206
rect 29932 19684 29988 20076
rect 29148 18946 29204 18956
rect 29260 19010 29316 19022
rect 29260 18958 29262 19010
rect 29314 18958 29316 19010
rect 29260 18900 29316 18958
rect 29708 18900 29764 19404
rect 29260 18844 29764 18900
rect 28700 18610 28756 18620
rect 29596 18676 29652 18686
rect 28364 18564 28420 18574
rect 28420 18508 28532 18564
rect 28364 18498 28420 18508
rect 27916 17890 28196 17892
rect 27916 17838 27918 17890
rect 27970 17838 28196 17890
rect 27916 17836 28196 17838
rect 28252 18450 28308 18462
rect 28252 18398 28254 18450
rect 28306 18398 28308 18450
rect 28252 18340 28308 18398
rect 27916 17826 27972 17836
rect 26908 14690 26964 14700
rect 27132 15092 27300 15148
rect 27356 16604 27636 16660
rect 27692 16940 27860 16996
rect 27916 17668 27972 17678
rect 26908 14084 26964 14094
rect 26572 13748 26628 13758
rect 26572 13654 26628 13692
rect 26908 13746 26964 14028
rect 26908 13694 26910 13746
rect 26962 13694 26964 13746
rect 26908 13682 26964 13694
rect 27132 13412 27188 15092
rect 26908 13356 27188 13412
rect 26684 13300 26740 13310
rect 26460 13076 26516 13086
rect 26460 12982 26516 13020
rect 26684 13076 26740 13244
rect 26684 13010 26740 13020
rect 26572 12852 26628 12862
rect 26572 12758 26628 12796
rect 26908 12850 26964 13356
rect 26908 12798 26910 12850
rect 26962 12798 26964 12850
rect 26908 12786 26964 12798
rect 26348 12740 26404 12750
rect 26348 12646 26404 12684
rect 27244 12738 27300 12750
rect 27244 12686 27246 12738
rect 27298 12686 27300 12738
rect 27244 12628 27300 12686
rect 27244 12562 27300 12572
rect 26012 12460 26292 12516
rect 25900 11844 25956 11854
rect 25788 11788 25900 11844
rect 25900 11778 25956 11788
rect 26012 11620 26068 12460
rect 27356 12292 27412 16604
rect 27468 16210 27524 16222
rect 27468 16158 27470 16210
rect 27522 16158 27524 16210
rect 27468 15764 27524 16158
rect 27468 15698 27524 15708
rect 27692 15986 27748 16940
rect 27804 16772 27860 16782
rect 27804 16678 27860 16716
rect 27692 15934 27694 15986
rect 27746 15934 27748 15986
rect 27580 15314 27636 15326
rect 27580 15262 27582 15314
rect 27634 15262 27636 15314
rect 27580 14868 27636 15262
rect 27580 14802 27636 14812
rect 27244 12236 27412 12292
rect 27468 13748 27524 13758
rect 26124 12068 26180 12078
rect 26124 12066 26292 12068
rect 26124 12014 26126 12066
rect 26178 12014 26292 12066
rect 26124 12012 26292 12014
rect 26124 12002 26180 12012
rect 26012 11554 26068 11564
rect 25452 11218 25508 11228
rect 25404 11004 25668 11014
rect 25460 10948 25508 11004
rect 25564 10948 25612 11004
rect 25404 10938 25668 10948
rect 26236 10834 26292 12012
rect 27244 11732 27300 12236
rect 26236 10782 26238 10834
rect 26290 10782 26292 10834
rect 26236 10770 26292 10782
rect 26908 11676 27300 11732
rect 27356 11844 27412 11854
rect 25564 10724 25620 10734
rect 25228 10558 25230 10610
rect 25282 10558 25284 10610
rect 25228 10052 25284 10558
rect 25452 10612 25508 10622
rect 25452 10518 25508 10556
rect 25340 10500 25396 10510
rect 25340 10406 25396 10444
rect 25228 9986 25284 9996
rect 25452 9940 25508 9950
rect 25564 9940 25620 10668
rect 25508 9884 25620 9940
rect 25676 10722 25732 10734
rect 25676 10670 25678 10722
rect 25730 10670 25732 10722
rect 25676 9940 25732 10670
rect 26460 10724 26516 10734
rect 26460 10630 26516 10668
rect 26124 10610 26180 10622
rect 26124 10558 26126 10610
rect 26178 10558 26180 10610
rect 26012 10500 26068 10510
rect 25676 9884 25956 9940
rect 25452 9826 25508 9884
rect 25676 9828 25732 9884
rect 25452 9774 25454 9826
rect 25506 9774 25508 9826
rect 25452 9762 25508 9774
rect 25564 9772 25732 9828
rect 25228 9716 25284 9726
rect 25228 9622 25284 9660
rect 25340 9604 25396 9614
rect 25564 9604 25620 9772
rect 25788 9714 25844 9726
rect 25788 9662 25790 9714
rect 25842 9662 25844 9714
rect 25396 9548 25620 9604
rect 25676 9604 25732 9642
rect 25340 9538 25396 9548
rect 25676 9538 25732 9548
rect 25404 9436 25668 9446
rect 25460 9380 25508 9436
rect 25564 9380 25612 9436
rect 25404 9370 25668 9380
rect 25564 9268 25620 9278
rect 25564 9174 25620 9212
rect 25228 9154 25284 9166
rect 25228 9102 25230 9154
rect 25282 9102 25284 9154
rect 25116 8708 25172 8718
rect 25004 8652 25116 8708
rect 25116 8642 25172 8652
rect 25228 8484 25284 9102
rect 25116 8428 25284 8484
rect 25340 8708 25396 8718
rect 25116 7700 25172 8428
rect 25340 8370 25396 8652
rect 25340 8318 25342 8370
rect 25394 8318 25396 8370
rect 25340 8306 25396 8318
rect 25788 8372 25844 9662
rect 25900 9492 25956 9884
rect 25900 9426 25956 9436
rect 25788 8306 25844 8316
rect 26012 9042 26068 10444
rect 26124 9940 26180 10558
rect 26348 10612 26404 10622
rect 26236 9940 26292 9950
rect 26124 9938 26292 9940
rect 26124 9886 26238 9938
rect 26290 9886 26292 9938
rect 26124 9884 26292 9886
rect 26236 9874 26292 9884
rect 26348 9826 26404 10556
rect 26572 10612 26628 10622
rect 26572 10500 26628 10556
rect 26348 9774 26350 9826
rect 26402 9774 26404 9826
rect 26348 9762 26404 9774
rect 26460 10444 26628 10500
rect 26684 10610 26740 10622
rect 26684 10558 26686 10610
rect 26738 10558 26740 10610
rect 26124 9602 26180 9614
rect 26124 9550 26126 9602
rect 26178 9550 26180 9602
rect 26124 9156 26180 9550
rect 26124 9090 26180 9100
rect 26012 8990 26014 9042
rect 26066 8990 26068 9042
rect 25900 8034 25956 8046
rect 25900 7982 25902 8034
rect 25954 7982 25956 8034
rect 25404 7868 25668 7878
rect 25460 7812 25508 7868
rect 25564 7812 25612 7868
rect 25404 7802 25668 7812
rect 25116 7634 25172 7644
rect 25564 7586 25620 7598
rect 25564 7534 25566 7586
rect 25618 7534 25620 7586
rect 25228 7474 25284 7486
rect 25228 7422 25230 7474
rect 25282 7422 25284 7474
rect 25228 7364 25284 7422
rect 25228 7298 25284 7308
rect 25116 6468 25172 6478
rect 25340 6468 25396 6506
rect 24892 6178 24948 6188
rect 25004 6466 25172 6468
rect 25004 6414 25118 6466
rect 25170 6414 25172 6466
rect 25004 6412 25172 6414
rect 24780 5070 24782 5122
rect 24834 5070 24836 5122
rect 24780 5058 24836 5070
rect 24892 5122 24948 5134
rect 24892 5070 24894 5122
rect 24946 5070 24948 5122
rect 24892 4900 24948 5070
rect 24668 4844 24948 4900
rect 24108 4510 24110 4562
rect 24162 4510 24164 4562
rect 24108 4498 24164 4510
rect 24444 4564 24500 4574
rect 24500 4508 24612 4564
rect 24444 4498 24500 4508
rect 24556 4450 24612 4508
rect 24556 4398 24558 4450
rect 24610 4398 24612 4450
rect 24556 4386 24612 4398
rect 25004 4452 25060 6412
rect 25116 6402 25172 6412
rect 25228 6412 25340 6468
rect 25004 4386 25060 4396
rect 25116 6244 25172 6254
rect 23772 4226 24052 4228
rect 23772 4174 23774 4226
rect 23826 4174 24052 4226
rect 23772 4172 24052 4174
rect 24220 4228 24276 4238
rect 24668 4228 24724 4238
rect 24220 4226 24500 4228
rect 24220 4174 24222 4226
rect 24274 4174 24500 4226
rect 24220 4172 24500 4174
rect 23772 4162 23828 4172
rect 24220 4162 24276 4172
rect 23660 3390 23662 3442
rect 23714 3390 23716 3442
rect 23660 3378 23716 3390
rect 23996 3444 24052 3482
rect 24444 3444 24500 4172
rect 24668 4134 24724 4172
rect 24780 3556 24836 3566
rect 24892 3556 24948 3566
rect 24836 3554 24948 3556
rect 24836 3502 24894 3554
rect 24946 3502 24948 3554
rect 24836 3500 24948 3502
rect 24668 3444 24724 3454
rect 24444 3442 24724 3444
rect 24444 3390 24670 3442
rect 24722 3390 24724 3442
rect 24444 3388 24724 3390
rect 23996 3378 24052 3388
rect 24668 3378 24724 3388
rect 24780 980 24836 3500
rect 24892 3490 24948 3500
rect 25116 1204 25172 6188
rect 25228 6132 25284 6412
rect 25340 6402 25396 6412
rect 25564 6468 25620 7534
rect 25900 6916 25956 7982
rect 25900 6850 25956 6860
rect 26012 6804 26068 8990
rect 26236 8260 26292 8270
rect 26460 8260 26516 10444
rect 26684 9940 26740 10558
rect 26684 9874 26740 9884
rect 26796 9826 26852 9838
rect 26796 9774 26798 9826
rect 26850 9774 26852 9826
rect 26572 9604 26628 9614
rect 26628 9548 26740 9604
rect 26572 9538 26628 9548
rect 26684 9154 26740 9548
rect 26684 9102 26686 9154
rect 26738 9102 26740 9154
rect 26684 9090 26740 9102
rect 26796 8932 26852 9774
rect 26908 9268 26964 11676
rect 27244 11508 27300 11518
rect 27132 11394 27188 11406
rect 27132 11342 27134 11394
rect 27186 11342 27188 11394
rect 27132 10612 27188 11342
rect 27132 10518 27188 10556
rect 27020 10052 27076 10062
rect 27020 9826 27076 9996
rect 27132 9940 27188 9950
rect 27132 9846 27188 9884
rect 27020 9774 27022 9826
rect 27074 9774 27076 9826
rect 27020 9762 27076 9774
rect 27244 9826 27300 11452
rect 27244 9774 27246 9826
rect 27298 9774 27300 9826
rect 27244 9762 27300 9774
rect 27356 9604 27412 11788
rect 27468 10612 27524 13692
rect 27692 12964 27748 15934
rect 27916 15876 27972 17612
rect 28140 17668 28196 17678
rect 28140 17332 28196 17612
rect 28140 17266 28196 17276
rect 28252 17220 28308 18284
rect 28476 17668 28532 18508
rect 29148 18508 29540 18564
rect 28588 18452 28644 18462
rect 28588 18338 28644 18396
rect 28588 18286 28590 18338
rect 28642 18286 28644 18338
rect 28588 18274 28644 18286
rect 28700 18450 28756 18462
rect 28700 18398 28702 18450
rect 28754 18398 28756 18450
rect 28700 18116 28756 18398
rect 28700 18050 28756 18060
rect 28812 18228 28868 18238
rect 28588 18004 28644 18014
rect 28588 17780 28644 17948
rect 28588 17778 28756 17780
rect 28588 17726 28590 17778
rect 28642 17726 28756 17778
rect 28588 17724 28756 17726
rect 28588 17714 28644 17724
rect 28476 17602 28532 17612
rect 28252 17154 28308 17164
rect 28476 17444 28532 17454
rect 28364 17108 28420 17118
rect 28364 17014 28420 17052
rect 28476 16884 28532 17388
rect 28364 16828 28532 16884
rect 28028 16100 28084 16110
rect 28252 16100 28308 16110
rect 28028 16098 28196 16100
rect 28028 16046 28030 16098
rect 28082 16046 28196 16098
rect 28028 16044 28196 16046
rect 28028 16034 28084 16044
rect 27916 15820 28084 15876
rect 27916 15426 27972 15438
rect 27916 15374 27918 15426
rect 27970 15374 27972 15426
rect 27916 15204 27972 15374
rect 27916 15138 27972 15148
rect 27804 14418 27860 14430
rect 27804 14366 27806 14418
rect 27858 14366 27860 14418
rect 27804 13524 27860 14366
rect 27916 13860 27972 13870
rect 27916 13766 27972 13804
rect 27804 13458 27860 13468
rect 28028 13074 28084 15820
rect 28140 15538 28196 16044
rect 28252 16006 28308 16044
rect 28140 15486 28142 15538
rect 28194 15486 28196 15538
rect 28140 15474 28196 15486
rect 28252 15764 28308 15774
rect 28252 15538 28308 15708
rect 28252 15486 28254 15538
rect 28306 15486 28308 15538
rect 28252 15474 28308 15486
rect 28364 14980 28420 16828
rect 28700 16212 28756 17724
rect 28812 17106 28868 18172
rect 28812 17054 28814 17106
rect 28866 17054 28868 17106
rect 28812 17042 28868 17054
rect 28700 16146 28756 16156
rect 29148 16770 29204 18508
rect 29484 18452 29540 18508
rect 29484 18386 29540 18396
rect 29596 18450 29652 18620
rect 29596 18398 29598 18450
rect 29650 18398 29652 18450
rect 29596 18386 29652 18398
rect 29260 18340 29316 18350
rect 29260 17668 29316 18284
rect 29708 18340 29764 18844
rect 29932 18564 29988 19628
rect 30044 19234 30100 25452
rect 30156 24500 30212 28252
rect 30268 27970 30324 28590
rect 30268 27918 30270 27970
rect 30322 27918 30324 27970
rect 30268 27074 30324 27918
rect 30268 27022 30270 27074
rect 30322 27022 30324 27074
rect 30268 25506 30324 27022
rect 30268 25454 30270 25506
rect 30322 25454 30324 25506
rect 30268 25442 30324 25454
rect 30380 28420 30436 28430
rect 30156 24444 30324 24500
rect 30268 24164 30324 24444
rect 30268 24098 30324 24108
rect 30268 23940 30324 23950
rect 30268 23846 30324 23884
rect 30268 22372 30324 22382
rect 30268 22278 30324 22316
rect 30044 19182 30046 19234
rect 30098 19182 30100 19234
rect 30044 19170 30100 19182
rect 30156 22258 30212 22270
rect 30156 22206 30158 22258
rect 30210 22206 30212 22258
rect 30156 18900 30212 22206
rect 30268 21588 30324 21598
rect 30268 21494 30324 21532
rect 30380 20914 30436 28364
rect 30492 23380 30548 31052
rect 30604 30100 30660 30110
rect 30604 29538 30660 30044
rect 30604 29486 30606 29538
rect 30658 29486 30660 29538
rect 30604 29474 30660 29486
rect 30492 23314 30548 23324
rect 30604 28196 30660 28206
rect 30604 22932 30660 28140
rect 30716 26402 30772 34200
rect 30716 26350 30718 26402
rect 30770 26350 30772 26402
rect 30716 26338 30772 26350
rect 30828 28532 30884 28542
rect 30716 24948 30772 24958
rect 30716 24834 30772 24892
rect 30716 24782 30718 24834
rect 30770 24782 30772 24834
rect 30716 24770 30772 24782
rect 30828 24162 30884 28476
rect 30828 24110 30830 24162
rect 30882 24110 30884 24162
rect 30828 24098 30884 24110
rect 30940 23378 30996 34300
rect 31500 34132 31556 34300
rect 31808 34200 31920 35000
rect 32928 34200 33040 35000
rect 34048 34200 34160 35000
rect 31836 34132 31892 34200
rect 31500 34076 31892 34132
rect 32284 30996 32340 31006
rect 32732 30996 32788 31006
rect 32284 30994 32452 30996
rect 32284 30942 32286 30994
rect 32338 30942 32452 30994
rect 32284 30940 32452 30942
rect 32284 30930 32340 30940
rect 31276 30882 31332 30894
rect 31276 30830 31278 30882
rect 31330 30830 31332 30882
rect 31052 30324 31108 30334
rect 31052 28754 31108 30268
rect 31276 30324 31332 30830
rect 32172 30884 32228 30894
rect 32172 30790 32228 30828
rect 32284 30770 32340 30782
rect 32284 30718 32286 30770
rect 32338 30718 32340 30770
rect 31276 30258 31332 30268
rect 32172 30324 32228 30334
rect 31388 29652 31444 29662
rect 31276 28868 31332 28878
rect 31052 28702 31054 28754
rect 31106 28702 31108 28754
rect 31052 28690 31108 28702
rect 31164 28812 31276 28868
rect 31052 27188 31108 27198
rect 31164 27188 31220 28812
rect 31276 28802 31332 28812
rect 31052 27186 31220 27188
rect 31052 27134 31054 27186
rect 31106 27134 31220 27186
rect 31052 27132 31220 27134
rect 31276 28644 31332 28654
rect 31052 27122 31108 27132
rect 31052 26068 31108 26078
rect 31052 25618 31108 26012
rect 31052 25566 31054 25618
rect 31106 25566 31108 25618
rect 31052 25554 31108 25566
rect 31276 24948 31332 28588
rect 31276 24882 31332 24892
rect 31388 24612 31444 29596
rect 31948 29428 32004 29438
rect 31948 29334 32004 29372
rect 32172 26290 32228 30268
rect 32284 28868 32340 30718
rect 32396 29092 32452 30940
rect 32956 30996 33012 34200
rect 33468 31388 33732 31398
rect 33524 31332 33572 31388
rect 33628 31332 33676 31388
rect 33468 31322 33732 31332
rect 32956 30940 33348 30996
rect 32732 30902 32788 30940
rect 32956 30772 33012 30782
rect 32956 30678 33012 30716
rect 32844 30436 32900 30446
rect 32508 30322 32564 30334
rect 32508 30270 32510 30322
rect 32562 30270 32564 30322
rect 32508 29652 32564 30270
rect 32844 30098 32900 30380
rect 32844 30046 32846 30098
rect 32898 30046 32900 30098
rect 32844 30034 32900 30046
rect 33068 30210 33124 30222
rect 33068 30158 33070 30210
rect 33122 30158 33124 30210
rect 32508 29586 32564 29596
rect 32396 29026 32452 29036
rect 33068 28980 33124 30158
rect 33180 29316 33236 29326
rect 33180 29222 33236 29260
rect 33068 28914 33124 28924
rect 32284 28802 32340 28812
rect 33180 28756 33236 28766
rect 33180 28662 33236 28700
rect 33180 27746 33236 27758
rect 33180 27694 33182 27746
rect 33234 27694 33236 27746
rect 33180 27636 33236 27694
rect 33180 27570 33236 27580
rect 32172 26238 32174 26290
rect 32226 26238 32228 26290
rect 30940 23326 30942 23378
rect 30994 23326 30996 23378
rect 30940 23314 30996 23326
rect 31052 24556 31444 24612
rect 31948 24612 32004 24622
rect 30604 22876 30884 22932
rect 30380 20862 30382 20914
rect 30434 20862 30436 20914
rect 30380 20850 30436 20862
rect 30716 21474 30772 21486
rect 30716 21422 30718 21474
rect 30770 21422 30772 21474
rect 30268 20132 30324 20142
rect 30268 20018 30324 20076
rect 30268 19966 30270 20018
rect 30322 19966 30324 20018
rect 30268 19954 30324 19966
rect 30492 20130 30548 20142
rect 30492 20078 30494 20130
rect 30546 20078 30548 20130
rect 30268 19124 30324 19134
rect 30324 19068 30436 19124
rect 30268 19058 30324 19068
rect 30156 18834 30212 18844
rect 30380 18564 30436 19068
rect 30492 18788 30548 20078
rect 30492 18722 30548 18732
rect 30604 19236 30660 19246
rect 30492 18564 30548 18574
rect 30380 18562 30548 18564
rect 30380 18510 30494 18562
rect 30546 18510 30548 18562
rect 30380 18508 30548 18510
rect 29932 18498 29988 18508
rect 30492 18498 30548 18508
rect 30268 18450 30324 18462
rect 30268 18398 30270 18450
rect 30322 18398 30324 18450
rect 30044 18340 30100 18350
rect 29708 18274 29764 18284
rect 29932 18338 30100 18340
rect 29932 18286 30046 18338
rect 30098 18286 30100 18338
rect 29932 18284 30100 18286
rect 29820 18228 29876 18238
rect 29820 18134 29876 18172
rect 29436 18060 29700 18070
rect 29492 18004 29540 18060
rect 29596 18004 29644 18060
rect 29436 17994 29700 18004
rect 29260 17602 29316 17612
rect 29372 17892 29428 17902
rect 29372 16996 29428 17836
rect 29372 16902 29428 16940
rect 29820 17108 29876 17118
rect 29148 16718 29150 16770
rect 29202 16718 29204 16770
rect 28924 16100 28980 16110
rect 28980 16044 29092 16100
rect 28924 16034 28980 16044
rect 28588 15930 28644 15942
rect 28476 15874 28532 15886
rect 28476 15822 28478 15874
rect 28530 15822 28532 15874
rect 28476 15652 28532 15822
rect 28476 15586 28532 15596
rect 28588 15878 28590 15930
rect 28642 15878 28644 15930
rect 28476 15316 28532 15326
rect 28476 15222 28532 15260
rect 28252 14644 28308 14654
rect 28252 13746 28308 14588
rect 28252 13694 28254 13746
rect 28306 13694 28308 13746
rect 28252 13682 28308 13694
rect 28364 13636 28420 14924
rect 28588 14980 28644 15878
rect 28588 14914 28644 14924
rect 28700 15428 28756 15438
rect 28364 13570 28420 13580
rect 28476 14868 28532 14878
rect 28476 13412 28532 14812
rect 28588 14756 28644 14766
rect 28588 14530 28644 14700
rect 28588 14478 28590 14530
rect 28642 14478 28644 14530
rect 28588 13748 28644 14478
rect 28588 13682 28644 13692
rect 28028 13022 28030 13074
rect 28082 13022 28084 13074
rect 28028 13010 28084 13022
rect 28364 13356 28532 13412
rect 27468 10546 27524 10556
rect 27580 12908 27748 12964
rect 26908 9202 26964 9212
rect 27244 9548 27412 9604
rect 27468 9604 27524 9614
rect 26796 8876 26964 8932
rect 26292 8204 26516 8260
rect 26908 8260 26964 8876
rect 26908 8204 27188 8260
rect 26236 8166 26292 8204
rect 26796 8036 26852 8046
rect 26796 7942 26852 7980
rect 27132 7924 27188 8204
rect 27244 8146 27300 9548
rect 27468 9510 27524 9548
rect 27580 8932 27636 12908
rect 27692 12740 27748 12750
rect 27692 12646 27748 12684
rect 28028 12068 28084 12078
rect 28028 9826 28084 12012
rect 28252 12066 28308 12078
rect 28252 12014 28254 12066
rect 28306 12014 28308 12066
rect 28252 11508 28308 12014
rect 28364 11732 28420 13356
rect 28476 13188 28532 13198
rect 28476 12962 28532 13132
rect 28476 12910 28478 12962
rect 28530 12910 28532 12962
rect 28476 12898 28532 12910
rect 28700 12740 28756 15372
rect 29036 14644 29092 16044
rect 29148 15986 29204 16718
rect 29436 16492 29700 16502
rect 29492 16436 29540 16492
rect 29596 16436 29644 16492
rect 29436 16426 29700 16436
rect 29372 16100 29428 16110
rect 29372 16006 29428 16044
rect 29148 15934 29150 15986
rect 29202 15934 29204 15986
rect 29148 15922 29204 15934
rect 29260 15764 29316 15774
rect 29148 15540 29204 15550
rect 29260 15540 29316 15708
rect 29148 15538 29316 15540
rect 29148 15486 29150 15538
rect 29202 15486 29316 15538
rect 29148 15484 29316 15486
rect 29148 15474 29204 15484
rect 29596 15316 29652 15326
rect 29260 15314 29652 15316
rect 29260 15262 29598 15314
rect 29650 15262 29652 15314
rect 29260 15260 29652 15262
rect 29148 14644 29204 14654
rect 29036 14642 29204 14644
rect 29036 14590 29150 14642
rect 29202 14590 29204 14642
rect 29036 14588 29204 14590
rect 29148 14578 29204 14588
rect 29036 14308 29092 14318
rect 28924 13858 28980 13870
rect 28924 13806 28926 13858
rect 28978 13806 28980 13858
rect 28924 13524 28980 13806
rect 28924 13458 28980 13468
rect 29036 13746 29092 14252
rect 29036 13694 29038 13746
rect 29090 13694 29092 13746
rect 29036 13186 29092 13694
rect 29036 13134 29038 13186
rect 29090 13134 29092 13186
rect 29036 13122 29092 13134
rect 29260 13188 29316 15260
rect 29596 15250 29652 15260
rect 29436 14924 29700 14934
rect 29492 14868 29540 14924
rect 29596 14868 29644 14924
rect 29436 14858 29700 14868
rect 29820 14532 29876 17052
rect 29932 16660 29988 18284
rect 30044 18274 30100 18284
rect 30268 18116 30324 18398
rect 30268 18050 30324 18060
rect 30380 18338 30436 18350
rect 30380 18286 30382 18338
rect 30434 18286 30436 18338
rect 30044 17668 30100 17678
rect 30044 16882 30100 17612
rect 30380 17220 30436 18286
rect 30604 17666 30660 19180
rect 30716 17778 30772 21422
rect 30828 19458 30884 22876
rect 30828 19406 30830 19458
rect 30882 19406 30884 19458
rect 30828 19394 30884 19406
rect 30940 22372 30996 22382
rect 30940 18676 30996 22316
rect 31052 22370 31108 24556
rect 31948 23940 32004 24556
rect 31948 23874 32004 23884
rect 31052 22318 31054 22370
rect 31106 22318 31108 22370
rect 31052 22306 31108 22318
rect 32060 21700 32116 21710
rect 31612 21698 32116 21700
rect 31612 21646 32062 21698
rect 32114 21646 32116 21698
rect 31612 21644 32116 21646
rect 31052 20356 31108 20366
rect 31108 20300 31220 20356
rect 31052 20290 31108 20300
rect 31052 20020 31108 20030
rect 31052 19926 31108 19964
rect 30716 17726 30718 17778
rect 30770 17726 30772 17778
rect 30716 17714 30772 17726
rect 30828 18620 30996 18676
rect 30604 17614 30606 17666
rect 30658 17614 30660 17666
rect 30604 17602 30660 17614
rect 30492 17220 30548 17230
rect 30380 17164 30492 17220
rect 30492 17154 30548 17164
rect 30268 16996 30324 17006
rect 30268 16994 30436 16996
rect 30268 16942 30270 16994
rect 30322 16942 30436 16994
rect 30268 16940 30436 16942
rect 30268 16930 30324 16940
rect 30044 16830 30046 16882
rect 30098 16830 30100 16882
rect 30044 16818 30100 16830
rect 30268 16772 30324 16782
rect 30268 16678 30324 16716
rect 29932 16604 30100 16660
rect 29932 15874 29988 15886
rect 29932 15822 29934 15874
rect 29986 15822 29988 15874
rect 29932 15540 29988 15822
rect 29932 15474 29988 15484
rect 29596 14476 29876 14532
rect 29596 13860 29652 14476
rect 29708 14308 29764 14318
rect 29708 14214 29764 14252
rect 29820 14196 29876 14206
rect 29820 13972 29876 14140
rect 30044 14196 30100 16604
rect 30268 16098 30324 16110
rect 30268 16046 30270 16098
rect 30322 16046 30324 16098
rect 30268 15652 30324 16046
rect 30268 15586 30324 15596
rect 30380 15428 30436 16940
rect 30828 16772 30884 18620
rect 30940 18452 30996 18462
rect 30940 18358 30996 18396
rect 30268 15372 30436 15428
rect 30492 16716 30884 16772
rect 31052 18340 31108 18350
rect 30268 14868 30324 15372
rect 30380 15204 30436 15242
rect 30380 15138 30436 15148
rect 30044 14130 30100 14140
rect 30156 14812 30324 14868
rect 30044 13972 30100 13982
rect 29820 13970 30100 13972
rect 29820 13918 30046 13970
rect 30098 13918 30100 13970
rect 29820 13916 30100 13918
rect 30044 13906 30100 13916
rect 29596 13804 29988 13860
rect 29596 13636 29652 13646
rect 29596 13542 29652 13580
rect 29820 13524 29876 13534
rect 29436 13356 29700 13366
rect 29492 13300 29540 13356
rect 29596 13300 29644 13356
rect 29436 13290 29700 13300
rect 29484 13188 29540 13198
rect 29260 13132 29428 13188
rect 29260 12850 29316 12862
rect 29260 12798 29262 12850
rect 29314 12798 29316 12850
rect 29148 12740 29204 12750
rect 29260 12740 29316 12798
rect 28700 12516 28756 12684
rect 28700 12450 28756 12460
rect 28812 12684 29148 12740
rect 29204 12684 29316 12740
rect 28588 12180 28644 12190
rect 28588 12178 28756 12180
rect 28588 12126 28590 12178
rect 28642 12126 28756 12178
rect 28588 12124 28756 12126
rect 28588 12114 28644 12124
rect 28588 11956 28644 11966
rect 28364 11676 28532 11732
rect 28140 11452 28252 11508
rect 28140 10052 28196 11452
rect 28252 11442 28308 11452
rect 28364 11284 28420 11294
rect 28252 11172 28308 11182
rect 28252 11078 28308 11116
rect 28140 9996 28308 10052
rect 28028 9774 28030 9826
rect 28082 9774 28084 9826
rect 28028 9762 28084 9774
rect 28140 9828 28196 9838
rect 28140 9734 28196 9772
rect 27244 8094 27246 8146
rect 27298 8094 27300 8146
rect 27244 8082 27300 8094
rect 27468 8876 27636 8932
rect 28028 9156 28084 9166
rect 27356 8034 27412 8046
rect 27356 7982 27358 8034
rect 27410 7982 27412 8034
rect 27356 7924 27412 7982
rect 27132 7868 27412 7924
rect 26796 7700 26852 7710
rect 26852 7644 27188 7700
rect 26796 7634 26852 7644
rect 26684 7588 26740 7598
rect 26684 7494 26740 7532
rect 26908 7476 26964 7486
rect 26460 7364 26516 7374
rect 26460 7362 26628 7364
rect 26460 7310 26462 7362
rect 26514 7310 26628 7362
rect 26460 7308 26628 7310
rect 26460 7298 26516 7308
rect 26460 6916 26516 6926
rect 26012 6748 26292 6804
rect 25676 6692 25732 6702
rect 25676 6598 25732 6636
rect 25564 6402 25620 6412
rect 26012 6466 26068 6478
rect 26012 6414 26014 6466
rect 26066 6414 26068 6466
rect 25404 6300 25668 6310
rect 25460 6244 25508 6300
rect 25564 6244 25612 6300
rect 25404 6234 25668 6244
rect 26012 6132 26068 6414
rect 26236 6356 26292 6748
rect 26348 6692 26404 6702
rect 26348 6598 26404 6636
rect 26236 6300 26404 6356
rect 26124 6132 26180 6142
rect 25228 6076 25620 6132
rect 25564 6018 25620 6076
rect 26068 6130 26180 6132
rect 26068 6078 26126 6130
rect 26178 6078 26180 6130
rect 26068 6076 26180 6078
rect 26012 6066 26068 6076
rect 26124 6066 26180 6076
rect 26348 6132 26404 6300
rect 26348 6066 26404 6076
rect 25564 5966 25566 6018
rect 25618 5966 25620 6018
rect 25564 5954 25620 5966
rect 25228 5906 25284 5918
rect 25228 5854 25230 5906
rect 25282 5854 25284 5906
rect 25228 5684 25284 5854
rect 25340 5908 25396 5946
rect 25340 5842 25396 5852
rect 25676 5908 25732 5918
rect 25228 5628 25508 5684
rect 25452 5234 25508 5628
rect 25452 5182 25454 5234
rect 25506 5182 25508 5234
rect 25452 5170 25508 5182
rect 25340 5124 25396 5134
rect 25340 5030 25396 5068
rect 25676 5012 25732 5852
rect 25788 5908 25844 5918
rect 26236 5908 26292 5918
rect 25788 5906 26292 5908
rect 25788 5854 25790 5906
rect 25842 5854 26238 5906
rect 26290 5854 26292 5906
rect 25788 5852 26292 5854
rect 25788 5842 25844 5852
rect 26236 5842 26292 5852
rect 26348 5908 26404 5918
rect 26348 5814 26404 5852
rect 26460 5684 26516 6860
rect 26236 5628 26516 5684
rect 26012 5180 26180 5236
rect 26012 5122 26068 5180
rect 26012 5070 26014 5122
rect 26066 5070 26068 5122
rect 26012 5058 26068 5070
rect 26124 5122 26180 5180
rect 26124 5070 26126 5122
rect 26178 5070 26180 5122
rect 26124 5058 26180 5070
rect 25676 4956 25956 5012
rect 25564 4900 25620 4938
rect 25564 4834 25620 4844
rect 25404 4732 25668 4742
rect 25460 4676 25508 4732
rect 25564 4676 25612 4732
rect 25404 4666 25668 4676
rect 25340 4564 25396 4574
rect 25340 4338 25396 4508
rect 25900 4452 25956 4956
rect 26012 4452 26068 4462
rect 25900 4450 26068 4452
rect 25900 4398 26014 4450
rect 26066 4398 26068 4450
rect 25900 4396 26068 4398
rect 26236 4452 26292 5628
rect 26460 5460 26516 5470
rect 26348 5348 26404 5358
rect 26348 5010 26404 5292
rect 26460 5122 26516 5404
rect 26460 5070 26462 5122
rect 26514 5070 26516 5122
rect 26460 5058 26516 5070
rect 26348 4958 26350 5010
rect 26402 4958 26404 5010
rect 26348 4946 26404 4958
rect 26236 4396 26404 4452
rect 26012 4386 26068 4396
rect 25340 4286 25342 4338
rect 25394 4286 25396 4338
rect 25340 4274 25396 4286
rect 25564 4340 25620 4350
rect 25564 3666 25620 4284
rect 26348 4340 26404 4396
rect 26348 4274 26404 4284
rect 25564 3614 25566 3666
rect 25618 3614 25620 3666
rect 25564 3602 25620 3614
rect 26236 4228 26292 4238
rect 25900 3444 25956 3482
rect 25900 3378 25956 3388
rect 26236 3442 26292 4172
rect 26572 3668 26628 7308
rect 26796 6804 26852 6814
rect 26796 6580 26852 6748
rect 26908 6692 26964 7420
rect 27020 7474 27076 7486
rect 27020 7422 27022 7474
rect 27074 7422 27076 7474
rect 27020 7028 27076 7422
rect 27132 7476 27188 7644
rect 27132 7410 27188 7420
rect 27468 7698 27524 8876
rect 28028 8258 28084 9100
rect 28028 8206 28030 8258
rect 28082 8206 28084 8258
rect 28028 8194 28084 8206
rect 28140 8260 28196 8270
rect 28140 8166 28196 8204
rect 28252 8258 28308 9996
rect 28364 9938 28420 11228
rect 28364 9886 28366 9938
rect 28418 9886 28420 9938
rect 28364 9874 28420 9886
rect 28252 8206 28254 8258
rect 28306 8206 28308 8258
rect 28252 8194 28308 8206
rect 27692 8146 27748 8158
rect 27692 8094 27694 8146
rect 27746 8094 27748 8146
rect 27468 7646 27470 7698
rect 27522 7646 27524 7698
rect 27020 6962 27076 6972
rect 27132 6692 27188 6702
rect 27468 6692 27524 7646
rect 26908 6636 27076 6692
rect 26796 6578 26964 6580
rect 26796 6526 26798 6578
rect 26850 6526 26964 6578
rect 26796 6524 26964 6526
rect 26796 6486 26852 6524
rect 26684 6468 26740 6478
rect 26684 5906 26740 6412
rect 26684 5854 26686 5906
rect 26738 5854 26740 5906
rect 26684 5842 26740 5854
rect 26796 6132 26852 6142
rect 26796 5572 26852 6076
rect 26684 5516 26852 5572
rect 26908 6020 26964 6524
rect 27020 6244 27076 6636
rect 27132 6690 27524 6692
rect 27132 6638 27134 6690
rect 27186 6638 27524 6690
rect 27132 6636 27524 6638
rect 27132 6626 27188 6636
rect 27468 6578 27524 6636
rect 27468 6526 27470 6578
rect 27522 6526 27524 6578
rect 27468 6514 27524 6526
rect 27580 8034 27636 8046
rect 27580 7982 27582 8034
rect 27634 7982 27636 8034
rect 27580 6356 27636 7982
rect 27692 7476 27748 8094
rect 28364 7700 28420 7710
rect 28476 7700 28532 11676
rect 28588 11282 28644 11900
rect 28588 11230 28590 11282
rect 28642 11230 28644 11282
rect 28588 11218 28644 11230
rect 28700 10388 28756 12124
rect 28700 10322 28756 10332
rect 28812 10836 28868 12684
rect 29148 12674 29204 12684
rect 29372 12628 29428 13132
rect 29484 13186 29764 13188
rect 29484 13134 29486 13186
rect 29538 13134 29764 13186
rect 29484 13132 29764 13134
rect 29484 13122 29540 13132
rect 29708 13074 29764 13132
rect 29708 13022 29710 13074
rect 29762 13022 29764 13074
rect 29708 13010 29764 13022
rect 29260 12572 29428 12628
rect 29596 12964 29652 12974
rect 28924 12180 28980 12190
rect 28924 12086 28980 12124
rect 29148 12178 29204 12190
rect 29148 12126 29150 12178
rect 29202 12126 29204 12178
rect 29036 12068 29092 12078
rect 29036 11974 29092 12012
rect 28812 10164 28868 10780
rect 28700 10108 28868 10164
rect 28588 9826 28644 9838
rect 28588 9774 28590 9826
rect 28642 9774 28644 9826
rect 28588 9268 28644 9774
rect 28588 9202 28644 9212
rect 28700 9044 28756 10108
rect 29148 10052 29204 12126
rect 29260 11620 29316 12572
rect 29596 12066 29652 12908
rect 29596 12014 29598 12066
rect 29650 12014 29652 12066
rect 29596 12002 29652 12014
rect 29436 11788 29700 11798
rect 29492 11732 29540 11788
rect 29596 11732 29644 11788
rect 29436 11722 29700 11732
rect 29260 11564 29428 11620
rect 29260 11394 29316 11406
rect 29260 11342 29262 11394
rect 29314 11342 29316 11394
rect 29260 10500 29316 11342
rect 29372 11172 29428 11564
rect 29372 11106 29428 11116
rect 29260 10434 29316 10444
rect 29436 10220 29700 10230
rect 29492 10164 29540 10220
rect 29596 10164 29644 10220
rect 29436 10154 29700 10164
rect 29820 10108 29876 13468
rect 29932 11508 29988 13804
rect 30156 13188 30212 14812
rect 30268 14642 30324 14654
rect 30268 14590 30270 14642
rect 30322 14590 30324 14642
rect 30268 13748 30324 14590
rect 30380 13748 30436 13758
rect 30268 13746 30436 13748
rect 30268 13694 30382 13746
rect 30434 13694 30436 13746
rect 30268 13692 30436 13694
rect 30380 13682 30436 13692
rect 30156 13122 30212 13132
rect 30156 12962 30212 12974
rect 30156 12910 30158 12962
rect 30210 12910 30212 12962
rect 30156 12852 30212 12910
rect 29932 11442 29988 11452
rect 30044 12516 30100 12526
rect 29932 11284 29988 11294
rect 29932 11190 29988 11228
rect 29820 10052 29988 10108
rect 29148 9826 29204 9996
rect 29148 9774 29150 9826
rect 29202 9774 29204 9826
rect 29148 9762 29204 9774
rect 29260 9716 29316 9726
rect 29260 9622 29316 9660
rect 29372 9602 29428 9614
rect 29372 9550 29374 9602
rect 29426 9550 29428 9602
rect 29260 9268 29316 9278
rect 29260 9174 29316 9212
rect 29372 9266 29428 9550
rect 29596 9604 29652 9614
rect 29596 9510 29652 9548
rect 29372 9214 29374 9266
rect 29426 9214 29428 9266
rect 29148 9156 29204 9166
rect 29148 9062 29204 9100
rect 28588 8988 28756 9044
rect 28588 8036 28644 8988
rect 28812 8930 28868 8942
rect 28812 8878 28814 8930
rect 28866 8878 28868 8930
rect 28812 8820 28868 8878
rect 29372 8820 29428 9214
rect 28812 8764 29428 8820
rect 29820 9042 29876 9054
rect 29820 8990 29822 9042
rect 29874 8990 29876 9042
rect 29436 8652 29700 8662
rect 29492 8596 29540 8652
rect 29596 8596 29644 8652
rect 29436 8586 29700 8596
rect 29484 8484 29540 8494
rect 28700 8260 28756 8270
rect 28700 8258 29316 8260
rect 28700 8206 28702 8258
rect 28754 8206 29316 8258
rect 28700 8204 29316 8206
rect 28700 8194 28756 8204
rect 28588 7970 28644 7980
rect 29148 8034 29204 8046
rect 29148 7982 29150 8034
rect 29202 7982 29204 8034
rect 28364 7698 28532 7700
rect 28364 7646 28366 7698
rect 28418 7646 28532 7698
rect 28364 7644 28532 7646
rect 29148 7700 29204 7982
rect 29260 7812 29316 8204
rect 29484 8146 29540 8428
rect 29484 8094 29486 8146
rect 29538 8094 29540 8146
rect 29484 8082 29540 8094
rect 29260 7756 29652 7812
rect 28364 7634 28420 7644
rect 29148 7634 29204 7644
rect 29596 7698 29652 7756
rect 29596 7646 29598 7698
rect 29650 7646 29652 7698
rect 29596 7634 29652 7646
rect 27804 7586 27860 7598
rect 27804 7534 27806 7586
rect 27858 7534 27860 7586
rect 27804 7476 27860 7534
rect 28588 7588 28644 7598
rect 28588 7494 28644 7532
rect 28924 7588 28980 7598
rect 27804 7420 28196 7476
rect 27692 7410 27748 7420
rect 27692 7028 27748 7038
rect 27748 6972 27860 7028
rect 27692 6962 27748 6972
rect 27580 6290 27636 6300
rect 27804 6578 27860 6972
rect 27804 6526 27806 6578
rect 27858 6526 27860 6578
rect 27020 6188 27412 6244
rect 27356 6130 27412 6188
rect 27356 6078 27358 6130
rect 27410 6078 27412 6130
rect 27244 6020 27300 6030
rect 26908 6018 27300 6020
rect 26908 5966 27246 6018
rect 27298 5966 27300 6018
rect 26908 5964 27300 5966
rect 26684 4564 26740 5516
rect 26908 5460 26964 5964
rect 27244 5954 27300 5964
rect 26908 5394 26964 5404
rect 26796 5348 26852 5358
rect 26796 5254 26852 5292
rect 27356 5348 27412 6078
rect 27804 6020 27860 6526
rect 28140 6804 28196 7420
rect 28252 7028 28308 7038
rect 28308 6972 28420 7028
rect 28252 6962 28308 6972
rect 27916 6020 27972 6030
rect 27804 6018 27972 6020
rect 27804 5966 27918 6018
rect 27970 5966 27972 6018
rect 27804 5964 27972 5966
rect 27916 5954 27972 5964
rect 28028 6018 28084 6030
rect 28028 5966 28030 6018
rect 28082 5966 28084 6018
rect 27356 5282 27412 5292
rect 27580 5906 27636 5918
rect 27580 5854 27582 5906
rect 27634 5854 27636 5906
rect 27580 5122 27636 5854
rect 27692 5908 27748 5918
rect 27748 5852 27860 5908
rect 27692 5842 27748 5852
rect 27580 5070 27582 5122
rect 27634 5070 27636 5122
rect 27580 5058 27636 5070
rect 26684 4498 26740 4508
rect 26908 5010 26964 5022
rect 26908 4958 26910 5010
rect 26962 4958 26964 5010
rect 26908 3778 26964 4958
rect 27804 5012 27860 5852
rect 28028 5684 28084 5966
rect 28028 5618 28084 5628
rect 28028 5124 28084 5134
rect 28028 5030 28084 5068
rect 28140 5122 28196 6748
rect 28364 6690 28420 6972
rect 28364 6638 28366 6690
rect 28418 6638 28420 6690
rect 28252 6132 28308 6142
rect 28252 6038 28308 6076
rect 28364 6020 28420 6638
rect 28700 6916 28756 6926
rect 28700 6690 28756 6860
rect 28700 6638 28702 6690
rect 28754 6638 28756 6690
rect 28700 6626 28756 6638
rect 28476 6466 28532 6478
rect 28476 6414 28478 6466
rect 28530 6414 28532 6466
rect 28476 6244 28532 6414
rect 28476 6178 28532 6188
rect 28588 6356 28644 6366
rect 28476 6020 28532 6030
rect 28364 6018 28532 6020
rect 28364 5966 28478 6018
rect 28530 5966 28532 6018
rect 28364 5964 28532 5966
rect 28476 5954 28532 5964
rect 28588 6018 28644 6300
rect 28588 5966 28590 6018
rect 28642 5966 28644 6018
rect 28364 5348 28420 5358
rect 28588 5348 28644 5966
rect 28812 5908 28868 5918
rect 28812 5814 28868 5852
rect 28420 5292 28532 5348
rect 28364 5282 28420 5292
rect 28476 5234 28532 5292
rect 28924 5348 28980 7532
rect 29372 7588 29428 7598
rect 29372 7586 29540 7588
rect 29372 7534 29374 7586
rect 29426 7534 29540 7586
rect 29372 7532 29540 7534
rect 29372 7522 29428 7532
rect 29148 7476 29204 7486
rect 29260 7476 29316 7486
rect 29204 7474 29316 7476
rect 29204 7422 29262 7474
rect 29314 7422 29316 7474
rect 29204 7420 29316 7422
rect 29148 7252 29204 7420
rect 29260 7410 29316 7420
rect 29484 7252 29540 7532
rect 29036 7196 29204 7252
rect 29260 7196 29540 7252
rect 29036 6018 29092 7196
rect 29148 6244 29204 6254
rect 29148 6130 29204 6188
rect 29148 6078 29150 6130
rect 29202 6078 29204 6130
rect 29148 6066 29204 6078
rect 29036 5966 29038 6018
rect 29090 5966 29092 6018
rect 29036 5954 29092 5966
rect 29260 5684 29316 7196
rect 29436 7084 29700 7094
rect 29492 7028 29540 7084
rect 29596 7028 29644 7084
rect 29436 7018 29700 7028
rect 29820 6916 29876 8990
rect 29372 6860 29876 6916
rect 29372 6130 29428 6860
rect 29932 6804 29988 10052
rect 30044 8370 30100 12460
rect 30156 11956 30212 12796
rect 30156 11890 30212 11900
rect 30044 8318 30046 8370
rect 30098 8318 30100 8370
rect 30044 8306 30100 8318
rect 30156 11172 30212 11182
rect 30044 7700 30100 7710
rect 30156 7700 30212 11116
rect 30492 10164 30548 16716
rect 31052 16212 31108 18284
rect 31164 18228 31220 20300
rect 31500 20132 31556 20142
rect 31500 20018 31556 20076
rect 31500 19966 31502 20018
rect 31554 19966 31556 20018
rect 31500 19954 31556 19966
rect 31612 19460 31668 21644
rect 32060 21634 32116 21644
rect 31612 19394 31668 19404
rect 31724 21474 31780 21486
rect 31724 21422 31726 21474
rect 31778 21422 31780 21474
rect 31276 18788 31332 18798
rect 31332 18732 31668 18788
rect 31276 18722 31332 18732
rect 31500 18450 31556 18462
rect 31500 18398 31502 18450
rect 31554 18398 31556 18450
rect 31164 18172 31444 18228
rect 31276 17666 31332 17678
rect 31276 17614 31278 17666
rect 31330 17614 31332 17666
rect 31164 17220 31220 17230
rect 31164 16882 31220 17164
rect 31276 16994 31332 17614
rect 31276 16942 31278 16994
rect 31330 16942 31332 16994
rect 31276 16930 31332 16942
rect 31164 16830 31166 16882
rect 31218 16830 31220 16882
rect 31164 16818 31220 16830
rect 31388 16882 31444 18172
rect 31500 17892 31556 18398
rect 31500 17826 31556 17836
rect 31388 16830 31390 16882
rect 31442 16830 31444 16882
rect 31388 16818 31444 16830
rect 31500 17666 31556 17678
rect 31500 17614 31502 17666
rect 31554 17614 31556 17666
rect 31500 16884 31556 17614
rect 31500 16818 31556 16828
rect 31500 16212 31556 16222
rect 31052 16210 31556 16212
rect 31052 16158 31502 16210
rect 31554 16158 31556 16210
rect 31052 16156 31556 16158
rect 31500 16146 31556 16156
rect 30604 15986 30660 15998
rect 30604 15934 30606 15986
rect 30658 15934 30660 15986
rect 30604 14308 30660 15934
rect 30828 15986 30884 15998
rect 30828 15934 30830 15986
rect 30882 15934 30884 15986
rect 30828 15204 30884 15934
rect 30828 15138 30884 15148
rect 30604 13858 30660 14252
rect 30604 13806 30606 13858
rect 30658 13806 30660 13858
rect 30604 13794 30660 13806
rect 31164 14084 31220 14094
rect 31164 13858 31220 14028
rect 31164 13806 31166 13858
rect 31218 13806 31220 13858
rect 31164 13794 31220 13806
rect 31612 13858 31668 18732
rect 31724 18562 31780 21422
rect 31836 21362 31892 21374
rect 31836 21310 31838 21362
rect 31890 21310 31892 21362
rect 31836 20130 31892 21310
rect 32060 20802 32116 20814
rect 32060 20750 32062 20802
rect 32114 20750 32116 20802
rect 32060 20244 32116 20750
rect 32172 20580 32228 26238
rect 33068 27300 33124 27310
rect 33068 27188 33124 27244
rect 33180 27188 33236 27198
rect 33068 27186 33236 27188
rect 33068 27134 33182 27186
rect 33234 27134 33236 27186
rect 33068 27132 33236 27134
rect 33068 24836 33124 27132
rect 33180 27122 33236 27132
rect 33180 26180 33236 26190
rect 33180 26086 33236 26124
rect 33180 25620 33236 25630
rect 33180 25526 33236 25564
rect 33180 24836 33236 24846
rect 33068 24834 33236 24836
rect 33068 24782 33182 24834
rect 33234 24782 33236 24834
rect 33068 24780 33236 24782
rect 33180 24770 33236 24780
rect 32508 24724 32564 24734
rect 32508 24630 32564 24668
rect 33068 24500 33124 24510
rect 32172 20514 32228 20524
rect 32284 24498 33124 24500
rect 32284 24446 33070 24498
rect 33122 24446 33124 24498
rect 32284 24444 33124 24446
rect 32060 20178 32116 20188
rect 31836 20078 31838 20130
rect 31890 20078 31892 20130
rect 31836 20066 31892 20078
rect 32172 20130 32228 20142
rect 32172 20078 32174 20130
rect 32226 20078 32228 20130
rect 32172 19908 32228 20078
rect 31724 18510 31726 18562
rect 31778 18510 31780 18562
rect 31724 18498 31780 18510
rect 32060 18900 32116 18910
rect 31724 18116 31780 18126
rect 31780 18060 31892 18116
rect 31724 18050 31780 18060
rect 31724 17890 31780 17902
rect 31724 17838 31726 17890
rect 31778 17838 31780 17890
rect 31724 14532 31780 17838
rect 31724 14466 31780 14476
rect 31724 13972 31780 13982
rect 31724 13878 31780 13916
rect 31612 13806 31614 13858
rect 31666 13806 31668 13858
rect 31612 13794 31668 13806
rect 30828 13748 30884 13758
rect 30268 10108 30492 10164
rect 30268 9938 30324 10108
rect 30492 10070 30548 10108
rect 30604 13636 30660 13646
rect 30268 9886 30270 9938
rect 30322 9886 30324 9938
rect 30268 9874 30324 9886
rect 30268 9268 30324 9278
rect 30604 9268 30660 13580
rect 30716 13076 30772 13086
rect 30716 12982 30772 13020
rect 30268 9266 30660 9268
rect 30268 9214 30270 9266
rect 30322 9214 30660 9266
rect 30268 9212 30660 9214
rect 30716 12628 30772 12638
rect 30268 9202 30324 9212
rect 30604 9044 30660 9054
rect 30716 9044 30772 12572
rect 30604 9042 30772 9044
rect 30604 8990 30606 9042
rect 30658 8990 30772 9042
rect 30604 8988 30772 8990
rect 30604 8978 30660 8988
rect 30828 8820 30884 13692
rect 31724 13524 31780 13534
rect 31836 13524 31892 18060
rect 32060 17556 32116 18844
rect 32172 18676 32228 19852
rect 32172 18562 32228 18620
rect 32172 18510 32174 18562
rect 32226 18510 32228 18562
rect 32172 18498 32228 18510
rect 32284 18450 32340 24444
rect 33068 24434 33124 24444
rect 33180 24500 33236 24510
rect 32732 23940 32788 23950
rect 32732 23826 32788 23884
rect 33180 23938 33236 24444
rect 33180 23886 33182 23938
rect 33234 23886 33236 23938
rect 33180 23874 33236 23886
rect 32732 23774 32734 23826
rect 32786 23774 32788 23826
rect 32620 23716 32676 23726
rect 32396 23714 32676 23716
rect 32396 23662 32622 23714
rect 32674 23662 32676 23714
rect 32396 23660 32676 23662
rect 32396 21476 32452 23660
rect 32620 23650 32676 23660
rect 32620 22932 32676 22942
rect 32396 21410 32452 21420
rect 32508 22876 32620 22932
rect 32396 20692 32452 20702
rect 32396 20598 32452 20636
rect 32508 20018 32564 22876
rect 32620 22866 32676 22876
rect 32508 19966 32510 20018
rect 32562 19966 32564 20018
rect 32508 19954 32564 19966
rect 32620 21924 32676 21934
rect 32284 18398 32286 18450
rect 32338 18398 32340 18450
rect 32284 18386 32340 18398
rect 32508 18452 32564 18462
rect 32508 17892 32564 18396
rect 31948 16996 32004 17006
rect 31948 16098 32004 16940
rect 32060 16882 32116 17500
rect 32060 16830 32062 16882
rect 32114 16830 32116 16882
rect 32060 16818 32116 16830
rect 32172 17836 32564 17892
rect 31948 16046 31950 16098
rect 32002 16046 32004 16098
rect 31948 16034 32004 16046
rect 32172 13970 32228 17836
rect 32620 16210 32676 21868
rect 32732 20690 32788 23774
rect 32956 23714 33012 23726
rect 32956 23662 32958 23714
rect 33010 23662 33012 23714
rect 32956 22820 33012 23662
rect 33180 23268 33236 23278
rect 33180 23174 33236 23212
rect 33068 22932 33124 22942
rect 33068 22838 33124 22876
rect 32732 20638 32734 20690
rect 32786 20638 32788 20690
rect 32732 20132 32788 20638
rect 32732 20066 32788 20076
rect 32844 22764 33012 22820
rect 32732 19908 32788 19918
rect 32844 19908 32900 22764
rect 32956 22596 33012 22606
rect 33292 22596 33348 30940
rect 33468 29820 33732 29830
rect 33524 29764 33572 29820
rect 33628 29764 33676 29820
rect 33468 29754 33732 29764
rect 34076 28644 34132 34200
rect 34076 28578 34132 28588
rect 33468 28252 33732 28262
rect 33524 28196 33572 28252
rect 33628 28196 33676 28252
rect 33468 28186 33732 28196
rect 33468 26684 33732 26694
rect 33524 26628 33572 26684
rect 33628 26628 33676 26684
rect 33468 26618 33732 26628
rect 33852 26180 33908 26190
rect 33468 25116 33732 25126
rect 33524 25060 33572 25116
rect 33628 25060 33676 25116
rect 33468 25050 33732 25060
rect 33468 23548 33732 23558
rect 33524 23492 33572 23548
rect 33628 23492 33676 23548
rect 33468 23482 33732 23492
rect 32956 22594 33348 22596
rect 32956 22542 32958 22594
rect 33010 22542 33348 22594
rect 32956 22540 33348 22542
rect 32956 22530 33012 22540
rect 33852 22148 33908 26124
rect 33292 22092 33908 22148
rect 33964 24724 34020 24734
rect 33180 21474 33236 21486
rect 33180 21422 33182 21474
rect 33234 21422 33236 21474
rect 32788 19852 32900 19908
rect 32956 20580 33012 20590
rect 32732 19842 32788 19852
rect 32844 19348 32900 19358
rect 32956 19348 33012 20524
rect 33180 20468 33236 21422
rect 33292 20914 33348 22092
rect 33468 21980 33732 21990
rect 33524 21924 33572 21980
rect 33628 21924 33676 21980
rect 33468 21914 33732 21924
rect 33292 20862 33294 20914
rect 33346 20862 33348 20914
rect 33292 20850 33348 20862
rect 33180 20188 33236 20412
rect 33468 20412 33732 20422
rect 33524 20356 33572 20412
rect 33628 20356 33676 20412
rect 33468 20346 33732 20356
rect 33180 20132 33348 20188
rect 33180 20018 33236 20030
rect 33180 19966 33182 20018
rect 33234 19966 33236 20018
rect 33068 19794 33124 19806
rect 33068 19742 33070 19794
rect 33122 19742 33124 19794
rect 33068 19460 33124 19742
rect 33180 19684 33236 19966
rect 33180 19618 33236 19628
rect 33068 19394 33124 19404
rect 32844 19346 33012 19348
rect 32844 19294 32846 19346
rect 32898 19294 33012 19346
rect 32844 19292 33012 19294
rect 32844 19282 32900 19292
rect 33068 19236 33124 19246
rect 33068 18674 33124 19180
rect 33068 18622 33070 18674
rect 33122 18622 33124 18674
rect 33068 18610 33124 18622
rect 33292 18452 33348 20132
rect 33852 19236 33908 19246
rect 33964 19236 34020 24668
rect 33908 19180 34020 19236
rect 33852 19170 33908 19180
rect 33468 18844 33732 18854
rect 33524 18788 33572 18844
rect 33628 18788 33676 18844
rect 33468 18778 33732 18788
rect 33292 18386 33348 18396
rect 33180 18340 33236 18350
rect 32620 16158 32622 16210
rect 32674 16158 32676 16210
rect 32620 16146 32676 16158
rect 32732 18338 33236 18340
rect 32732 18286 33182 18338
rect 33234 18286 33236 18338
rect 32732 18284 33236 18286
rect 32732 15988 32788 18284
rect 33180 18274 33236 18284
rect 32956 17556 33012 17566
rect 33012 17500 33124 17556
rect 32956 17490 33012 17500
rect 33068 17442 33124 17500
rect 33068 17390 33070 17442
rect 33122 17390 33124 17442
rect 33068 17378 33124 17390
rect 33180 17554 33236 17566
rect 33180 17502 33182 17554
rect 33234 17502 33236 17554
rect 33180 16996 33236 17502
rect 33468 17276 33732 17286
rect 33524 17220 33572 17276
rect 33628 17220 33676 17276
rect 33468 17210 33732 17220
rect 33236 16940 33348 16996
rect 33180 16902 33236 16940
rect 32956 16100 33012 16110
rect 32956 16006 33012 16044
rect 32172 13918 32174 13970
rect 32226 13918 32228 13970
rect 32172 13906 32228 13918
rect 32284 15932 32788 15988
rect 31724 13522 31892 13524
rect 31724 13470 31726 13522
rect 31778 13470 31892 13522
rect 31724 13468 31892 13470
rect 31724 13458 31780 13468
rect 31052 12964 31108 12974
rect 31052 12870 31108 12908
rect 31276 12852 31332 12862
rect 31276 12758 31332 12796
rect 31724 12850 31780 12862
rect 31724 12798 31726 12850
rect 31778 12798 31780 12850
rect 31724 12066 31780 12798
rect 32284 12628 32340 15932
rect 32508 15652 32564 15662
rect 32508 15202 32564 15596
rect 33180 15428 33236 15438
rect 33180 15334 33236 15372
rect 32508 15150 32510 15202
rect 32562 15150 32564 15202
rect 32508 15138 32564 15150
rect 33068 14532 33124 14542
rect 32956 14530 33124 14532
rect 32956 14478 33070 14530
rect 33122 14478 33124 14530
rect 32956 14476 33124 14478
rect 32396 14418 32452 14430
rect 32396 14366 32398 14418
rect 32450 14366 32452 14418
rect 32396 14084 32452 14366
rect 32396 13972 32452 14028
rect 32396 13916 32676 13972
rect 32508 13746 32564 13758
rect 32508 13694 32510 13746
rect 32562 13694 32564 13746
rect 32396 13412 32452 13422
rect 32396 13074 32452 13356
rect 32396 13022 32398 13074
rect 32450 13022 32452 13074
rect 32396 13010 32452 13022
rect 32284 12562 32340 12572
rect 32396 12852 32452 12862
rect 31724 12014 31726 12066
rect 31778 12014 31780 12066
rect 31724 11788 31780 12014
rect 32060 12180 32116 12190
rect 31724 11732 32004 11788
rect 31836 10612 31892 10622
rect 31724 10500 31780 10510
rect 31724 10406 31780 10444
rect 31052 10164 31108 10174
rect 31108 10108 31332 10164
rect 31052 10098 31108 10108
rect 31276 9266 31332 10108
rect 31836 9492 31892 10556
rect 31836 9426 31892 9436
rect 31276 9214 31278 9266
rect 31330 9214 31332 9266
rect 31276 9202 31332 9214
rect 31388 9268 31444 9278
rect 31948 9268 32004 11732
rect 32060 11506 32116 12124
rect 32396 12178 32452 12796
rect 32396 12126 32398 12178
rect 32450 12126 32452 12178
rect 32396 12114 32452 12126
rect 32508 12740 32564 13694
rect 32060 11454 32062 11506
rect 32114 11454 32116 11506
rect 32060 11442 32116 11454
rect 32396 11284 32452 11294
rect 32508 11284 32564 12684
rect 32620 11844 32676 13916
rect 32732 12962 32788 12974
rect 32732 12910 32734 12962
rect 32786 12910 32788 12962
rect 32732 12740 32788 12910
rect 32956 12852 33012 14476
rect 33068 14466 33124 14476
rect 32956 12786 33012 12796
rect 33068 14196 33124 14206
rect 32732 12674 32788 12684
rect 33068 12402 33124 14140
rect 33180 13636 33236 13646
rect 33292 13636 33348 16940
rect 33468 15708 33732 15718
rect 33524 15652 33572 15708
rect 33628 15652 33676 15708
rect 33468 15642 33732 15652
rect 33468 14140 33732 14150
rect 33524 14084 33572 14140
rect 33628 14084 33676 14140
rect 33468 14074 33732 14084
rect 33180 13634 33348 13636
rect 33180 13582 33182 13634
rect 33234 13582 33348 13634
rect 33180 13580 33348 13582
rect 33180 13570 33236 13580
rect 33068 12350 33070 12402
rect 33122 12350 33124 12402
rect 33068 12338 33124 12350
rect 33180 12180 33236 12190
rect 33180 12086 33236 12124
rect 32620 11788 32900 11844
rect 32620 11396 32676 11406
rect 32620 11302 32676 11340
rect 32396 11282 32564 11284
rect 32396 11230 32398 11282
rect 32450 11230 32564 11282
rect 32396 11228 32564 11230
rect 32396 11218 32452 11228
rect 32396 9716 32452 9726
rect 32284 9714 32452 9716
rect 32284 9662 32398 9714
rect 32450 9662 32452 9714
rect 32284 9660 32452 9662
rect 31388 9266 31892 9268
rect 31388 9214 31390 9266
rect 31442 9214 31892 9266
rect 31388 9212 31892 9214
rect 31948 9212 32228 9268
rect 31388 9202 31444 9212
rect 31836 9154 31892 9212
rect 31836 9102 31838 9154
rect 31890 9102 31892 9154
rect 31836 9090 31892 9102
rect 30940 9044 30996 9054
rect 30940 8950 30996 8988
rect 31500 9044 31556 9054
rect 32060 9044 32116 9054
rect 31500 9042 31780 9044
rect 31500 8990 31502 9042
rect 31554 8990 31780 9042
rect 31500 8988 31780 8990
rect 31500 8978 31556 8988
rect 30380 8764 30884 8820
rect 30044 7698 30212 7700
rect 30044 7646 30046 7698
rect 30098 7646 30212 7698
rect 30044 7644 30212 7646
rect 30268 8370 30324 8382
rect 30268 8318 30270 8370
rect 30322 8318 30324 8370
rect 30268 7700 30324 8318
rect 30044 7634 30100 7644
rect 30268 7634 30324 7644
rect 30380 7586 30436 8764
rect 31612 8596 31668 8606
rect 31500 8540 31612 8596
rect 31052 7700 31108 7710
rect 31108 7644 31444 7700
rect 31052 7606 31108 7644
rect 30380 7534 30382 7586
rect 30434 7534 30436 7586
rect 30380 7522 30436 7534
rect 29484 6748 29988 6804
rect 30492 7476 30548 7486
rect 29484 6578 29540 6748
rect 30044 6690 30100 6702
rect 30044 6638 30046 6690
rect 30098 6638 30100 6690
rect 29484 6526 29486 6578
rect 29538 6526 29540 6578
rect 29484 6514 29540 6526
rect 29820 6580 29876 6590
rect 29820 6486 29876 6524
rect 29372 6078 29374 6130
rect 29426 6078 29428 6130
rect 29372 6066 29428 6078
rect 29596 6356 29652 6366
rect 29596 6130 29652 6300
rect 29596 6078 29598 6130
rect 29650 6078 29652 6130
rect 29596 6066 29652 6078
rect 30044 6132 30100 6638
rect 30492 6692 30548 7420
rect 30604 7474 30660 7486
rect 30604 7422 30606 7474
rect 30658 7422 30660 7474
rect 30604 6916 30660 7422
rect 31276 7474 31332 7486
rect 31276 7422 31278 7474
rect 31330 7422 31332 7474
rect 31164 7364 31220 7374
rect 31164 7270 31220 7308
rect 30604 6850 30660 6860
rect 30716 6804 30772 6814
rect 30604 6692 30660 6702
rect 30492 6690 30660 6692
rect 30492 6638 30606 6690
rect 30658 6638 30660 6690
rect 30492 6636 30660 6638
rect 30604 6626 30660 6636
rect 30716 6692 30772 6748
rect 31276 6692 31332 7422
rect 30716 6690 31332 6692
rect 30716 6638 30718 6690
rect 30770 6638 31332 6690
rect 30716 6636 31332 6638
rect 31388 6690 31444 7644
rect 31500 7364 31556 8540
rect 31612 8530 31668 8540
rect 31724 8484 31780 8988
rect 31500 7298 31556 7308
rect 31612 7474 31668 7486
rect 31612 7422 31614 7474
rect 31666 7422 31668 7474
rect 31500 6804 31556 6814
rect 31612 6804 31668 7422
rect 31500 6802 31668 6804
rect 31500 6750 31502 6802
rect 31554 6750 31668 6802
rect 31500 6748 31668 6750
rect 31500 6738 31556 6748
rect 31388 6638 31390 6690
rect 31442 6638 31444 6690
rect 30716 6626 30772 6636
rect 30044 6066 30100 6076
rect 30156 6468 30212 6478
rect 29820 6020 29876 6030
rect 29820 5926 29876 5964
rect 30156 5906 30212 6412
rect 30492 6466 30548 6478
rect 30492 6414 30494 6466
rect 30546 6414 30548 6466
rect 30492 6132 30548 6414
rect 30156 5854 30158 5906
rect 30210 5854 30212 5906
rect 30156 5842 30212 5854
rect 30380 5908 30436 5918
rect 30380 5814 30436 5852
rect 29708 5794 29764 5806
rect 29708 5742 29710 5794
rect 29762 5742 29764 5794
rect 29372 5684 29428 5694
rect 29260 5628 29372 5684
rect 29708 5684 29764 5742
rect 29708 5628 29876 5684
rect 29372 5618 29428 5628
rect 29436 5516 29700 5526
rect 29492 5460 29540 5516
rect 29596 5460 29644 5516
rect 29436 5450 29700 5460
rect 28924 5292 29428 5348
rect 28588 5282 28644 5292
rect 28476 5182 28478 5234
rect 28530 5182 28532 5234
rect 28476 5170 28532 5182
rect 28140 5070 28142 5122
rect 28194 5070 28196 5122
rect 28140 5058 28196 5070
rect 29036 5124 29092 5134
rect 29036 5030 29092 5068
rect 29372 5122 29428 5292
rect 29372 5070 29374 5122
rect 29426 5070 29428 5122
rect 29372 5058 29428 5070
rect 29708 5124 29764 5134
rect 29820 5124 29876 5628
rect 30268 5236 30324 5246
rect 30492 5236 30548 6076
rect 30828 6020 30884 6030
rect 30828 5906 30884 5964
rect 31052 6018 31108 6636
rect 31388 6626 31444 6638
rect 31612 6580 31668 6590
rect 31724 6580 31780 8428
rect 31948 9042 32116 9044
rect 31948 8990 32062 9042
rect 32114 8990 32116 9042
rect 31948 8988 32116 8990
rect 31948 7588 32004 8988
rect 32060 8978 32116 8988
rect 32060 7924 32116 7934
rect 32060 7698 32116 7868
rect 32060 7646 32062 7698
rect 32114 7646 32116 7698
rect 32060 7634 32116 7646
rect 32172 7700 32228 9212
rect 32284 9266 32340 9660
rect 32396 9650 32452 9660
rect 32284 9214 32286 9266
rect 32338 9214 32340 9266
rect 32284 9202 32340 9214
rect 32732 9492 32788 9502
rect 32508 9156 32564 9166
rect 32396 9042 32452 9054
rect 32396 8990 32398 9042
rect 32450 8990 32452 9042
rect 32396 8596 32452 8990
rect 32396 8530 32452 8540
rect 32396 8146 32452 8158
rect 32396 8094 32398 8146
rect 32450 8094 32452 8146
rect 32396 7924 32452 8094
rect 32396 7858 32452 7868
rect 32508 8148 32564 9100
rect 32172 7644 32340 7700
rect 31948 7476 32004 7532
rect 32172 7476 32228 7486
rect 31948 7474 32116 7476
rect 31948 7422 31950 7474
rect 32002 7422 32116 7474
rect 31948 7420 32116 7422
rect 31948 7410 32004 7420
rect 31612 6578 32004 6580
rect 31612 6526 31614 6578
rect 31666 6526 32004 6578
rect 31612 6524 32004 6526
rect 31612 6514 31668 6524
rect 31052 5966 31054 6018
rect 31106 5966 31108 6018
rect 31052 5954 31108 5966
rect 31164 6468 31220 6478
rect 30828 5854 30830 5906
rect 30882 5854 30884 5906
rect 30268 5234 30548 5236
rect 30268 5182 30270 5234
rect 30322 5182 30548 5234
rect 30268 5180 30548 5182
rect 30604 5796 30660 5806
rect 30268 5170 30324 5180
rect 29708 5122 29876 5124
rect 29708 5070 29710 5122
rect 29762 5070 29876 5122
rect 29708 5068 29876 5070
rect 29708 5058 29764 5068
rect 27916 5012 27972 5022
rect 27804 5010 27972 5012
rect 27804 4958 27918 5010
rect 27970 4958 27972 5010
rect 27804 4956 27972 4958
rect 27916 4228 27972 4956
rect 28588 5012 28644 5022
rect 28588 5010 28756 5012
rect 28588 4958 28590 5010
rect 28642 4958 28756 5010
rect 28588 4956 28756 4958
rect 28588 4946 28644 4956
rect 28588 4340 28644 4350
rect 28588 4246 28644 4284
rect 28140 4228 28196 4238
rect 27916 4226 28196 4228
rect 27916 4174 28142 4226
rect 28194 4174 28196 4226
rect 27916 4172 28196 4174
rect 28140 4162 28196 4172
rect 26908 3726 26910 3778
rect 26962 3726 26964 3778
rect 26908 3714 26964 3726
rect 27580 3780 27636 3790
rect 26572 3602 26628 3612
rect 26460 3554 26516 3566
rect 26460 3502 26462 3554
rect 26514 3502 26516 3554
rect 26236 3390 26238 3442
rect 26290 3390 26292 3442
rect 26236 3378 26292 3390
rect 26348 3444 26404 3454
rect 26460 3444 26516 3502
rect 27020 3556 27076 3566
rect 27020 3462 27076 3500
rect 26404 3388 26516 3444
rect 27468 3444 27524 3482
rect 25404 3164 25668 3174
rect 25460 3108 25508 3164
rect 25564 3108 25612 3164
rect 25404 3098 25668 3108
rect 25116 1138 25172 1148
rect 26348 980 26404 3388
rect 27468 3378 27524 3388
rect 24444 924 24836 980
rect 26012 924 26404 980
rect 24444 800 24500 924
rect 26012 800 26068 924
rect 27580 800 27636 3724
rect 27916 3780 27972 3790
rect 28588 3780 28644 3790
rect 27916 3778 28420 3780
rect 27916 3726 27918 3778
rect 27970 3726 28420 3778
rect 27916 3724 28420 3726
rect 27916 3714 27972 3724
rect 28364 3442 28420 3724
rect 28588 3554 28644 3724
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 28364 3390 28366 3442
rect 28418 3390 28420 3442
rect 28364 3378 28420 3390
rect 28700 3444 28756 4956
rect 29260 4898 29316 4910
rect 29260 4846 29262 4898
rect 29314 4846 29316 4898
rect 29260 4450 29316 4846
rect 29260 4398 29262 4450
rect 29314 4398 29316 4450
rect 29260 4386 29316 4398
rect 30268 4228 30324 4238
rect 29436 3948 29700 3958
rect 29492 3892 29540 3948
rect 29596 3892 29644 3948
rect 29436 3882 29700 3892
rect 28700 3378 28756 3388
rect 29148 3556 29204 3566
rect 29148 800 29204 3500
rect 29596 3556 29652 3566
rect 29596 3462 29652 3500
rect 30268 3556 30324 4172
rect 30268 3462 30324 3500
rect 29372 3444 29428 3454
rect 29372 3350 29428 3388
rect 30604 3442 30660 5740
rect 30828 4900 30884 5854
rect 31164 5908 31220 6412
rect 31948 6356 32004 6524
rect 31724 6132 31780 6142
rect 31724 6038 31780 6076
rect 31948 6130 32004 6300
rect 31948 6078 31950 6130
rect 32002 6078 32004 6130
rect 31948 6066 32004 6078
rect 31276 5908 31332 5918
rect 31164 5906 31332 5908
rect 31164 5854 31278 5906
rect 31330 5854 31332 5906
rect 31164 5852 31332 5854
rect 31276 5842 31332 5852
rect 30940 5794 30996 5806
rect 30940 5742 30942 5794
rect 30994 5742 30996 5794
rect 30940 5012 30996 5742
rect 31836 5794 31892 5806
rect 31836 5742 31838 5794
rect 31890 5742 31892 5794
rect 31836 5236 31892 5742
rect 31724 5180 31892 5236
rect 30940 4956 31668 5012
rect 30828 4844 31444 4900
rect 31276 4228 31332 4238
rect 30604 3390 30606 3442
rect 30658 3390 30660 3442
rect 30604 3378 30660 3390
rect 30716 3668 30772 3678
rect 30716 3444 30772 3612
rect 30940 3444 30996 3454
rect 30716 3442 30996 3444
rect 30716 3390 30942 3442
rect 30994 3390 30996 3442
rect 30716 3388 30996 3390
rect 30716 800 30772 3388
rect 30940 3378 30996 3388
rect 31276 3442 31332 4172
rect 31388 4226 31444 4844
rect 31612 4338 31668 4956
rect 31724 4452 31780 5180
rect 31948 5124 32004 5134
rect 31836 5068 31948 5124
rect 31836 4562 31892 5068
rect 31948 5058 32004 5068
rect 31836 4510 31838 4562
rect 31890 4510 31892 4562
rect 31836 4498 31892 4510
rect 31724 4386 31780 4396
rect 32060 4450 32116 7420
rect 32172 7382 32228 7420
rect 32172 6580 32228 6590
rect 32284 6580 32340 7644
rect 32508 6690 32564 8092
rect 32508 6638 32510 6690
rect 32562 6638 32564 6690
rect 32508 6626 32564 6638
rect 32172 6578 32340 6580
rect 32172 6526 32174 6578
rect 32226 6526 32340 6578
rect 32172 6524 32340 6526
rect 32172 6514 32228 6524
rect 32396 5796 32452 5806
rect 32396 5794 32564 5796
rect 32396 5742 32398 5794
rect 32450 5742 32564 5794
rect 32396 5740 32564 5742
rect 32396 5730 32452 5740
rect 32284 5684 32340 5694
rect 32284 5590 32340 5628
rect 32396 5124 32452 5134
rect 32396 5030 32452 5068
rect 32060 4398 32062 4450
rect 32114 4398 32116 4450
rect 32060 4386 32116 4398
rect 32172 4452 32228 4462
rect 31612 4286 31614 4338
rect 31666 4286 31668 4338
rect 31612 4274 31668 4286
rect 32172 4338 32228 4396
rect 32172 4286 32174 4338
rect 32226 4286 32228 4338
rect 32172 4274 32228 4286
rect 31388 4174 31390 4226
rect 31442 4174 31444 4226
rect 31388 4162 31444 4174
rect 31276 3390 31278 3442
rect 31330 3390 31332 3442
rect 31276 3378 31332 3390
rect 32284 3780 32340 3790
rect 32284 3554 32340 3724
rect 32284 3502 32286 3554
rect 32338 3502 32340 3554
rect 32284 800 32340 3502
rect 32508 3442 32564 5740
rect 32508 3390 32510 3442
rect 32562 3390 32564 3442
rect 32508 3378 32564 3390
rect 32732 3444 32788 9436
rect 32844 6578 32900 11788
rect 33180 11508 33236 11518
rect 33180 11414 33236 11452
rect 32956 10836 33012 10846
rect 33180 10836 33236 10846
rect 33012 10834 33236 10836
rect 33012 10782 33182 10834
rect 33234 10782 33236 10834
rect 33012 10780 33236 10782
rect 32956 10770 33012 10780
rect 33180 10770 33236 10780
rect 33068 10500 33124 10510
rect 33068 9826 33124 10444
rect 33292 10276 33348 13580
rect 33468 12572 33732 12582
rect 33524 12516 33572 12572
rect 33628 12516 33676 12572
rect 33468 12506 33732 12516
rect 33852 11956 33908 11966
rect 33468 11004 33732 11014
rect 33524 10948 33572 11004
rect 33628 10948 33676 11004
rect 33468 10938 33732 10948
rect 33068 9774 33070 9826
rect 33122 9774 33124 9826
rect 33068 8260 33124 9774
rect 32844 6526 32846 6578
rect 32898 6526 32900 6578
rect 32844 6514 32900 6526
rect 32956 8258 33124 8260
rect 32956 8206 33070 8258
rect 33122 8206 33124 8258
rect 32956 8204 33124 8206
rect 32844 5348 32900 5358
rect 32844 4564 32900 5292
rect 32956 5124 33012 8204
rect 33068 8194 33124 8204
rect 33180 10220 33348 10276
rect 33180 7698 33236 10220
rect 33468 9436 33732 9446
rect 33524 9380 33572 9436
rect 33628 9380 33676 9436
rect 33468 9370 33732 9380
rect 33292 9268 33348 9278
rect 33292 9174 33348 9212
rect 33852 8372 33908 11900
rect 33468 7868 33732 7878
rect 33524 7812 33572 7868
rect 33628 7812 33676 7868
rect 33468 7802 33732 7812
rect 33180 7646 33182 7698
rect 33234 7646 33236 7698
rect 33180 7634 33236 7646
rect 33180 7476 33236 7486
rect 33180 6690 33236 7420
rect 33852 7476 33908 8316
rect 33852 7410 33908 7420
rect 33180 6638 33182 6690
rect 33234 6638 33236 6690
rect 33180 6626 33236 6638
rect 33468 6300 33732 6310
rect 33068 6244 33124 6254
rect 33524 6244 33572 6300
rect 33628 6244 33676 6300
rect 33468 6234 33732 6244
rect 33068 6130 33124 6188
rect 33068 6078 33070 6130
rect 33122 6078 33124 6130
rect 33068 6066 33124 6078
rect 33180 5796 33236 5806
rect 33180 5702 33236 5740
rect 33068 5124 33124 5134
rect 32956 5122 33124 5124
rect 32956 5070 33070 5122
rect 33122 5070 33124 5122
rect 32956 5068 33124 5070
rect 33068 5058 33124 5068
rect 33468 4732 33732 4742
rect 33524 4676 33572 4732
rect 33628 4676 33676 4732
rect 33468 4666 33732 4676
rect 33068 4564 33124 4574
rect 32844 4562 33124 4564
rect 32844 4510 33070 4562
rect 33122 4510 33124 4562
rect 32844 4508 33124 4510
rect 33068 4498 33124 4508
rect 33180 4228 33236 4238
rect 33180 4134 33236 4172
rect 33180 4004 33236 4014
rect 33180 3554 33236 3948
rect 33180 3502 33182 3554
rect 33234 3502 33236 3554
rect 33180 3490 33236 3502
rect 33852 3556 33908 3566
rect 32844 3444 32900 3454
rect 32732 3442 32900 3444
rect 32732 3390 32846 3442
rect 32898 3390 32900 3442
rect 32732 3388 32900 3390
rect 32844 3378 32900 3388
rect 33468 3164 33732 3174
rect 33524 3108 33572 3164
rect 33628 3108 33676 3164
rect 33468 3098 33732 3108
rect 33852 800 33908 3500
rect 13804 700 14308 756
rect 15008 0 15120 800
rect 16576 0 16688 800
rect 18144 0 18256 800
rect 19712 0 19824 800
rect 21280 0 21392 800
rect 22848 0 22960 800
rect 24416 0 24528 800
rect 25984 0 26096 800
rect 27552 0 27664 800
rect 29120 0 29232 800
rect 30688 0 30800 800
rect 32256 0 32368 800
rect 33824 0 33936 800
<< via2 >>
rect 4956 31836 5012 31892
rect 6076 31836 6132 31892
rect 6860 31724 6916 31780
rect 5068 31500 5124 31556
rect 3724 31106 3780 31108
rect 3724 31054 3726 31106
rect 3726 31054 3778 31106
rect 3778 31054 3780 31106
rect 3724 31052 3780 31054
rect 5852 31218 5908 31220
rect 5852 31166 5854 31218
rect 5854 31166 5906 31218
rect 5906 31166 5908 31218
rect 5852 31164 5908 31166
rect 5244 30602 5300 30604
rect 5244 30550 5246 30602
rect 5246 30550 5298 30602
rect 5298 30550 5300 30602
rect 5244 30548 5300 30550
rect 5348 30602 5404 30604
rect 5348 30550 5350 30602
rect 5350 30550 5402 30602
rect 5402 30550 5404 30602
rect 5348 30548 5404 30550
rect 5452 30602 5508 30604
rect 5452 30550 5454 30602
rect 5454 30550 5506 30602
rect 5506 30550 5508 30602
rect 5452 30548 5508 30550
rect 1708 29260 1764 29316
rect 2940 30098 2996 30100
rect 2940 30046 2942 30098
rect 2942 30046 2994 30098
rect 2994 30046 2996 30098
rect 2940 30044 2996 30046
rect 3948 30044 4004 30100
rect 2268 29260 2324 29316
rect 5516 29650 5572 29652
rect 5516 29598 5518 29650
rect 5518 29598 5570 29650
rect 5570 29598 5572 29650
rect 5516 29596 5572 29598
rect 4508 29314 4564 29316
rect 4508 29262 4510 29314
rect 4510 29262 4562 29314
rect 4562 29262 4564 29314
rect 4508 29260 4564 29262
rect 5292 29260 5348 29316
rect 4060 28700 4116 28756
rect 4620 29036 4676 29092
rect 4844 28812 4900 28868
rect 4620 27580 4676 27636
rect 2940 27186 2996 27188
rect 2940 27134 2942 27186
rect 2942 27134 2994 27186
rect 2994 27134 2996 27186
rect 2940 27132 2996 27134
rect 5244 29034 5300 29036
rect 5244 28982 5246 29034
rect 5246 28982 5298 29034
rect 5298 28982 5300 29034
rect 5244 28980 5300 28982
rect 5348 29034 5404 29036
rect 5348 28982 5350 29034
rect 5350 28982 5402 29034
rect 5402 28982 5404 29034
rect 5348 28980 5404 28982
rect 5452 29034 5508 29036
rect 5452 28982 5454 29034
rect 5454 28982 5506 29034
rect 5506 28982 5508 29034
rect 5452 28980 5508 28982
rect 5180 28642 5236 28644
rect 5180 28590 5182 28642
rect 5182 28590 5234 28642
rect 5234 28590 5236 28642
rect 5180 28588 5236 28590
rect 6412 30098 6468 30100
rect 6412 30046 6414 30098
rect 6414 30046 6466 30098
rect 6466 30046 6468 30098
rect 6412 30044 6468 30046
rect 7196 31164 7252 31220
rect 7980 31836 8036 31892
rect 6860 29596 6916 29652
rect 7196 30268 7252 30324
rect 7644 30044 7700 30100
rect 5852 29148 5908 29204
rect 6076 28754 6132 28756
rect 6076 28702 6078 28754
rect 6078 28702 6130 28754
rect 6130 28702 6132 28754
rect 6076 28700 6132 28702
rect 5244 27466 5300 27468
rect 5244 27414 5246 27466
rect 5246 27414 5298 27466
rect 5298 27414 5300 27466
rect 5244 27412 5300 27414
rect 5348 27466 5404 27468
rect 5348 27414 5350 27466
rect 5350 27414 5402 27466
rect 5402 27414 5404 27466
rect 5348 27412 5404 27414
rect 5452 27466 5508 27468
rect 5452 27414 5454 27466
rect 5454 27414 5506 27466
rect 5506 27414 5508 27466
rect 5452 27412 5508 27414
rect 3388 26012 3444 26068
rect 4732 25676 4788 25732
rect 2492 25228 2548 25284
rect 4060 25282 4116 25284
rect 4060 25230 4062 25282
rect 4062 25230 4114 25282
rect 4114 25230 4116 25282
rect 4060 25228 4116 25230
rect 4508 24780 4564 24836
rect 4620 24610 4676 24612
rect 4620 24558 4622 24610
rect 4622 24558 4674 24610
rect 4674 24558 4676 24610
rect 4620 24556 4676 24558
rect 3948 23996 4004 24052
rect 4956 26572 5012 26628
rect 5068 26348 5124 26404
rect 4844 23884 4900 23940
rect 4956 26236 5012 26292
rect 5516 26178 5572 26180
rect 5516 26126 5518 26178
rect 5518 26126 5570 26178
rect 5570 26126 5572 26178
rect 5516 26124 5572 26126
rect 5244 25898 5300 25900
rect 5244 25846 5246 25898
rect 5246 25846 5298 25898
rect 5298 25846 5300 25898
rect 5244 25844 5300 25846
rect 5348 25898 5404 25900
rect 5348 25846 5350 25898
rect 5350 25846 5402 25898
rect 5402 25846 5404 25898
rect 5348 25844 5404 25846
rect 5452 25898 5508 25900
rect 5452 25846 5454 25898
rect 5454 25846 5506 25898
rect 5506 25846 5508 25898
rect 5452 25844 5508 25846
rect 2492 23324 2548 23380
rect 5068 25676 5124 25732
rect 1820 22092 1876 22148
rect 4620 21868 4676 21924
rect 2492 21756 2548 21812
rect 2492 21474 2548 21476
rect 2492 21422 2494 21474
rect 2494 21422 2546 21474
rect 2546 21422 2548 21474
rect 2492 21420 2548 21422
rect 4172 21420 4228 21476
rect 4620 20802 4676 20804
rect 4620 20750 4622 20802
rect 4622 20750 4674 20802
rect 4674 20750 4676 20802
rect 4620 20748 4676 20750
rect 4620 20524 4676 20580
rect 4620 20018 4676 20020
rect 4620 19966 4622 20018
rect 4622 19966 4674 20018
rect 4674 19966 4676 20018
rect 4620 19964 4676 19966
rect 4060 19404 4116 19460
rect 3612 19068 3668 19124
rect 4508 18956 4564 19012
rect 4620 19068 4676 19124
rect 3612 18732 3668 18788
rect 3052 18674 3108 18676
rect 3052 18622 3054 18674
rect 3054 18622 3106 18674
rect 3106 18622 3108 18674
rect 3052 18620 3108 18622
rect 3724 18620 3780 18676
rect 2492 18284 2548 18340
rect 3276 18450 3332 18452
rect 3276 18398 3278 18450
rect 3278 18398 3330 18450
rect 3330 18398 3332 18450
rect 3276 18396 3332 18398
rect 3948 18450 4004 18452
rect 3948 18398 3950 18450
rect 3950 18398 4002 18450
rect 4002 18398 4004 18450
rect 3948 18396 4004 18398
rect 4396 18450 4452 18452
rect 4396 18398 4398 18450
rect 4398 18398 4450 18450
rect 4450 18398 4452 18450
rect 4396 18396 4452 18398
rect 4172 18338 4228 18340
rect 4172 18286 4174 18338
rect 4174 18286 4226 18338
rect 4226 18286 4228 18338
rect 4172 18284 4228 18286
rect 3500 18172 3556 18228
rect 2492 17554 2548 17556
rect 2492 17502 2494 17554
rect 2494 17502 2546 17554
rect 2546 17502 2548 17554
rect 2492 17500 2548 17502
rect 3948 17724 4004 17780
rect 4508 17724 4564 17780
rect 4508 17500 4564 17556
rect 4956 23324 5012 23380
rect 6636 29484 6692 29540
rect 6524 29260 6580 29316
rect 6524 28924 6580 28980
rect 6300 28588 6356 28644
rect 6300 28028 6356 28084
rect 6300 27858 6356 27860
rect 6300 27806 6302 27858
rect 6302 27806 6354 27858
rect 6354 27806 6356 27858
rect 6300 27804 6356 27806
rect 6188 27468 6244 27524
rect 5964 26962 6020 26964
rect 5964 26910 5966 26962
rect 5966 26910 6018 26962
rect 6018 26910 6020 26962
rect 5964 26908 6020 26910
rect 6748 29314 6804 29316
rect 6748 29262 6750 29314
rect 6750 29262 6802 29314
rect 6802 29262 6804 29314
rect 6748 29260 6804 29262
rect 6636 28812 6692 28868
rect 6636 27804 6692 27860
rect 6748 27746 6804 27748
rect 6748 27694 6750 27746
rect 6750 27694 6802 27746
rect 6802 27694 6804 27746
rect 6748 27692 6804 27694
rect 6748 27468 6804 27524
rect 6636 26684 6692 26740
rect 6300 26124 6356 26180
rect 6076 25788 6132 25844
rect 6188 26012 6244 26068
rect 5180 24892 5236 24948
rect 5292 24834 5348 24836
rect 5292 24782 5294 24834
rect 5294 24782 5346 24834
rect 5346 24782 5348 24834
rect 5292 24780 5348 24782
rect 5516 24722 5572 24724
rect 5516 24670 5518 24722
rect 5518 24670 5570 24722
rect 5570 24670 5572 24722
rect 5516 24668 5572 24670
rect 5244 24330 5300 24332
rect 5244 24278 5246 24330
rect 5246 24278 5298 24330
rect 5298 24278 5300 24330
rect 5244 24276 5300 24278
rect 5348 24330 5404 24332
rect 5348 24278 5350 24330
rect 5350 24278 5402 24330
rect 5402 24278 5404 24330
rect 5348 24276 5404 24278
rect 5452 24330 5508 24332
rect 5452 24278 5454 24330
rect 5454 24278 5506 24330
rect 5506 24278 5508 24330
rect 5452 24276 5508 24278
rect 5404 23436 5460 23492
rect 5068 23212 5124 23268
rect 6524 25788 6580 25844
rect 6076 25228 6132 25284
rect 5964 24892 6020 24948
rect 5964 24050 6020 24052
rect 5964 23998 5966 24050
rect 5966 23998 6018 24050
rect 6018 23998 6020 24050
rect 5964 23996 6020 23998
rect 6300 25228 6356 25284
rect 6748 26460 6804 26516
rect 6748 26290 6804 26292
rect 6748 26238 6750 26290
rect 6750 26238 6802 26290
rect 6802 26238 6804 26290
rect 6748 26236 6804 26238
rect 6748 26012 6804 26068
rect 7084 27020 7140 27076
rect 6972 26962 7028 26964
rect 6972 26910 6974 26962
rect 6974 26910 7026 26962
rect 7026 26910 7028 26962
rect 6972 26908 7028 26910
rect 7196 26962 7252 26964
rect 7196 26910 7198 26962
rect 7198 26910 7250 26962
rect 7250 26910 7252 26962
rect 7196 26908 7252 26910
rect 7308 26850 7364 26852
rect 7308 26798 7310 26850
rect 7310 26798 7362 26850
rect 7362 26798 7364 26850
rect 7308 26796 7364 26798
rect 8764 32060 8820 32116
rect 8316 29932 8372 29988
rect 7756 29426 7812 29428
rect 7756 29374 7758 29426
rect 7758 29374 7810 29426
rect 7810 29374 7812 29426
rect 7756 29372 7812 29374
rect 8092 28924 8148 28980
rect 7308 26572 7364 26628
rect 7196 26348 7252 26404
rect 6412 25116 6468 25172
rect 6300 24892 6356 24948
rect 6636 25004 6692 25060
rect 7084 25452 7140 25508
rect 7420 26402 7476 26404
rect 7420 26350 7422 26402
rect 7422 26350 7474 26402
rect 7474 26350 7476 26402
rect 7420 26348 7476 26350
rect 6636 24668 6692 24724
rect 6524 24556 6580 24612
rect 6412 24444 6468 24500
rect 6300 23996 6356 24052
rect 5852 23436 5908 23492
rect 5740 23324 5796 23380
rect 5292 23100 5348 23156
rect 5244 22762 5300 22764
rect 5244 22710 5246 22762
rect 5246 22710 5298 22762
rect 5298 22710 5300 22762
rect 5244 22708 5300 22710
rect 5348 22762 5404 22764
rect 5348 22710 5350 22762
rect 5350 22710 5402 22762
rect 5402 22710 5404 22762
rect 5348 22708 5404 22710
rect 5452 22762 5508 22764
rect 5452 22710 5454 22762
rect 5454 22710 5506 22762
rect 5506 22710 5508 22762
rect 5452 22708 5508 22710
rect 5852 23266 5908 23268
rect 5852 23214 5854 23266
rect 5854 23214 5906 23266
rect 5906 23214 5908 23266
rect 5852 23212 5908 23214
rect 5068 22092 5124 22148
rect 4956 20748 5012 20804
rect 5292 21810 5348 21812
rect 5292 21758 5294 21810
rect 5294 21758 5346 21810
rect 5346 21758 5348 21810
rect 5292 21756 5348 21758
rect 5852 21644 5908 21700
rect 5292 21586 5348 21588
rect 5292 21534 5294 21586
rect 5294 21534 5346 21586
rect 5346 21534 5348 21586
rect 5292 21532 5348 21534
rect 5244 21194 5300 21196
rect 5244 21142 5246 21194
rect 5246 21142 5298 21194
rect 5298 21142 5300 21194
rect 5244 21140 5300 21142
rect 5348 21194 5404 21196
rect 5348 21142 5350 21194
rect 5350 21142 5402 21194
rect 5402 21142 5404 21194
rect 5348 21140 5404 21142
rect 5452 21194 5508 21196
rect 5452 21142 5454 21194
rect 5454 21142 5506 21194
rect 5506 21142 5508 21194
rect 5452 21140 5508 21142
rect 5068 20300 5124 20356
rect 5740 20578 5796 20580
rect 5740 20526 5742 20578
rect 5742 20526 5794 20578
rect 5794 20526 5796 20578
rect 5740 20524 5796 20526
rect 5404 20076 5460 20132
rect 5740 20300 5796 20356
rect 5180 19740 5236 19796
rect 5244 19626 5300 19628
rect 5244 19574 5246 19626
rect 5246 19574 5298 19626
rect 5298 19574 5300 19626
rect 5244 19572 5300 19574
rect 5348 19626 5404 19628
rect 5348 19574 5350 19626
rect 5350 19574 5402 19626
rect 5402 19574 5404 19626
rect 5348 19572 5404 19574
rect 5452 19626 5508 19628
rect 5452 19574 5454 19626
rect 5454 19574 5506 19626
rect 5506 19574 5508 19626
rect 5452 19572 5508 19574
rect 5740 19458 5796 19460
rect 5740 19406 5742 19458
rect 5742 19406 5794 19458
rect 5794 19406 5796 19458
rect 5740 19404 5796 19406
rect 5292 18956 5348 19012
rect 4844 18450 4900 18452
rect 4844 18398 4846 18450
rect 4846 18398 4898 18450
rect 4898 18398 4900 18450
rect 4844 18396 4900 18398
rect 5180 18620 5236 18676
rect 5068 18562 5124 18564
rect 5068 18510 5070 18562
rect 5070 18510 5122 18562
rect 5122 18510 5124 18562
rect 5068 18508 5124 18510
rect 5292 18508 5348 18564
rect 4732 17052 4788 17108
rect 6972 24722 7028 24724
rect 6972 24670 6974 24722
rect 6974 24670 7026 24722
rect 7026 24670 7028 24722
rect 6972 24668 7028 24670
rect 7308 24780 7364 24836
rect 6636 23996 6692 24052
rect 7308 24332 7364 24388
rect 7868 28364 7924 28420
rect 8092 28082 8148 28084
rect 8092 28030 8094 28082
rect 8094 28030 8146 28082
rect 8146 28030 8148 28082
rect 8092 28028 8148 28030
rect 7756 27970 7812 27972
rect 7756 27918 7758 27970
rect 7758 27918 7810 27970
rect 7810 27918 7812 27970
rect 7756 27916 7812 27918
rect 8540 29372 8596 29428
rect 8652 29484 8708 29540
rect 7756 27468 7812 27524
rect 8540 28028 8596 28084
rect 9436 31836 9492 31892
rect 9276 31386 9332 31388
rect 9276 31334 9278 31386
rect 9278 31334 9330 31386
rect 9330 31334 9332 31386
rect 9276 31332 9332 31334
rect 9380 31386 9436 31388
rect 9380 31334 9382 31386
rect 9382 31334 9434 31386
rect 9434 31334 9436 31386
rect 9380 31332 9436 31334
rect 9484 31386 9540 31388
rect 9484 31334 9486 31386
rect 9486 31334 9538 31386
rect 9538 31334 9540 31386
rect 9484 31332 9540 31334
rect 8876 29986 8932 29988
rect 8876 29934 8878 29986
rect 8878 29934 8930 29986
rect 8930 29934 8932 29986
rect 8876 29932 8932 29934
rect 9436 29986 9492 29988
rect 9436 29934 9438 29986
rect 9438 29934 9490 29986
rect 9490 29934 9492 29986
rect 9436 29932 9492 29934
rect 9276 29818 9332 29820
rect 9276 29766 9278 29818
rect 9278 29766 9330 29818
rect 9330 29766 9332 29818
rect 9276 29764 9332 29766
rect 9380 29818 9436 29820
rect 9380 29766 9382 29818
rect 9382 29766 9434 29818
rect 9434 29766 9436 29818
rect 9380 29764 9436 29766
rect 9484 29818 9540 29820
rect 9484 29766 9486 29818
rect 9486 29766 9538 29818
rect 9538 29766 9540 29818
rect 9484 29764 9540 29766
rect 9100 29650 9156 29652
rect 9100 29598 9102 29650
rect 9102 29598 9154 29650
rect 9154 29598 9156 29650
rect 9100 29596 9156 29598
rect 9660 29484 9716 29540
rect 9100 29036 9156 29092
rect 9324 29260 9380 29316
rect 8764 27916 8820 27972
rect 9212 28812 9268 28868
rect 7980 27186 8036 27188
rect 7980 27134 7982 27186
rect 7982 27134 8034 27186
rect 8034 27134 8036 27186
rect 7980 27132 8036 27134
rect 8428 27356 8484 27412
rect 7868 26460 7924 26516
rect 7868 26012 7924 26068
rect 7980 26796 8036 26852
rect 8204 27020 8260 27076
rect 8092 26348 8148 26404
rect 7980 26124 8036 26180
rect 8540 27244 8596 27300
rect 8652 27580 8708 27636
rect 9660 29314 9716 29316
rect 9660 29262 9662 29314
rect 9662 29262 9714 29314
rect 9714 29262 9716 29314
rect 9660 29260 9716 29262
rect 9772 29036 9828 29092
rect 9772 28418 9828 28420
rect 9772 28366 9774 28418
rect 9774 28366 9826 28418
rect 9826 28366 9828 28418
rect 9772 28364 9828 28366
rect 9276 28250 9332 28252
rect 9276 28198 9278 28250
rect 9278 28198 9330 28250
rect 9330 28198 9332 28250
rect 9276 28196 9332 28198
rect 9380 28250 9436 28252
rect 9380 28198 9382 28250
rect 9382 28198 9434 28250
rect 9434 28198 9436 28250
rect 9380 28196 9436 28198
rect 9484 28250 9540 28252
rect 9484 28198 9486 28250
rect 9486 28198 9538 28250
rect 9538 28198 9540 28250
rect 9484 28196 9540 28198
rect 9660 28140 9716 28196
rect 9212 27916 9268 27972
rect 9100 27132 9156 27188
rect 9548 27916 9604 27972
rect 8876 27020 8932 27076
rect 9996 28530 10052 28532
rect 9996 28478 9998 28530
rect 9998 28478 10050 28530
rect 10050 28478 10052 28530
rect 9996 28476 10052 28478
rect 10556 29484 10612 29540
rect 10332 29372 10388 29428
rect 10892 29314 10948 29316
rect 10892 29262 10894 29314
rect 10894 29262 10946 29314
rect 10946 29262 10948 29314
rect 10892 29260 10948 29262
rect 11004 28700 11060 28756
rect 10220 28364 10276 28420
rect 10892 28476 10948 28532
rect 10780 28252 10836 28308
rect 9772 27580 9828 27636
rect 9660 27356 9716 27412
rect 10780 27970 10836 27972
rect 10780 27918 10782 27970
rect 10782 27918 10834 27970
rect 10834 27918 10836 27970
rect 10780 27916 10836 27918
rect 9772 26908 9828 26964
rect 8540 26684 8596 26740
rect 9276 26682 9332 26684
rect 9276 26630 9278 26682
rect 9278 26630 9330 26682
rect 9330 26630 9332 26682
rect 9276 26628 9332 26630
rect 9380 26682 9436 26684
rect 9380 26630 9382 26682
rect 9382 26630 9434 26682
rect 9434 26630 9436 26682
rect 9380 26628 9436 26630
rect 9484 26682 9540 26684
rect 9484 26630 9486 26682
rect 9486 26630 9538 26682
rect 9538 26630 9540 26682
rect 9484 26628 9540 26630
rect 9212 26236 9268 26292
rect 8428 25676 8484 25732
rect 8876 25676 8932 25732
rect 7756 25116 7812 25172
rect 7420 24220 7476 24276
rect 8540 25116 8596 25172
rect 7868 24220 7924 24276
rect 7196 23938 7252 23940
rect 7196 23886 7198 23938
rect 7198 23886 7250 23938
rect 7250 23886 7252 23938
rect 7196 23884 7252 23886
rect 7644 23714 7700 23716
rect 7644 23662 7646 23714
rect 7646 23662 7698 23714
rect 7698 23662 7700 23714
rect 7644 23660 7700 23662
rect 6636 23436 6692 23492
rect 6972 23378 7028 23380
rect 6972 23326 6974 23378
rect 6974 23326 7026 23378
rect 7026 23326 7028 23378
rect 6972 23324 7028 23326
rect 6636 22988 6692 23044
rect 6188 21810 6244 21812
rect 6188 21758 6190 21810
rect 6190 21758 6242 21810
rect 6242 21758 6244 21810
rect 6188 21756 6244 21758
rect 6076 21698 6132 21700
rect 6076 21646 6078 21698
rect 6078 21646 6130 21698
rect 6130 21646 6132 21698
rect 6076 21644 6132 21646
rect 5740 19010 5796 19012
rect 5740 18958 5742 19010
rect 5742 18958 5794 19010
rect 5794 18958 5796 19010
rect 5740 18956 5796 18958
rect 6076 19964 6132 20020
rect 5628 18172 5684 18228
rect 5244 18058 5300 18060
rect 5244 18006 5246 18058
rect 5246 18006 5298 18058
rect 5298 18006 5300 18058
rect 5244 18004 5300 18006
rect 5348 18058 5404 18060
rect 5348 18006 5350 18058
rect 5350 18006 5402 18058
rect 5402 18006 5404 18058
rect 5348 18004 5404 18006
rect 5452 18058 5508 18060
rect 5452 18006 5454 18058
rect 5454 18006 5506 18058
rect 5506 18006 5508 18058
rect 5452 18004 5508 18006
rect 4172 16604 4228 16660
rect 4844 16604 4900 16660
rect 4956 16098 5012 16100
rect 4956 16046 4958 16098
rect 4958 16046 5010 16098
rect 5010 16046 5012 16098
rect 4956 16044 5012 16046
rect 2492 15820 2548 15876
rect 4508 15874 4564 15876
rect 4508 15822 4510 15874
rect 4510 15822 4562 15874
rect 4562 15822 4564 15874
rect 4508 15820 4564 15822
rect 3948 15708 4004 15764
rect 2492 15148 2548 15204
rect 5180 17164 5236 17220
rect 5404 17164 5460 17220
rect 8540 24220 8596 24276
rect 8652 24892 8708 24948
rect 7308 23154 7364 23156
rect 7308 23102 7310 23154
rect 7310 23102 7362 23154
rect 7362 23102 7364 23154
rect 7308 23100 7364 23102
rect 7196 22988 7252 23044
rect 6748 21810 6804 21812
rect 6748 21758 6750 21810
rect 6750 21758 6802 21810
rect 6802 21758 6804 21810
rect 6748 21756 6804 21758
rect 6972 21586 7028 21588
rect 6972 21534 6974 21586
rect 6974 21534 7026 21586
rect 7026 21534 7028 21586
rect 6972 21532 7028 21534
rect 6636 20972 6692 21028
rect 7308 20972 7364 21028
rect 6860 20802 6916 20804
rect 6860 20750 6862 20802
rect 6862 20750 6914 20802
rect 6914 20750 6916 20802
rect 6860 20748 6916 20750
rect 7196 20300 7252 20356
rect 7308 20748 7364 20804
rect 6412 19964 6468 20020
rect 6300 19068 6356 19124
rect 5964 18674 6020 18676
rect 5964 18622 5966 18674
rect 5966 18622 6018 18674
rect 6018 18622 6020 18674
rect 5964 18620 6020 18622
rect 7644 19852 7700 19908
rect 7532 19740 7588 19796
rect 6300 18450 6356 18452
rect 6300 18398 6302 18450
rect 6302 18398 6354 18450
rect 6354 18398 6356 18450
rect 6300 18396 6356 18398
rect 6748 18450 6804 18452
rect 6748 18398 6750 18450
rect 6750 18398 6802 18450
rect 6802 18398 6804 18450
rect 6748 18396 6804 18398
rect 6748 17724 6804 17780
rect 5852 17666 5908 17668
rect 5852 17614 5854 17666
rect 5854 17614 5906 17666
rect 5906 17614 5908 17666
rect 5852 17612 5908 17614
rect 6636 17106 6692 17108
rect 6636 17054 6638 17106
rect 6638 17054 6690 17106
rect 6690 17054 6692 17106
rect 6636 17052 6692 17054
rect 5244 16490 5300 16492
rect 5244 16438 5246 16490
rect 5246 16438 5298 16490
rect 5298 16438 5300 16490
rect 5244 16436 5300 16438
rect 5348 16490 5404 16492
rect 5348 16438 5350 16490
rect 5350 16438 5402 16490
rect 5402 16438 5404 16490
rect 5348 16436 5404 16438
rect 5452 16490 5508 16492
rect 5452 16438 5454 16490
rect 5454 16438 5506 16490
rect 5506 16438 5508 16490
rect 5452 16436 5508 16438
rect 5628 16098 5684 16100
rect 5628 16046 5630 16098
rect 5630 16046 5682 16098
rect 5682 16046 5684 16098
rect 5628 16044 5684 16046
rect 4620 15484 4676 15540
rect 5292 15538 5348 15540
rect 5292 15486 5294 15538
rect 5294 15486 5346 15538
rect 5346 15486 5348 15538
rect 5292 15484 5348 15486
rect 5404 15314 5460 15316
rect 5404 15262 5406 15314
rect 5406 15262 5458 15314
rect 5458 15262 5460 15314
rect 5404 15260 5460 15262
rect 6300 16994 6356 16996
rect 6300 16942 6302 16994
rect 6302 16942 6354 16994
rect 6354 16942 6356 16994
rect 6300 16940 6356 16942
rect 5852 15708 5908 15764
rect 5740 15484 5796 15540
rect 5244 14922 5300 14924
rect 5244 14870 5246 14922
rect 5246 14870 5298 14922
rect 5298 14870 5300 14922
rect 5244 14868 5300 14870
rect 5348 14922 5404 14924
rect 5348 14870 5350 14922
rect 5350 14870 5402 14922
rect 5402 14870 5404 14922
rect 5348 14868 5404 14870
rect 5452 14922 5508 14924
rect 5452 14870 5454 14922
rect 5454 14870 5506 14922
rect 5506 14870 5508 14922
rect 5452 14868 5508 14870
rect 7196 17836 7252 17892
rect 7980 20076 8036 20132
rect 7980 19852 8036 19908
rect 8764 24780 8820 24836
rect 9996 26850 10052 26852
rect 9996 26798 9998 26850
rect 9998 26798 10050 26850
rect 10050 26798 10052 26850
rect 9996 26796 10052 26798
rect 9772 26402 9828 26404
rect 9772 26350 9774 26402
rect 9774 26350 9826 26402
rect 9826 26350 9828 26402
rect 9772 26348 9828 26350
rect 9996 26290 10052 26292
rect 9996 26238 9998 26290
rect 9998 26238 10050 26290
rect 10050 26238 10052 26290
rect 9996 26236 10052 26238
rect 9884 26012 9940 26068
rect 9996 25676 10052 25732
rect 9212 25618 9268 25620
rect 9212 25566 9214 25618
rect 9214 25566 9266 25618
rect 9266 25566 9268 25618
rect 9212 25564 9268 25566
rect 10332 26684 10388 26740
rect 9660 25394 9716 25396
rect 9660 25342 9662 25394
rect 9662 25342 9714 25394
rect 9714 25342 9716 25394
rect 9660 25340 9716 25342
rect 9548 25282 9604 25284
rect 9548 25230 9550 25282
rect 9550 25230 9602 25282
rect 9602 25230 9604 25282
rect 9548 25228 9604 25230
rect 9276 25114 9332 25116
rect 9276 25062 9278 25114
rect 9278 25062 9330 25114
rect 9330 25062 9332 25114
rect 9276 25060 9332 25062
rect 9380 25114 9436 25116
rect 9380 25062 9382 25114
rect 9382 25062 9434 25114
rect 9434 25062 9436 25114
rect 9380 25060 9436 25062
rect 9484 25114 9540 25116
rect 9484 25062 9486 25114
rect 9486 25062 9538 25114
rect 9538 25062 9540 25114
rect 9484 25060 9540 25062
rect 9996 25282 10052 25284
rect 9996 25230 9998 25282
rect 9998 25230 10050 25282
rect 10050 25230 10052 25282
rect 9996 25228 10052 25230
rect 9996 24780 10052 24836
rect 8428 23714 8484 23716
rect 8428 23662 8430 23714
rect 8430 23662 8482 23714
rect 8482 23662 8484 23714
rect 8428 23660 8484 23662
rect 8876 24220 8932 24276
rect 10108 24498 10164 24500
rect 10108 24446 10110 24498
rect 10110 24446 10162 24498
rect 10162 24446 10164 24498
rect 10108 24444 10164 24446
rect 9276 23546 9332 23548
rect 9276 23494 9278 23546
rect 9278 23494 9330 23546
rect 9330 23494 9332 23546
rect 9276 23492 9332 23494
rect 9380 23546 9436 23548
rect 9380 23494 9382 23546
rect 9382 23494 9434 23546
rect 9434 23494 9436 23546
rect 9380 23492 9436 23494
rect 9484 23546 9540 23548
rect 9484 23494 9486 23546
rect 9486 23494 9538 23546
rect 9538 23494 9540 23546
rect 9484 23492 9540 23494
rect 8428 20748 8484 20804
rect 8652 19906 8708 19908
rect 8652 19854 8654 19906
rect 8654 19854 8706 19906
rect 8706 19854 8708 19906
rect 8652 19852 8708 19854
rect 8204 18732 8260 18788
rect 7084 17388 7140 17444
rect 7084 16882 7140 16884
rect 7084 16830 7086 16882
rect 7086 16830 7138 16882
rect 7138 16830 7140 16882
rect 7084 16828 7140 16830
rect 6188 15484 6244 15540
rect 6636 15874 6692 15876
rect 6636 15822 6638 15874
rect 6638 15822 6690 15874
rect 6690 15822 6692 15874
rect 6636 15820 6692 15822
rect 6748 15538 6804 15540
rect 6748 15486 6750 15538
rect 6750 15486 6802 15538
rect 6802 15486 6804 15538
rect 6748 15484 6804 15486
rect 6412 15426 6468 15428
rect 6412 15374 6414 15426
rect 6414 15374 6466 15426
rect 6466 15374 6468 15426
rect 6412 15372 6468 15374
rect 6300 15314 6356 15316
rect 6300 15262 6302 15314
rect 6302 15262 6354 15314
rect 6354 15262 6356 15314
rect 6300 15260 6356 15262
rect 5964 15148 6020 15204
rect 6524 15260 6580 15316
rect 6972 15426 7028 15428
rect 6972 15374 6974 15426
rect 6974 15374 7026 15426
rect 7026 15374 7028 15426
rect 6972 15372 7028 15374
rect 7196 15372 7252 15428
rect 6748 15148 6804 15204
rect 7196 14530 7252 14532
rect 7196 14478 7198 14530
rect 7198 14478 7250 14530
rect 7250 14478 7252 14530
rect 7196 14476 7252 14478
rect 5244 13354 5300 13356
rect 5244 13302 5246 13354
rect 5246 13302 5298 13354
rect 5298 13302 5300 13354
rect 5244 13300 5300 13302
rect 5348 13354 5404 13356
rect 5348 13302 5350 13354
rect 5350 13302 5402 13354
rect 5402 13302 5404 13354
rect 5348 13300 5404 13302
rect 5452 13354 5508 13356
rect 5452 13302 5454 13354
rect 5454 13302 5506 13354
rect 5506 13302 5508 13354
rect 5452 13300 5508 13302
rect 6188 12908 6244 12964
rect 5244 11786 5300 11788
rect 5244 11734 5246 11786
rect 5246 11734 5298 11786
rect 5298 11734 5300 11786
rect 5244 11732 5300 11734
rect 5348 11786 5404 11788
rect 5348 11734 5350 11786
rect 5350 11734 5402 11786
rect 5402 11734 5404 11786
rect 5348 11732 5404 11734
rect 5452 11786 5508 11788
rect 5452 11734 5454 11786
rect 5454 11734 5506 11786
rect 5506 11734 5508 11786
rect 5452 11732 5508 11734
rect 7532 17164 7588 17220
rect 7756 17388 7812 17444
rect 8204 17442 8260 17444
rect 8204 17390 8206 17442
rect 8206 17390 8258 17442
rect 8258 17390 8260 17442
rect 8204 17388 8260 17390
rect 7644 16940 7700 16996
rect 7532 16828 7588 16884
rect 10108 23772 10164 23828
rect 9276 21978 9332 21980
rect 9276 21926 9278 21978
rect 9278 21926 9330 21978
rect 9330 21926 9332 21978
rect 9276 21924 9332 21926
rect 9380 21978 9436 21980
rect 9380 21926 9382 21978
rect 9382 21926 9434 21978
rect 9434 21926 9436 21978
rect 9380 21924 9436 21926
rect 9484 21978 9540 21980
rect 9484 21926 9486 21978
rect 9486 21926 9538 21978
rect 9538 21926 9540 21978
rect 9484 21924 9540 21926
rect 9548 21698 9604 21700
rect 9548 21646 9550 21698
rect 9550 21646 9602 21698
rect 9602 21646 9604 21698
rect 9548 21644 9604 21646
rect 8988 20860 9044 20916
rect 9660 20860 9716 20916
rect 9884 20412 9940 20468
rect 9276 20410 9332 20412
rect 9276 20358 9278 20410
rect 9278 20358 9330 20410
rect 9330 20358 9332 20410
rect 9276 20356 9332 20358
rect 9380 20410 9436 20412
rect 9380 20358 9382 20410
rect 9382 20358 9434 20410
rect 9434 20358 9436 20410
rect 9380 20356 9436 20358
rect 9484 20410 9540 20412
rect 9484 20358 9486 20410
rect 9486 20358 9538 20410
rect 9538 20358 9540 20410
rect 9484 20356 9540 20358
rect 9548 20188 9604 20244
rect 9772 20018 9828 20020
rect 9772 19966 9774 20018
rect 9774 19966 9826 20018
rect 9826 19966 9828 20018
rect 9772 19964 9828 19966
rect 9660 19180 9716 19236
rect 9100 19122 9156 19124
rect 9100 19070 9102 19122
rect 9102 19070 9154 19122
rect 9154 19070 9156 19122
rect 9100 19068 9156 19070
rect 8876 18956 8932 19012
rect 9100 18732 9156 18788
rect 9276 18842 9332 18844
rect 9276 18790 9278 18842
rect 9278 18790 9330 18842
rect 9330 18790 9332 18842
rect 9276 18788 9332 18790
rect 9380 18842 9436 18844
rect 9380 18790 9382 18842
rect 9382 18790 9434 18842
rect 9434 18790 9436 18842
rect 9380 18788 9436 18790
rect 9484 18842 9540 18844
rect 9484 18790 9486 18842
rect 9486 18790 9538 18842
rect 9538 18790 9540 18842
rect 9484 18788 9540 18790
rect 9212 18620 9268 18676
rect 8540 18508 8596 18564
rect 8988 18508 9044 18564
rect 9772 18732 9828 18788
rect 10668 26962 10724 26964
rect 10668 26910 10670 26962
rect 10670 26910 10722 26962
rect 10722 26910 10724 26962
rect 10668 26908 10724 26910
rect 12236 30940 12292 30996
rect 11676 29650 11732 29652
rect 11676 29598 11678 29650
rect 11678 29598 11730 29650
rect 11730 29598 11732 29650
rect 11676 29596 11732 29598
rect 12124 29426 12180 29428
rect 12124 29374 12126 29426
rect 12126 29374 12178 29426
rect 12178 29374 12180 29426
rect 12124 29372 12180 29374
rect 11452 27580 11508 27636
rect 11564 28588 11620 28644
rect 11228 27468 11284 27524
rect 11228 26962 11284 26964
rect 11228 26910 11230 26962
rect 11230 26910 11282 26962
rect 11282 26910 11284 26962
rect 11228 26908 11284 26910
rect 11116 26796 11172 26852
rect 10668 26124 10724 26180
rect 10892 26012 10948 26068
rect 10556 25506 10612 25508
rect 10556 25454 10558 25506
rect 10558 25454 10610 25506
rect 10610 25454 10612 25506
rect 10556 25452 10612 25454
rect 10556 25004 10612 25060
rect 10892 24892 10948 24948
rect 11004 24780 11060 24836
rect 11340 25506 11396 25508
rect 11340 25454 11342 25506
rect 11342 25454 11394 25506
rect 11394 25454 11396 25506
rect 11340 25452 11396 25454
rect 11340 25004 11396 25060
rect 12124 28588 12180 28644
rect 13356 30882 13412 30884
rect 13356 30830 13358 30882
rect 13358 30830 13410 30882
rect 13410 30830 13412 30882
rect 13356 30828 13412 30830
rect 13468 30770 13524 30772
rect 13468 30718 13470 30770
rect 13470 30718 13522 30770
rect 13522 30718 13524 30770
rect 13468 30716 13524 30718
rect 13308 30602 13364 30604
rect 13308 30550 13310 30602
rect 13310 30550 13362 30602
rect 13362 30550 13364 30602
rect 13308 30548 13364 30550
rect 13412 30602 13468 30604
rect 13412 30550 13414 30602
rect 13414 30550 13466 30602
rect 13466 30550 13468 30602
rect 13412 30548 13468 30550
rect 13516 30602 13572 30604
rect 13516 30550 13518 30602
rect 13518 30550 13570 30602
rect 13570 30550 13572 30602
rect 13516 30548 13572 30550
rect 12236 28252 12292 28308
rect 12348 30044 12404 30100
rect 12684 29932 12740 29988
rect 11788 27804 11844 27860
rect 12572 29372 12628 29428
rect 12012 27244 12068 27300
rect 11900 26962 11956 26964
rect 11900 26910 11902 26962
rect 11902 26910 11954 26962
rect 11954 26910 11956 26962
rect 11900 26908 11956 26910
rect 11900 26012 11956 26068
rect 12348 27580 12404 27636
rect 12796 28924 12852 28980
rect 12460 26908 12516 26964
rect 12124 26684 12180 26740
rect 12908 28700 12964 28756
rect 13308 29034 13364 29036
rect 13308 28982 13310 29034
rect 13310 28982 13362 29034
rect 13362 28982 13364 29034
rect 13308 28980 13364 28982
rect 13412 29034 13468 29036
rect 13412 28982 13414 29034
rect 13414 28982 13466 29034
rect 13466 28982 13468 29034
rect 13412 28980 13468 28982
rect 13516 29034 13572 29036
rect 13516 28982 13518 29034
rect 13518 28982 13570 29034
rect 13570 28982 13572 29034
rect 13516 28980 13572 28982
rect 13804 30994 13860 30996
rect 13804 30942 13806 30994
rect 13806 30942 13858 30994
rect 13858 30942 13860 30994
rect 13804 30940 13860 30942
rect 14812 30492 14868 30548
rect 14028 30380 14084 30436
rect 15260 30716 15316 30772
rect 14924 30210 14980 30212
rect 14924 30158 14926 30210
rect 14926 30158 14978 30210
rect 14978 30158 14980 30210
rect 14924 30156 14980 30158
rect 15036 30098 15092 30100
rect 15036 30046 15038 30098
rect 15038 30046 15090 30098
rect 15090 30046 15092 30098
rect 15036 30044 15092 30046
rect 15036 29484 15092 29540
rect 14364 29372 14420 29428
rect 13468 28754 13524 28756
rect 13468 28702 13470 28754
rect 13470 28702 13522 28754
rect 13522 28702 13524 28754
rect 13468 28700 13524 28702
rect 14140 29148 14196 29204
rect 13132 28476 13188 28532
rect 13580 28364 13636 28420
rect 13692 28252 13748 28308
rect 13804 28140 13860 28196
rect 14028 28476 14084 28532
rect 13692 27916 13748 27972
rect 13308 27466 13364 27468
rect 13308 27414 13310 27466
rect 13310 27414 13362 27466
rect 13362 27414 13364 27466
rect 13308 27412 13364 27414
rect 13412 27466 13468 27468
rect 13412 27414 13414 27466
rect 13414 27414 13466 27466
rect 13466 27414 13468 27466
rect 13412 27412 13468 27414
rect 13516 27466 13572 27468
rect 13516 27414 13518 27466
rect 13518 27414 13570 27466
rect 13570 27414 13572 27466
rect 13516 27412 13572 27414
rect 12908 27298 12964 27300
rect 12908 27246 12910 27298
rect 12910 27246 12962 27298
rect 12962 27246 12964 27298
rect 12908 27244 12964 27246
rect 13468 26962 13524 26964
rect 13468 26910 13470 26962
rect 13470 26910 13522 26962
rect 13522 26910 13524 26962
rect 13468 26908 13524 26910
rect 12572 26514 12628 26516
rect 12572 26462 12574 26514
rect 12574 26462 12626 26514
rect 12626 26462 12628 26514
rect 12572 26460 12628 26462
rect 11676 25394 11732 25396
rect 11676 25342 11678 25394
rect 11678 25342 11730 25394
rect 11730 25342 11732 25394
rect 11676 25340 11732 25342
rect 10444 24108 10500 24164
rect 10668 23826 10724 23828
rect 10668 23774 10670 23826
rect 10670 23774 10722 23826
rect 10722 23774 10724 23826
rect 10668 23772 10724 23774
rect 10332 22540 10388 22596
rect 10108 20914 10164 20916
rect 10108 20862 10110 20914
rect 10110 20862 10162 20914
rect 10162 20862 10164 20914
rect 10108 20860 10164 20862
rect 10332 20188 10388 20244
rect 11228 23714 11284 23716
rect 11228 23662 11230 23714
rect 11230 23662 11282 23714
rect 11282 23662 11284 23714
rect 11228 23660 11284 23662
rect 10892 23100 10948 23156
rect 11564 23826 11620 23828
rect 11564 23774 11566 23826
rect 11566 23774 11618 23826
rect 11618 23774 11620 23826
rect 11564 23772 11620 23774
rect 12572 26236 12628 26292
rect 12348 26124 12404 26180
rect 12236 26012 12292 26068
rect 11900 25116 11956 25172
rect 12460 25452 12516 25508
rect 11900 24332 11956 24388
rect 13804 26572 13860 26628
rect 14700 28812 14756 28868
rect 14140 27356 14196 27412
rect 14252 27244 14308 27300
rect 15036 28700 15092 28756
rect 15148 28082 15204 28084
rect 15148 28030 15150 28082
rect 15150 28030 15202 28082
rect 15202 28030 15204 28082
rect 15148 28028 15204 28030
rect 14812 27356 14868 27412
rect 14252 27020 14308 27076
rect 14812 26962 14868 26964
rect 14812 26910 14814 26962
rect 14814 26910 14866 26962
rect 14866 26910 14868 26962
rect 14812 26908 14868 26910
rect 14140 26684 14196 26740
rect 14028 26236 14084 26292
rect 12684 25788 12740 25844
rect 13308 25898 13364 25900
rect 13308 25846 13310 25898
rect 13310 25846 13362 25898
rect 13362 25846 13364 25898
rect 13308 25844 13364 25846
rect 13412 25898 13468 25900
rect 13412 25846 13414 25898
rect 13414 25846 13466 25898
rect 13466 25846 13468 25898
rect 13412 25844 13468 25846
rect 13516 25898 13572 25900
rect 13516 25846 13518 25898
rect 13518 25846 13570 25898
rect 13570 25846 13572 25898
rect 13516 25844 13572 25846
rect 13916 25788 13972 25844
rect 12684 25564 12740 25620
rect 12572 24946 12628 24948
rect 12572 24894 12574 24946
rect 12574 24894 12626 24946
rect 12626 24894 12628 24946
rect 12572 24892 12628 24894
rect 13244 25004 13300 25060
rect 13020 24892 13076 24948
rect 13356 24946 13412 24948
rect 13356 24894 13358 24946
rect 13358 24894 13410 24946
rect 13410 24894 13412 24946
rect 13356 24892 13412 24894
rect 13468 24834 13524 24836
rect 13468 24782 13470 24834
rect 13470 24782 13522 24834
rect 13522 24782 13524 24834
rect 13468 24780 13524 24782
rect 12348 24108 12404 24164
rect 12236 23714 12292 23716
rect 12236 23662 12238 23714
rect 12238 23662 12290 23714
rect 12290 23662 12292 23714
rect 12236 23660 12292 23662
rect 11788 23436 11844 23492
rect 11676 23212 11732 23268
rect 12236 23436 12292 23492
rect 11564 23154 11620 23156
rect 11564 23102 11566 23154
rect 11566 23102 11618 23154
rect 11618 23102 11620 23154
rect 11564 23100 11620 23102
rect 11452 22876 11508 22932
rect 11116 21586 11172 21588
rect 11116 21534 11118 21586
rect 11118 21534 11170 21586
rect 11170 21534 11172 21586
rect 11116 21532 11172 21534
rect 10892 20076 10948 20132
rect 10780 19852 10836 19908
rect 9660 18508 9716 18564
rect 8540 17554 8596 17556
rect 8540 17502 8542 17554
rect 8542 17502 8594 17554
rect 8594 17502 8596 17554
rect 8540 17500 8596 17502
rect 7868 16994 7924 16996
rect 7868 16942 7870 16994
rect 7870 16942 7922 16994
rect 7922 16942 7924 16994
rect 7868 16940 7924 16942
rect 7308 14252 7364 14308
rect 7196 14140 7252 14196
rect 6748 12796 6804 12852
rect 3724 11004 3780 11060
rect 2828 10556 2884 10612
rect 3276 9660 3332 9716
rect 1708 8764 1764 8820
rect 2156 8316 2212 8372
rect 1820 8258 1876 8260
rect 1820 8206 1822 8258
rect 1822 8206 1874 8258
rect 1874 8206 1876 8258
rect 1820 8204 1876 8206
rect 2044 7868 2100 7924
rect 2716 8316 2772 8372
rect 2156 7644 2212 7700
rect 2492 7586 2548 7588
rect 2492 7534 2494 7586
rect 2494 7534 2546 7586
rect 2546 7534 2548 7586
rect 2492 7532 2548 7534
rect 1708 5404 1764 5460
rect 2044 5404 2100 5460
rect 1932 5010 1988 5012
rect 1932 4958 1934 5010
rect 1934 4958 1986 5010
rect 1986 4958 1988 5010
rect 1932 4956 1988 4958
rect 924 3500 980 3556
rect 3164 8092 3220 8148
rect 2604 7196 2660 7252
rect 2380 6524 2436 6580
rect 2380 5404 2436 5460
rect 2268 5292 2324 5348
rect 2044 3388 2100 3444
rect 2156 3330 2212 3332
rect 2156 3278 2158 3330
rect 2158 3278 2210 3330
rect 2210 3278 2212 3330
rect 2156 3276 2212 3278
rect 4508 10834 4564 10836
rect 4508 10782 4510 10834
rect 4510 10782 4562 10834
rect 4562 10782 4564 10834
rect 4508 10780 4564 10782
rect 3724 10610 3780 10612
rect 3724 10558 3726 10610
rect 3726 10558 3778 10610
rect 3778 10558 3780 10610
rect 3724 10556 3780 10558
rect 5964 10834 6020 10836
rect 5964 10782 5966 10834
rect 5966 10782 6018 10834
rect 6018 10782 6020 10834
rect 5964 10780 6020 10782
rect 5404 10386 5460 10388
rect 5404 10334 5406 10386
rect 5406 10334 5458 10386
rect 5458 10334 5460 10386
rect 5404 10332 5460 10334
rect 5244 10218 5300 10220
rect 5244 10166 5246 10218
rect 5246 10166 5298 10218
rect 5298 10166 5300 10218
rect 5244 10164 5300 10166
rect 5348 10218 5404 10220
rect 5348 10166 5350 10218
rect 5350 10166 5402 10218
rect 5402 10166 5404 10218
rect 5348 10164 5404 10166
rect 5452 10218 5508 10220
rect 5452 10166 5454 10218
rect 5454 10166 5506 10218
rect 5506 10166 5508 10218
rect 5452 10164 5508 10166
rect 4844 9996 4900 10052
rect 5516 9996 5572 10052
rect 4060 9602 4116 9604
rect 4060 9550 4062 9602
rect 4062 9550 4114 9602
rect 4114 9550 4116 9602
rect 4060 9548 4116 9550
rect 3500 8876 3556 8932
rect 3948 8652 4004 8708
rect 4956 9548 5012 9604
rect 4620 9100 4676 9156
rect 4284 8764 4340 8820
rect 3836 7868 3892 7924
rect 3836 6860 3892 6916
rect 5068 8930 5124 8932
rect 5068 8878 5070 8930
rect 5070 8878 5122 8930
rect 5122 8878 5124 8930
rect 5068 8876 5124 8878
rect 4508 8204 4564 8260
rect 4396 7980 4452 8036
rect 4172 7698 4228 7700
rect 4172 7646 4174 7698
rect 4174 7646 4226 7698
rect 4226 7646 4228 7698
rect 4172 7644 4228 7646
rect 4284 7474 4340 7476
rect 4284 7422 4286 7474
rect 4286 7422 4338 7474
rect 4338 7422 4340 7474
rect 4284 7420 4340 7422
rect 4396 7196 4452 7252
rect 3836 6412 3892 6468
rect 3836 5628 3892 5684
rect 4620 8764 4676 8820
rect 5740 9826 5796 9828
rect 5740 9774 5742 9826
rect 5742 9774 5794 9826
rect 5794 9774 5796 9826
rect 5740 9772 5796 9774
rect 6076 9602 6132 9604
rect 6076 9550 6078 9602
rect 6078 9550 6130 9602
rect 6130 9550 6132 9602
rect 6076 9548 6132 9550
rect 6412 11340 6468 11396
rect 6412 10834 6468 10836
rect 6412 10782 6414 10834
rect 6414 10782 6466 10834
rect 6466 10782 6468 10834
rect 6412 10780 6468 10782
rect 8428 16994 8484 16996
rect 8428 16942 8430 16994
rect 8430 16942 8482 16994
rect 8482 16942 8484 16994
rect 8428 16940 8484 16942
rect 7532 15148 7588 15204
rect 7644 14530 7700 14532
rect 7644 14478 7646 14530
rect 7646 14478 7698 14530
rect 7698 14478 7700 14530
rect 7644 14476 7700 14478
rect 7980 15314 8036 15316
rect 7980 15262 7982 15314
rect 7982 15262 8034 15314
rect 8034 15262 8036 15314
rect 7980 15260 8036 15262
rect 8316 15426 8372 15428
rect 8316 15374 8318 15426
rect 8318 15374 8370 15426
rect 8370 15374 8372 15426
rect 8316 15372 8372 15374
rect 7868 14140 7924 14196
rect 9276 17274 9332 17276
rect 9276 17222 9278 17274
rect 9278 17222 9330 17274
rect 9330 17222 9332 17274
rect 9276 17220 9332 17222
rect 9380 17274 9436 17276
rect 9380 17222 9382 17274
rect 9382 17222 9434 17274
rect 9434 17222 9436 17274
rect 9380 17220 9436 17222
rect 9484 17274 9540 17276
rect 9484 17222 9486 17274
rect 9486 17222 9538 17274
rect 9538 17222 9540 17274
rect 9484 17220 9540 17222
rect 12012 23100 12068 23156
rect 11452 21980 11508 22036
rect 12348 23266 12404 23268
rect 12348 23214 12350 23266
rect 12350 23214 12402 23266
rect 12402 23214 12404 23266
rect 12348 23212 12404 23214
rect 12236 21644 12292 21700
rect 11228 20524 11284 20580
rect 11116 20412 11172 20468
rect 11564 20412 11620 20468
rect 11004 19068 11060 19124
rect 11452 20076 11508 20132
rect 11564 19122 11620 19124
rect 11564 19070 11566 19122
rect 11566 19070 11618 19122
rect 11618 19070 11620 19122
rect 11564 19068 11620 19070
rect 11676 18956 11732 19012
rect 13308 24330 13364 24332
rect 13308 24278 13310 24330
rect 13310 24278 13362 24330
rect 13362 24278 13364 24330
rect 13308 24276 13364 24278
rect 13412 24330 13468 24332
rect 13412 24278 13414 24330
rect 13414 24278 13466 24330
rect 13466 24278 13468 24330
rect 13412 24276 13468 24278
rect 13516 24330 13572 24332
rect 13516 24278 13518 24330
rect 13518 24278 13570 24330
rect 13570 24278 13572 24330
rect 13516 24276 13572 24278
rect 13804 24668 13860 24724
rect 13916 24444 13972 24500
rect 13804 24220 13860 24276
rect 12684 22988 12740 23044
rect 14140 25676 14196 25732
rect 14252 25506 14308 25508
rect 14252 25454 14254 25506
rect 14254 25454 14306 25506
rect 14306 25454 14308 25506
rect 14252 25452 14308 25454
rect 14700 26850 14756 26852
rect 14700 26798 14702 26850
rect 14702 26798 14754 26850
rect 14754 26798 14756 26850
rect 14700 26796 14756 26798
rect 14588 25676 14644 25732
rect 14812 26684 14868 26740
rect 14588 25340 14644 25396
rect 14476 24892 14532 24948
rect 14140 24668 14196 24724
rect 14364 24332 14420 24388
rect 12908 22428 12964 22484
rect 12908 21756 12964 21812
rect 13692 23100 13748 23156
rect 13308 22762 13364 22764
rect 13308 22710 13310 22762
rect 13310 22710 13362 22762
rect 13362 22710 13364 22762
rect 13308 22708 13364 22710
rect 13412 22762 13468 22764
rect 13412 22710 13414 22762
rect 13414 22710 13466 22762
rect 13466 22710 13468 22762
rect 13412 22708 13468 22710
rect 13516 22762 13572 22764
rect 13516 22710 13518 22762
rect 13518 22710 13570 22762
rect 13570 22710 13572 22762
rect 13516 22708 13572 22710
rect 13580 22540 13636 22596
rect 12572 21644 12628 21700
rect 12460 21420 12516 21476
rect 12124 18844 12180 18900
rect 12236 20524 12292 20580
rect 11788 18674 11844 18676
rect 11788 18622 11790 18674
rect 11790 18622 11842 18674
rect 11842 18622 11844 18674
rect 11788 18620 11844 18622
rect 12012 18620 12068 18676
rect 9884 18284 9940 18340
rect 11116 18450 11172 18452
rect 11116 18398 11118 18450
rect 11118 18398 11170 18450
rect 11170 18398 11172 18450
rect 11116 18396 11172 18398
rect 12012 18450 12068 18452
rect 12012 18398 12014 18450
rect 12014 18398 12066 18450
rect 12066 18398 12068 18450
rect 12012 18396 12068 18398
rect 11228 18338 11284 18340
rect 11228 18286 11230 18338
rect 11230 18286 11282 18338
rect 11282 18286 11284 18338
rect 11228 18284 11284 18286
rect 10892 18172 10948 18228
rect 10668 17388 10724 17444
rect 11340 17612 11396 17668
rect 10892 16098 10948 16100
rect 10892 16046 10894 16098
rect 10894 16046 10946 16098
rect 10946 16046 10948 16098
rect 10892 16044 10948 16046
rect 14140 23660 14196 23716
rect 13804 22428 13860 22484
rect 14252 23100 14308 23156
rect 13692 21868 13748 21924
rect 14028 22092 14084 22148
rect 13580 21756 13636 21812
rect 13468 21532 13524 21588
rect 13308 21194 13364 21196
rect 13308 21142 13310 21194
rect 13310 21142 13362 21194
rect 13362 21142 13364 21194
rect 13308 21140 13364 21142
rect 13412 21194 13468 21196
rect 13412 21142 13414 21194
rect 13414 21142 13466 21194
rect 13466 21142 13468 21194
rect 13412 21140 13468 21142
rect 13516 21194 13572 21196
rect 13516 21142 13518 21194
rect 13518 21142 13570 21194
rect 13570 21142 13572 21194
rect 13516 21140 13572 21142
rect 13804 20972 13860 21028
rect 13468 20860 13524 20916
rect 12572 20076 12628 20132
rect 13692 20130 13748 20132
rect 13692 20078 13694 20130
rect 13694 20078 13746 20130
rect 13746 20078 13748 20130
rect 13692 20076 13748 20078
rect 12908 19964 12964 20020
rect 13308 19626 13364 19628
rect 13308 19574 13310 19626
rect 13310 19574 13362 19626
rect 13362 19574 13364 19626
rect 13308 19572 13364 19574
rect 13412 19626 13468 19628
rect 13412 19574 13414 19626
rect 13414 19574 13466 19626
rect 13466 19574 13468 19626
rect 13412 19572 13468 19574
rect 13516 19626 13572 19628
rect 13516 19574 13518 19626
rect 13518 19574 13570 19626
rect 13570 19574 13572 19626
rect 13516 19572 13572 19574
rect 12908 19346 12964 19348
rect 12908 19294 12910 19346
rect 12910 19294 12962 19346
rect 12962 19294 12964 19346
rect 12908 19292 12964 19294
rect 12236 17500 12292 17556
rect 12348 19068 12404 19124
rect 12460 17612 12516 17668
rect 13020 19068 13076 19124
rect 13692 18844 13748 18900
rect 13132 18674 13188 18676
rect 13132 18622 13134 18674
rect 13134 18622 13186 18674
rect 13186 18622 13188 18674
rect 13132 18620 13188 18622
rect 15372 30492 15428 30548
rect 16492 30380 16548 30436
rect 16940 29932 16996 29988
rect 15932 29596 15988 29652
rect 15708 29484 15764 29540
rect 16492 29596 16548 29652
rect 15708 29148 15764 29204
rect 16156 29426 16212 29428
rect 16156 29374 16158 29426
rect 16158 29374 16210 29426
rect 16210 29374 16212 29426
rect 16156 29372 16212 29374
rect 15820 28812 15876 28868
rect 16044 29036 16100 29092
rect 15484 28642 15540 28644
rect 15484 28590 15486 28642
rect 15486 28590 15538 28642
rect 15538 28590 15540 28642
rect 15484 28588 15540 28590
rect 15260 26460 15316 26516
rect 15372 26012 15428 26068
rect 15148 25900 15204 25956
rect 15372 25788 15428 25844
rect 15260 25564 15316 25620
rect 15036 25340 15092 25396
rect 15148 24780 15204 24836
rect 14588 22428 14644 22484
rect 14700 23324 14756 23380
rect 14476 22258 14532 22260
rect 14476 22206 14478 22258
rect 14478 22206 14530 22258
rect 14530 22206 14532 22258
rect 14476 22204 14532 22206
rect 15036 24220 15092 24276
rect 14812 22876 14868 22932
rect 14924 24108 14980 24164
rect 14812 22652 14868 22708
rect 14700 22092 14756 22148
rect 15036 23884 15092 23940
rect 15036 23100 15092 23156
rect 15484 25116 15540 25172
rect 15708 25564 15764 25620
rect 15820 26908 15876 26964
rect 15932 26684 15988 26740
rect 15932 25676 15988 25732
rect 16492 29036 16548 29092
rect 16828 28476 16884 28532
rect 17340 31386 17396 31388
rect 17340 31334 17342 31386
rect 17342 31334 17394 31386
rect 17394 31334 17396 31386
rect 17340 31332 17396 31334
rect 17444 31386 17500 31388
rect 17444 31334 17446 31386
rect 17446 31334 17498 31386
rect 17498 31334 17500 31386
rect 17444 31332 17500 31334
rect 17548 31386 17604 31388
rect 17548 31334 17550 31386
rect 17550 31334 17602 31386
rect 17602 31334 17604 31386
rect 17548 31332 17604 31334
rect 20636 33068 20692 33124
rect 20748 32060 20804 32116
rect 19516 31164 19572 31220
rect 19628 31948 19684 32004
rect 19628 31500 19684 31556
rect 17276 29932 17332 29988
rect 17836 30156 17892 30212
rect 17340 29818 17396 29820
rect 17340 29766 17342 29818
rect 17342 29766 17394 29818
rect 17394 29766 17396 29818
rect 17340 29764 17396 29766
rect 17444 29818 17500 29820
rect 17444 29766 17446 29818
rect 17446 29766 17498 29818
rect 17498 29766 17500 29818
rect 17444 29764 17500 29766
rect 17548 29818 17604 29820
rect 17548 29766 17550 29818
rect 17550 29766 17602 29818
rect 17602 29766 17604 29818
rect 17548 29764 17604 29766
rect 17836 29260 17892 29316
rect 17388 29036 17444 29092
rect 17500 28364 17556 28420
rect 17724 28924 17780 28980
rect 17340 28250 17396 28252
rect 17340 28198 17342 28250
rect 17342 28198 17394 28250
rect 17394 28198 17396 28250
rect 17340 28196 17396 28198
rect 17444 28250 17500 28252
rect 17444 28198 17446 28250
rect 17446 28198 17498 28250
rect 17498 28198 17500 28250
rect 17444 28196 17500 28198
rect 17548 28250 17604 28252
rect 17548 28198 17550 28250
rect 17550 28198 17602 28250
rect 17602 28198 17604 28250
rect 17548 28196 17604 28198
rect 17276 28028 17332 28084
rect 17052 27804 17108 27860
rect 17052 27020 17108 27076
rect 17340 26682 17396 26684
rect 17340 26630 17342 26682
rect 17342 26630 17394 26682
rect 17394 26630 17396 26682
rect 17340 26628 17396 26630
rect 17444 26682 17500 26684
rect 17444 26630 17446 26682
rect 17446 26630 17498 26682
rect 17498 26630 17500 26682
rect 17444 26628 17500 26630
rect 17548 26682 17604 26684
rect 17548 26630 17550 26682
rect 17550 26630 17602 26682
rect 17602 26630 17604 26682
rect 17548 26628 17604 26630
rect 17052 26460 17108 26516
rect 16156 26124 16212 26180
rect 16604 26178 16660 26180
rect 16604 26126 16606 26178
rect 16606 26126 16658 26178
rect 16658 26126 16660 26178
rect 16604 26124 16660 26126
rect 16156 25900 16212 25956
rect 15260 24556 15316 24612
rect 15260 24220 15316 24276
rect 15932 24722 15988 24724
rect 15932 24670 15934 24722
rect 15934 24670 15986 24722
rect 15986 24670 15988 24722
rect 15932 24668 15988 24670
rect 16940 25900 16996 25956
rect 16380 25452 16436 25508
rect 16268 25116 16324 25172
rect 16268 24834 16324 24836
rect 16268 24782 16270 24834
rect 16270 24782 16322 24834
rect 16322 24782 16324 24834
rect 16268 24780 16324 24782
rect 16828 25340 16884 25396
rect 16716 24834 16772 24836
rect 16716 24782 16718 24834
rect 16718 24782 16770 24834
rect 16770 24782 16772 24834
rect 16716 24780 16772 24782
rect 16828 24556 16884 24612
rect 15372 23996 15428 24052
rect 16604 23996 16660 24052
rect 15148 22540 15204 22596
rect 15708 23324 15764 23380
rect 15820 22930 15876 22932
rect 15820 22878 15822 22930
rect 15822 22878 15874 22930
rect 15874 22878 15876 22930
rect 15820 22876 15876 22878
rect 15708 22764 15764 22820
rect 15036 21980 15092 22036
rect 14364 21810 14420 21812
rect 14364 21758 14366 21810
rect 14366 21758 14418 21810
rect 14418 21758 14420 21810
rect 14364 21756 14420 21758
rect 15820 21868 15876 21924
rect 14252 20860 14308 20916
rect 14476 20076 14532 20132
rect 14364 20018 14420 20020
rect 14364 19966 14366 20018
rect 14366 19966 14418 20018
rect 14418 19966 14420 20018
rect 14364 19964 14420 19966
rect 14140 19292 14196 19348
rect 13916 18732 13972 18788
rect 13804 18620 13860 18676
rect 13916 18450 13972 18452
rect 13916 18398 13918 18450
rect 13918 18398 13970 18450
rect 13970 18398 13972 18450
rect 13916 18396 13972 18398
rect 13308 18058 13364 18060
rect 13308 18006 13310 18058
rect 13310 18006 13362 18058
rect 13362 18006 13364 18058
rect 13308 18004 13364 18006
rect 13412 18058 13468 18060
rect 13412 18006 13414 18058
rect 13414 18006 13466 18058
rect 13466 18006 13468 18058
rect 13412 18004 13468 18006
rect 13516 18058 13572 18060
rect 13516 18006 13518 18058
rect 13518 18006 13570 18058
rect 13570 18006 13572 18058
rect 13516 18004 13572 18006
rect 14028 18172 14084 18228
rect 12908 17612 12964 17668
rect 13580 17666 13636 17668
rect 13580 17614 13582 17666
rect 13582 17614 13634 17666
rect 13634 17614 13636 17666
rect 13580 17612 13636 17614
rect 14476 18620 14532 18676
rect 14476 18172 14532 18228
rect 11788 17164 11844 17220
rect 11564 16882 11620 16884
rect 11564 16830 11566 16882
rect 11566 16830 11618 16882
rect 11618 16830 11620 16882
rect 11564 16828 11620 16830
rect 12684 17164 12740 17220
rect 12572 16940 12628 16996
rect 11676 16098 11732 16100
rect 11676 16046 11678 16098
rect 11678 16046 11730 16098
rect 11730 16046 11732 16098
rect 11676 16044 11732 16046
rect 12460 16828 12516 16884
rect 9276 15706 9332 15708
rect 9276 15654 9278 15706
rect 9278 15654 9330 15706
rect 9330 15654 9332 15706
rect 9276 15652 9332 15654
rect 9380 15706 9436 15708
rect 9380 15654 9382 15706
rect 9382 15654 9434 15706
rect 9434 15654 9436 15706
rect 9380 15652 9436 15654
rect 9484 15706 9540 15708
rect 9484 15654 9486 15706
rect 9486 15654 9538 15706
rect 9538 15654 9540 15706
rect 9484 15652 9540 15654
rect 8540 14476 8596 14532
rect 8652 15372 8708 15428
rect 10220 15426 10276 15428
rect 10220 15374 10222 15426
rect 10222 15374 10274 15426
rect 10274 15374 10276 15426
rect 10220 15372 10276 15374
rect 10556 15314 10612 15316
rect 10556 15262 10558 15314
rect 10558 15262 10610 15314
rect 10610 15262 10612 15314
rect 10556 15260 10612 15262
rect 10556 14924 10612 14980
rect 8540 14306 8596 14308
rect 8540 14254 8542 14306
rect 8542 14254 8594 14306
rect 8594 14254 8596 14306
rect 8540 14252 8596 14254
rect 9276 14138 9332 14140
rect 9276 14086 9278 14138
rect 9278 14086 9330 14138
rect 9330 14086 9332 14138
rect 9276 14084 9332 14086
rect 9380 14138 9436 14140
rect 9380 14086 9382 14138
rect 9382 14086 9434 14138
rect 9434 14086 9436 14138
rect 9380 14084 9436 14086
rect 9484 14138 9540 14140
rect 9484 14086 9486 14138
rect 9486 14086 9538 14138
rect 9538 14086 9540 14138
rect 9484 14084 9540 14086
rect 8988 13916 9044 13972
rect 11228 15314 11284 15316
rect 11228 15262 11230 15314
rect 11230 15262 11282 15314
rect 11282 15262 11284 15314
rect 11228 15260 11284 15262
rect 11340 14924 11396 14980
rect 11452 15260 11508 15316
rect 10780 13970 10836 13972
rect 10780 13918 10782 13970
rect 10782 13918 10834 13970
rect 10834 13918 10836 13970
rect 10780 13916 10836 13918
rect 8540 12962 8596 12964
rect 8540 12910 8542 12962
rect 8542 12910 8594 12962
rect 8594 12910 8596 12962
rect 8540 12908 8596 12910
rect 9212 12908 9268 12964
rect 7756 12850 7812 12852
rect 7756 12798 7758 12850
rect 7758 12798 7810 12850
rect 7810 12798 7812 12850
rect 7756 12796 7812 12798
rect 7532 12012 7588 12068
rect 8092 12066 8148 12068
rect 8092 12014 8094 12066
rect 8094 12014 8146 12066
rect 8146 12014 8148 12066
rect 8092 12012 8148 12014
rect 7644 11004 7700 11060
rect 7868 11452 7924 11508
rect 6412 9826 6468 9828
rect 6412 9774 6414 9826
rect 6414 9774 6466 9826
rect 6466 9774 6468 9826
rect 6412 9772 6468 9774
rect 6188 9100 6244 9156
rect 5180 8764 5236 8820
rect 5244 8650 5300 8652
rect 5244 8598 5246 8650
rect 5246 8598 5298 8650
rect 5298 8598 5300 8650
rect 5244 8596 5300 8598
rect 5348 8650 5404 8652
rect 5348 8598 5350 8650
rect 5350 8598 5402 8650
rect 5402 8598 5404 8650
rect 5348 8596 5404 8598
rect 5452 8650 5508 8652
rect 5452 8598 5454 8650
rect 5454 8598 5506 8650
rect 5506 8598 5508 8650
rect 5452 8596 5508 8598
rect 5740 8146 5796 8148
rect 5740 8094 5742 8146
rect 5742 8094 5794 8146
rect 5794 8094 5796 8146
rect 5740 8092 5796 8094
rect 5180 7868 5236 7924
rect 5516 7756 5572 7812
rect 4956 7644 5012 7700
rect 4844 7196 4900 7252
rect 4844 6524 4900 6580
rect 5244 7082 5300 7084
rect 5244 7030 5246 7082
rect 5246 7030 5298 7082
rect 5298 7030 5300 7082
rect 5244 7028 5300 7030
rect 5348 7082 5404 7084
rect 5348 7030 5350 7082
rect 5350 7030 5402 7082
rect 5402 7030 5404 7082
rect 5348 7028 5404 7030
rect 5452 7082 5508 7084
rect 5452 7030 5454 7082
rect 5454 7030 5506 7082
rect 5506 7030 5508 7082
rect 5452 7028 5508 7030
rect 5516 6748 5572 6804
rect 5180 6076 5236 6132
rect 5292 6188 5348 6244
rect 5068 6018 5124 6020
rect 5068 5966 5070 6018
rect 5070 5966 5122 6018
rect 5122 5966 5124 6018
rect 5068 5964 5124 5966
rect 5244 5514 5300 5516
rect 5244 5462 5246 5514
rect 5246 5462 5298 5514
rect 5298 5462 5300 5514
rect 5244 5460 5300 5462
rect 5348 5514 5404 5516
rect 5348 5462 5350 5514
rect 5350 5462 5402 5514
rect 5402 5462 5404 5514
rect 5348 5460 5404 5462
rect 5452 5514 5508 5516
rect 5452 5462 5454 5514
rect 5454 5462 5506 5514
rect 5506 5462 5508 5514
rect 5452 5460 5508 5462
rect 5964 7644 6020 7700
rect 6188 8316 6244 8372
rect 6076 7474 6132 7476
rect 6076 7422 6078 7474
rect 6078 7422 6130 7474
rect 6130 7422 6132 7474
rect 6076 7420 6132 7422
rect 5964 7308 6020 7364
rect 5852 6690 5908 6692
rect 5852 6638 5854 6690
rect 5854 6638 5906 6690
rect 5906 6638 5908 6690
rect 5852 6636 5908 6638
rect 5740 6412 5796 6468
rect 5628 5292 5684 5348
rect 5740 6076 5796 6132
rect 6300 7532 6356 7588
rect 5964 5180 6020 5236
rect 6076 5068 6132 5124
rect 5244 3946 5300 3948
rect 5244 3894 5246 3946
rect 5246 3894 5298 3946
rect 5298 3894 5300 3946
rect 5244 3892 5300 3894
rect 5348 3946 5404 3948
rect 5348 3894 5350 3946
rect 5350 3894 5402 3946
rect 5402 3894 5404 3946
rect 5348 3892 5404 3894
rect 5452 3946 5508 3948
rect 5452 3894 5454 3946
rect 5454 3894 5506 3946
rect 5506 3894 5508 3946
rect 5452 3892 5508 3894
rect 3276 3500 3332 3556
rect 3164 3276 3220 3332
rect 5516 3330 5572 3332
rect 5516 3278 5518 3330
rect 5518 3278 5570 3330
rect 5570 3278 5572 3330
rect 5516 3276 5572 3278
rect 8652 11452 8708 11508
rect 8428 11340 8484 11396
rect 8204 10780 8260 10836
rect 7196 9996 7252 10052
rect 7084 9826 7140 9828
rect 7084 9774 7086 9826
rect 7086 9774 7138 9826
rect 7138 9774 7140 9826
rect 7084 9772 7140 9774
rect 6748 9714 6804 9716
rect 6748 9662 6750 9714
rect 6750 9662 6802 9714
rect 6802 9662 6804 9714
rect 6748 9660 6804 9662
rect 7420 9714 7476 9716
rect 7420 9662 7422 9714
rect 7422 9662 7474 9714
rect 7474 9662 7476 9714
rect 7420 9660 7476 9662
rect 7308 9324 7364 9380
rect 7532 9548 7588 9604
rect 6748 7980 6804 8036
rect 6748 7474 6804 7476
rect 6748 7422 6750 7474
rect 6750 7422 6802 7474
rect 6802 7422 6804 7474
rect 6748 7420 6804 7422
rect 6524 6860 6580 6916
rect 6300 5628 6356 5684
rect 6412 6636 6468 6692
rect 6412 5180 6468 5236
rect 6972 7308 7028 7364
rect 6860 6748 6916 6804
rect 7980 9602 8036 9604
rect 7980 9550 7982 9602
rect 7982 9550 8034 9602
rect 8034 9550 8036 9602
rect 7980 9548 8036 9550
rect 7756 9324 7812 9380
rect 7868 8316 7924 8372
rect 8316 11004 8372 11060
rect 8316 9714 8372 9716
rect 8316 9662 8318 9714
rect 8318 9662 8370 9714
rect 8370 9662 8372 9714
rect 8316 9660 8372 9662
rect 8988 11506 9044 11508
rect 8988 11454 8990 11506
rect 8990 11454 9042 11506
rect 9042 11454 9044 11506
rect 8988 11452 9044 11454
rect 8652 10834 8708 10836
rect 8652 10782 8654 10834
rect 8654 10782 8706 10834
rect 8706 10782 8708 10834
rect 8652 10780 8708 10782
rect 9996 12962 10052 12964
rect 9996 12910 9998 12962
rect 9998 12910 10050 12962
rect 10050 12910 10052 12962
rect 9996 12908 10052 12910
rect 9276 12570 9332 12572
rect 9276 12518 9278 12570
rect 9278 12518 9330 12570
rect 9330 12518 9332 12570
rect 9276 12516 9332 12518
rect 9380 12570 9436 12572
rect 9380 12518 9382 12570
rect 9382 12518 9434 12570
rect 9434 12518 9436 12570
rect 9380 12516 9436 12518
rect 9484 12570 9540 12572
rect 9484 12518 9486 12570
rect 9486 12518 9538 12570
rect 9538 12518 9540 12570
rect 9484 12516 9540 12518
rect 9436 11506 9492 11508
rect 9436 11454 9438 11506
rect 9438 11454 9490 11506
rect 9490 11454 9492 11506
rect 9436 11452 9492 11454
rect 10780 13468 10836 13524
rect 13132 16828 13188 16884
rect 13916 16882 13972 16884
rect 13916 16830 13918 16882
rect 13918 16830 13970 16882
rect 13970 16830 13972 16882
rect 13916 16828 13972 16830
rect 13308 16490 13364 16492
rect 13308 16438 13310 16490
rect 13310 16438 13362 16490
rect 13362 16438 13364 16490
rect 13308 16436 13364 16438
rect 13412 16490 13468 16492
rect 13412 16438 13414 16490
rect 13414 16438 13466 16490
rect 13466 16438 13468 16490
rect 13412 16436 13468 16438
rect 13516 16490 13572 16492
rect 13516 16438 13518 16490
rect 13518 16438 13570 16490
rect 13570 16438 13572 16490
rect 13516 16436 13572 16438
rect 13356 15426 13412 15428
rect 13356 15374 13358 15426
rect 13358 15374 13410 15426
rect 13410 15374 13412 15426
rect 13356 15372 13412 15374
rect 14812 21586 14868 21588
rect 14812 21534 14814 21586
rect 14814 21534 14866 21586
rect 14866 21534 14868 21586
rect 14812 21532 14868 21534
rect 15484 21308 15540 21364
rect 14812 20412 14868 20468
rect 15260 20242 15316 20244
rect 15260 20190 15262 20242
rect 15262 20190 15314 20242
rect 15314 20190 15316 20242
rect 15260 20188 15316 20190
rect 16268 23938 16324 23940
rect 16268 23886 16270 23938
rect 16270 23886 16322 23938
rect 16322 23886 16324 23938
rect 16268 23884 16324 23886
rect 16156 23826 16212 23828
rect 16156 23774 16158 23826
rect 16158 23774 16210 23826
rect 16210 23774 16212 23826
rect 16156 23772 16212 23774
rect 16380 23660 16436 23716
rect 16156 23324 16212 23380
rect 16380 23212 16436 23268
rect 17724 26514 17780 26516
rect 17724 26462 17726 26514
rect 17726 26462 17778 26514
rect 17778 26462 17780 26514
rect 17724 26460 17780 26462
rect 17388 26348 17444 26404
rect 18620 30940 18676 30996
rect 18508 30156 18564 30212
rect 18396 29650 18452 29652
rect 18396 29598 18398 29650
rect 18398 29598 18450 29650
rect 18450 29598 18452 29650
rect 18396 29596 18452 29598
rect 18284 29148 18340 29204
rect 18620 29484 18676 29540
rect 18732 30044 18788 30100
rect 17948 28700 18004 28756
rect 18284 28754 18340 28756
rect 18284 28702 18286 28754
rect 18286 28702 18338 28754
rect 18338 28702 18340 28754
rect 18284 28700 18340 28702
rect 18396 28588 18452 28644
rect 18844 29426 18900 29428
rect 18844 29374 18846 29426
rect 18846 29374 18898 29426
rect 18898 29374 18900 29426
rect 18844 29372 18900 29374
rect 18844 28530 18900 28532
rect 18844 28478 18846 28530
rect 18846 28478 18898 28530
rect 18898 28478 18900 28530
rect 18844 28476 18900 28478
rect 18508 28252 18564 28308
rect 18620 28364 18676 28420
rect 18508 28082 18564 28084
rect 18508 28030 18510 28082
rect 18510 28030 18562 28082
rect 18562 28030 18564 28082
rect 18508 28028 18564 28030
rect 20860 31276 20916 31332
rect 20748 30994 20804 30996
rect 20748 30942 20750 30994
rect 20750 30942 20802 30994
rect 20802 30942 20804 30994
rect 20748 30940 20804 30942
rect 20412 30380 20468 30436
rect 20076 30268 20132 30324
rect 20076 29932 20132 29988
rect 19516 29314 19572 29316
rect 19516 29262 19518 29314
rect 19518 29262 19570 29314
rect 19570 29262 19572 29314
rect 19516 29260 19572 29262
rect 20300 30156 20356 30212
rect 20636 30322 20692 30324
rect 20636 30270 20638 30322
rect 20638 30270 20690 30322
rect 20690 30270 20692 30322
rect 20636 30268 20692 30270
rect 20524 29260 20580 29316
rect 20076 29036 20132 29092
rect 19964 28700 20020 28756
rect 19292 28642 19348 28644
rect 19292 28590 19294 28642
rect 19294 28590 19346 28642
rect 19346 28590 19348 28642
rect 19292 28588 19348 28590
rect 19628 28588 19684 28644
rect 18732 27298 18788 27300
rect 18732 27246 18734 27298
rect 18734 27246 18786 27298
rect 18786 27246 18788 27298
rect 18732 27244 18788 27246
rect 18956 27692 19012 27748
rect 19180 27580 19236 27636
rect 19404 28418 19460 28420
rect 19404 28366 19406 28418
rect 19406 28366 19458 28418
rect 19458 28366 19460 28418
rect 19404 28364 19460 28366
rect 19292 27074 19348 27076
rect 19292 27022 19294 27074
rect 19294 27022 19346 27074
rect 19346 27022 19348 27074
rect 19292 27020 19348 27022
rect 18844 26572 18900 26628
rect 18732 26460 18788 26516
rect 18508 26348 18564 26404
rect 18172 26290 18228 26292
rect 18172 26238 18174 26290
rect 18174 26238 18226 26290
rect 18226 26238 18228 26290
rect 18172 26236 18228 26238
rect 17500 26066 17556 26068
rect 17500 26014 17502 26066
rect 17502 26014 17554 26066
rect 17554 26014 17556 26066
rect 17500 26012 17556 26014
rect 17724 25618 17780 25620
rect 17724 25566 17726 25618
rect 17726 25566 17778 25618
rect 17778 25566 17780 25618
rect 17724 25564 17780 25566
rect 17836 25506 17892 25508
rect 17836 25454 17838 25506
rect 17838 25454 17890 25506
rect 17890 25454 17892 25506
rect 17836 25452 17892 25454
rect 17052 24108 17108 24164
rect 16716 23212 16772 23268
rect 16940 23996 16996 24052
rect 16492 22652 16548 22708
rect 16604 22876 16660 22932
rect 16828 22876 16884 22932
rect 16380 22428 16436 22484
rect 16268 22370 16324 22372
rect 16268 22318 16270 22370
rect 16270 22318 16322 22370
rect 16322 22318 16324 22370
rect 16268 22316 16324 22318
rect 16044 21980 16100 22036
rect 16716 22092 16772 22148
rect 17052 23884 17108 23940
rect 17340 25114 17396 25116
rect 17340 25062 17342 25114
rect 17342 25062 17394 25114
rect 17394 25062 17396 25114
rect 17340 25060 17396 25062
rect 17444 25114 17500 25116
rect 17444 25062 17446 25114
rect 17446 25062 17498 25114
rect 17498 25062 17500 25114
rect 17444 25060 17500 25062
rect 17548 25114 17604 25116
rect 17548 25062 17550 25114
rect 17550 25062 17602 25114
rect 17602 25062 17604 25114
rect 17548 25060 17604 25062
rect 17388 24892 17444 24948
rect 17500 24556 17556 24612
rect 17612 24444 17668 24500
rect 17500 24220 17556 24276
rect 17164 23660 17220 23716
rect 17612 23714 17668 23716
rect 17612 23662 17614 23714
rect 17614 23662 17666 23714
rect 17666 23662 17668 23714
rect 17612 23660 17668 23662
rect 17340 23546 17396 23548
rect 17340 23494 17342 23546
rect 17342 23494 17394 23546
rect 17394 23494 17396 23546
rect 17340 23492 17396 23494
rect 17444 23546 17500 23548
rect 17444 23494 17446 23546
rect 17446 23494 17498 23546
rect 17498 23494 17500 23546
rect 17444 23492 17500 23494
rect 17548 23546 17604 23548
rect 17548 23494 17550 23546
rect 17550 23494 17602 23546
rect 17602 23494 17604 23546
rect 17548 23492 17604 23494
rect 18732 26236 18788 26292
rect 18620 26124 18676 26180
rect 18060 26012 18116 26068
rect 18508 25506 18564 25508
rect 18508 25454 18510 25506
rect 18510 25454 18562 25506
rect 18562 25454 18564 25506
rect 18508 25452 18564 25454
rect 17948 23772 18004 23828
rect 18284 25340 18340 25396
rect 17836 23548 17892 23604
rect 17500 22764 17556 22820
rect 17836 22652 17892 22708
rect 18508 25004 18564 25060
rect 18396 24946 18452 24948
rect 18396 24894 18398 24946
rect 18398 24894 18450 24946
rect 18450 24894 18452 24946
rect 18396 24892 18452 24894
rect 18172 24668 18228 24724
rect 18508 24332 18564 24388
rect 18060 23660 18116 23716
rect 19292 26348 19348 26404
rect 19180 26124 19236 26180
rect 18956 25618 19012 25620
rect 18956 25566 18958 25618
rect 18958 25566 19010 25618
rect 19010 25566 19012 25618
rect 18956 25564 19012 25566
rect 18844 25228 18900 25284
rect 20412 28700 20468 28756
rect 20300 28642 20356 28644
rect 20300 28590 20302 28642
rect 20302 28590 20354 28642
rect 20354 28590 20356 28642
rect 20300 28588 20356 28590
rect 20636 28530 20692 28532
rect 20636 28478 20638 28530
rect 20638 28478 20690 28530
rect 20690 28478 20692 28530
rect 20636 28476 20692 28478
rect 20188 27244 20244 27300
rect 20524 28082 20580 28084
rect 20524 28030 20526 28082
rect 20526 28030 20578 28082
rect 20578 28030 20580 28082
rect 20524 28028 20580 28030
rect 20412 27858 20468 27860
rect 20412 27806 20414 27858
rect 20414 27806 20466 27858
rect 20466 27806 20468 27858
rect 20412 27804 20468 27806
rect 20524 27634 20580 27636
rect 20524 27582 20526 27634
rect 20526 27582 20578 27634
rect 20578 27582 20580 27634
rect 20524 27580 20580 27582
rect 20524 27074 20580 27076
rect 20524 27022 20526 27074
rect 20526 27022 20578 27074
rect 20578 27022 20580 27074
rect 20524 27020 20580 27022
rect 20412 26908 20468 26964
rect 20972 31052 21028 31108
rect 20860 28812 20916 28868
rect 20972 29372 21028 29428
rect 20860 28476 20916 28532
rect 20860 27804 20916 27860
rect 21084 28476 21140 28532
rect 21756 31218 21812 31220
rect 21756 31166 21758 31218
rect 21758 31166 21810 31218
rect 21810 31166 21812 31218
rect 21756 31164 21812 31166
rect 22876 31164 22932 31220
rect 23884 33404 23940 33460
rect 23884 31612 23940 31668
rect 23660 31106 23716 31108
rect 23660 31054 23662 31106
rect 23662 31054 23714 31106
rect 23714 31054 23716 31106
rect 23660 31052 23716 31054
rect 21868 30716 21924 30772
rect 21372 30602 21428 30604
rect 21372 30550 21374 30602
rect 21374 30550 21426 30602
rect 21426 30550 21428 30602
rect 21372 30548 21428 30550
rect 21476 30602 21532 30604
rect 21476 30550 21478 30602
rect 21478 30550 21530 30602
rect 21530 30550 21532 30602
rect 21476 30548 21532 30550
rect 21580 30602 21636 30604
rect 21580 30550 21582 30602
rect 21582 30550 21634 30602
rect 21634 30550 21636 30602
rect 21580 30548 21636 30550
rect 21308 29372 21364 29428
rect 21372 29034 21428 29036
rect 21372 28982 21374 29034
rect 21374 28982 21426 29034
rect 21426 28982 21428 29034
rect 21372 28980 21428 28982
rect 21476 29034 21532 29036
rect 21476 28982 21478 29034
rect 21478 28982 21530 29034
rect 21530 28982 21532 29034
rect 21476 28980 21532 28982
rect 21580 29034 21636 29036
rect 21580 28982 21582 29034
rect 21582 28982 21634 29034
rect 21634 28982 21636 29034
rect 21580 28980 21636 28982
rect 21308 28812 21364 28868
rect 21644 28700 21700 28756
rect 23436 30380 23492 30436
rect 23436 30156 23492 30212
rect 21196 28364 21252 28420
rect 21644 28476 21700 28532
rect 21868 28530 21924 28532
rect 21868 28478 21870 28530
rect 21870 28478 21922 28530
rect 21922 28478 21924 28530
rect 21868 28476 21924 28478
rect 21756 27746 21812 27748
rect 21756 27694 21758 27746
rect 21758 27694 21810 27746
rect 21810 27694 21812 27746
rect 21756 27692 21812 27694
rect 21372 27466 21428 27468
rect 21372 27414 21374 27466
rect 21374 27414 21426 27466
rect 21426 27414 21428 27466
rect 21372 27412 21428 27414
rect 21476 27466 21532 27468
rect 21476 27414 21478 27466
rect 21478 27414 21530 27466
rect 21530 27414 21532 27466
rect 21476 27412 21532 27414
rect 21580 27466 21636 27468
rect 21580 27414 21582 27466
rect 21582 27414 21634 27466
rect 21634 27414 21636 27466
rect 21580 27412 21636 27414
rect 20860 27020 20916 27076
rect 19628 26348 19684 26404
rect 19740 26460 19796 26516
rect 19628 26178 19684 26180
rect 19628 26126 19630 26178
rect 19630 26126 19682 26178
rect 19682 26126 19684 26178
rect 19628 26124 19684 26126
rect 19740 25452 19796 25508
rect 19180 25228 19236 25284
rect 19068 25116 19124 25172
rect 18732 23938 18788 23940
rect 18732 23886 18734 23938
rect 18734 23886 18786 23938
rect 18786 23886 18788 23938
rect 18732 23884 18788 23886
rect 18620 23436 18676 23492
rect 18508 23324 18564 23380
rect 16492 21644 16548 21700
rect 16156 20242 16212 20244
rect 16156 20190 16158 20242
rect 16158 20190 16210 20242
rect 16210 20190 16212 20242
rect 16156 20188 16212 20190
rect 16604 20748 16660 20804
rect 15820 20076 15876 20132
rect 15036 20018 15092 20020
rect 15036 19966 15038 20018
rect 15038 19966 15090 20018
rect 15090 19966 15092 20018
rect 15036 19964 15092 19966
rect 15036 19516 15092 19572
rect 15036 18732 15092 18788
rect 14812 18450 14868 18452
rect 14812 18398 14814 18450
rect 14814 18398 14866 18450
rect 14866 18398 14868 18450
rect 14812 18396 14868 18398
rect 15484 18674 15540 18676
rect 15484 18622 15486 18674
rect 15486 18622 15538 18674
rect 15538 18622 15540 18674
rect 15484 18620 15540 18622
rect 15596 18562 15652 18564
rect 15596 18510 15598 18562
rect 15598 18510 15650 18562
rect 15650 18510 15652 18562
rect 15596 18508 15652 18510
rect 16156 19068 16212 19124
rect 15260 18450 15316 18452
rect 15260 18398 15262 18450
rect 15262 18398 15314 18450
rect 15314 18398 15316 18450
rect 15260 18396 15316 18398
rect 15820 18450 15876 18452
rect 15820 18398 15822 18450
rect 15822 18398 15874 18450
rect 15874 18398 15876 18450
rect 15820 18396 15876 18398
rect 16156 18562 16212 18564
rect 16156 18510 16158 18562
rect 16158 18510 16210 18562
rect 16210 18510 16212 18562
rect 16156 18508 16212 18510
rect 16044 18396 16100 18452
rect 15932 17724 15988 17780
rect 16940 20860 16996 20916
rect 17052 19516 17108 19572
rect 16828 19180 16884 19236
rect 17388 22316 17444 22372
rect 17948 22204 18004 22260
rect 17340 21978 17396 21980
rect 17340 21926 17342 21978
rect 17342 21926 17394 21978
rect 17394 21926 17396 21978
rect 17340 21924 17396 21926
rect 17444 21978 17500 21980
rect 17444 21926 17446 21978
rect 17446 21926 17498 21978
rect 17498 21926 17500 21978
rect 17444 21924 17500 21926
rect 17548 21978 17604 21980
rect 17548 21926 17550 21978
rect 17550 21926 17602 21978
rect 17602 21926 17604 21978
rect 17548 21924 17604 21926
rect 17388 21308 17444 21364
rect 18284 21868 18340 21924
rect 18732 23266 18788 23268
rect 18732 23214 18734 23266
rect 18734 23214 18786 23266
rect 18786 23214 18788 23266
rect 18732 23212 18788 23214
rect 19068 24556 19124 24612
rect 19516 25116 19572 25172
rect 19964 26514 20020 26516
rect 19964 26462 19966 26514
rect 19966 26462 20018 26514
rect 20018 26462 20020 26514
rect 19964 26460 20020 26462
rect 20412 26178 20468 26180
rect 20412 26126 20414 26178
rect 20414 26126 20466 26178
rect 20466 26126 20468 26178
rect 20412 26124 20468 26126
rect 20524 25788 20580 25844
rect 20524 25564 20580 25620
rect 20748 26290 20804 26292
rect 20748 26238 20750 26290
rect 20750 26238 20802 26290
rect 20802 26238 20804 26290
rect 20748 26236 20804 26238
rect 20300 25452 20356 25508
rect 20188 25004 20244 25060
rect 19628 24892 19684 24948
rect 19292 24722 19348 24724
rect 19292 24670 19294 24722
rect 19294 24670 19346 24722
rect 19346 24670 19348 24722
rect 19292 24668 19348 24670
rect 19516 24780 19572 24836
rect 19404 24108 19460 24164
rect 18956 23324 19012 23380
rect 19180 23996 19236 24052
rect 19292 23884 19348 23940
rect 19292 23100 19348 23156
rect 19852 24892 19908 24948
rect 19740 24668 19796 24724
rect 19852 24108 19908 24164
rect 18396 21756 18452 21812
rect 18508 22764 18564 22820
rect 18396 21474 18452 21476
rect 18396 21422 18398 21474
rect 18398 21422 18450 21474
rect 18450 21422 18452 21474
rect 18396 21420 18452 21422
rect 17836 20802 17892 20804
rect 17836 20750 17838 20802
rect 17838 20750 17890 20802
rect 17890 20750 17892 20802
rect 17836 20748 17892 20750
rect 17612 20524 17668 20580
rect 17340 20410 17396 20412
rect 17340 20358 17342 20410
rect 17342 20358 17394 20410
rect 17394 20358 17396 20410
rect 17340 20356 17396 20358
rect 17444 20410 17500 20412
rect 17444 20358 17446 20410
rect 17446 20358 17498 20410
rect 17498 20358 17500 20410
rect 17444 20356 17500 20358
rect 17548 20410 17604 20412
rect 17548 20358 17550 20410
rect 17550 20358 17602 20410
rect 17602 20358 17604 20410
rect 17548 20356 17604 20358
rect 17500 20188 17556 20244
rect 18284 20524 18340 20580
rect 17724 19122 17780 19124
rect 17724 19070 17726 19122
rect 17726 19070 17778 19122
rect 17778 19070 17780 19122
rect 17724 19068 17780 19070
rect 17500 18956 17556 19012
rect 18284 19010 18340 19012
rect 18284 18958 18286 19010
rect 18286 18958 18338 19010
rect 18338 18958 18340 19010
rect 18284 18956 18340 18958
rect 17340 18842 17396 18844
rect 17340 18790 17342 18842
rect 17342 18790 17394 18842
rect 17394 18790 17396 18842
rect 17340 18788 17396 18790
rect 17444 18842 17500 18844
rect 17444 18790 17446 18842
rect 17446 18790 17498 18842
rect 17498 18790 17500 18842
rect 17444 18788 17500 18790
rect 17548 18842 17604 18844
rect 17548 18790 17550 18842
rect 17550 18790 17602 18842
rect 17602 18790 17604 18842
rect 18396 18844 18452 18900
rect 17548 18788 17604 18790
rect 17052 18620 17108 18676
rect 17612 17836 17668 17892
rect 18844 22370 18900 22372
rect 18844 22318 18846 22370
rect 18846 22318 18898 22370
rect 18898 22318 18900 22370
rect 18844 22316 18900 22318
rect 19068 22764 19124 22820
rect 19180 22540 19236 22596
rect 19852 23436 19908 23492
rect 20636 25394 20692 25396
rect 20636 25342 20638 25394
rect 20638 25342 20690 25394
rect 20690 25342 20692 25394
rect 20636 25340 20692 25342
rect 20636 25116 20692 25172
rect 20300 24780 20356 24836
rect 20412 24722 20468 24724
rect 20412 24670 20414 24722
rect 20414 24670 20466 24722
rect 20466 24670 20468 24722
rect 20412 24668 20468 24670
rect 20300 24610 20356 24612
rect 20300 24558 20302 24610
rect 20302 24558 20354 24610
rect 20354 24558 20356 24610
rect 20300 24556 20356 24558
rect 20188 24444 20244 24500
rect 20076 23938 20132 23940
rect 20076 23886 20078 23938
rect 20078 23886 20130 23938
rect 20130 23886 20132 23938
rect 20076 23884 20132 23886
rect 20076 23714 20132 23716
rect 20076 23662 20078 23714
rect 20078 23662 20130 23714
rect 20130 23662 20132 23714
rect 20076 23660 20132 23662
rect 19964 23548 20020 23604
rect 20636 23772 20692 23828
rect 20412 23378 20468 23380
rect 20412 23326 20414 23378
rect 20414 23326 20466 23378
rect 20466 23326 20468 23378
rect 20412 23324 20468 23326
rect 20188 23100 20244 23156
rect 19852 22930 19908 22932
rect 19852 22878 19854 22930
rect 19854 22878 19906 22930
rect 19906 22878 19908 22930
rect 19852 22876 19908 22878
rect 20188 22764 20244 22820
rect 19740 22540 19796 22596
rect 19068 21644 19124 21700
rect 19180 21756 19236 21812
rect 18732 21586 18788 21588
rect 18732 21534 18734 21586
rect 18734 21534 18786 21586
rect 18786 21534 18788 21586
rect 18732 21532 18788 21534
rect 19404 21644 19460 21700
rect 18844 20690 18900 20692
rect 18844 20638 18846 20690
rect 18846 20638 18898 20690
rect 18898 20638 18900 20690
rect 18844 20636 18900 20638
rect 19852 22428 19908 22484
rect 19628 20578 19684 20580
rect 19628 20526 19630 20578
rect 19630 20526 19682 20578
rect 19682 20526 19684 20578
rect 19628 20524 19684 20526
rect 20636 23324 20692 23380
rect 21084 26684 21140 26740
rect 20972 26572 21028 26628
rect 20972 23772 21028 23828
rect 21644 26684 21700 26740
rect 21372 25898 21428 25900
rect 21372 25846 21374 25898
rect 21374 25846 21426 25898
rect 21426 25846 21428 25898
rect 21372 25844 21428 25846
rect 21476 25898 21532 25900
rect 21476 25846 21478 25898
rect 21478 25846 21530 25898
rect 21530 25846 21532 25898
rect 21476 25844 21532 25846
rect 21580 25898 21636 25900
rect 21580 25846 21582 25898
rect 21582 25846 21634 25898
rect 21634 25846 21636 25898
rect 21580 25844 21636 25846
rect 21196 25228 21252 25284
rect 22316 29708 22372 29764
rect 22652 29372 22708 29428
rect 22204 27244 22260 27300
rect 22316 28364 22372 28420
rect 22876 29426 22932 29428
rect 22876 29374 22878 29426
rect 22878 29374 22930 29426
rect 22930 29374 22932 29426
rect 22876 29372 22932 29374
rect 22988 29260 23044 29316
rect 23436 29148 23492 29204
rect 22428 27132 22484 27188
rect 23436 27132 23492 27188
rect 22092 26460 22148 26516
rect 23100 26348 23156 26404
rect 21868 26124 21924 26180
rect 22204 26124 22260 26180
rect 22316 26012 22372 26068
rect 22092 25676 22148 25732
rect 21980 25228 22036 25284
rect 21196 24444 21252 24500
rect 21372 24330 21428 24332
rect 21196 24220 21252 24276
rect 21372 24278 21374 24330
rect 21374 24278 21426 24330
rect 21426 24278 21428 24330
rect 21372 24276 21428 24278
rect 21476 24330 21532 24332
rect 21476 24278 21478 24330
rect 21478 24278 21530 24330
rect 21530 24278 21532 24330
rect 21476 24276 21532 24278
rect 21580 24330 21636 24332
rect 21580 24278 21582 24330
rect 21582 24278 21634 24330
rect 21634 24278 21636 24330
rect 21580 24276 21636 24278
rect 20860 23436 20916 23492
rect 20860 22988 20916 23044
rect 20748 22594 20804 22596
rect 20748 22542 20750 22594
rect 20750 22542 20802 22594
rect 20802 22542 20804 22594
rect 20748 22540 20804 22542
rect 20636 22428 20692 22484
rect 20524 22316 20580 22372
rect 20636 22258 20692 22260
rect 20636 22206 20638 22258
rect 20638 22206 20690 22258
rect 20690 22206 20692 22258
rect 20636 22204 20692 22206
rect 19964 21868 20020 21924
rect 20524 21420 20580 21476
rect 18732 20188 18788 20244
rect 19404 19852 19460 19908
rect 19068 19346 19124 19348
rect 19068 19294 19070 19346
rect 19070 19294 19122 19346
rect 19122 19294 19124 19346
rect 19068 19292 19124 19294
rect 18620 18674 18676 18676
rect 18620 18622 18622 18674
rect 18622 18622 18674 18674
rect 18674 18622 18676 18674
rect 18620 18620 18676 18622
rect 19404 18620 19460 18676
rect 19068 18508 19124 18564
rect 18620 17836 18676 17892
rect 16716 17500 16772 17556
rect 17340 17274 17396 17276
rect 17340 17222 17342 17274
rect 17342 17222 17394 17274
rect 17394 17222 17396 17274
rect 17340 17220 17396 17222
rect 17444 17274 17500 17276
rect 17444 17222 17446 17274
rect 17446 17222 17498 17274
rect 17498 17222 17500 17274
rect 17444 17220 17500 17222
rect 17548 17274 17604 17276
rect 17548 17222 17550 17274
rect 17550 17222 17602 17274
rect 17602 17222 17604 17274
rect 17548 17220 17604 17222
rect 16828 16882 16884 16884
rect 16828 16830 16830 16882
rect 16830 16830 16882 16882
rect 16882 16830 16884 16882
rect 16828 16828 16884 16830
rect 15036 16268 15092 16324
rect 14028 15372 14084 15428
rect 14700 15372 14756 15428
rect 11564 14252 11620 14308
rect 12012 13916 12068 13972
rect 11676 13468 11732 13524
rect 12236 14306 12292 14308
rect 12236 14254 12238 14306
rect 12238 14254 12290 14306
rect 12290 14254 12292 14306
rect 12236 14252 12292 14254
rect 11452 12348 11508 12404
rect 10892 11676 10948 11732
rect 9884 11170 9940 11172
rect 9884 11118 9886 11170
rect 9886 11118 9938 11170
rect 9938 11118 9940 11170
rect 9884 11116 9940 11118
rect 9276 11002 9332 11004
rect 9276 10950 9278 11002
rect 9278 10950 9330 11002
rect 9330 10950 9332 11002
rect 9276 10948 9332 10950
rect 9380 11002 9436 11004
rect 9380 10950 9382 11002
rect 9382 10950 9434 11002
rect 9434 10950 9436 11002
rect 9380 10948 9436 10950
rect 9484 11002 9540 11004
rect 9484 10950 9486 11002
rect 9486 10950 9538 11002
rect 9538 10950 9540 11002
rect 9484 10948 9540 10950
rect 9660 10722 9716 10724
rect 9660 10670 9662 10722
rect 9662 10670 9714 10722
rect 9714 10670 9716 10722
rect 9660 10668 9716 10670
rect 8764 9772 8820 9828
rect 8652 9714 8708 9716
rect 8652 9662 8654 9714
rect 8654 9662 8706 9714
rect 8706 9662 8708 9714
rect 8652 9660 8708 9662
rect 8316 7420 8372 7476
rect 7420 6972 7476 7028
rect 9100 9548 9156 9604
rect 7420 6748 7476 6804
rect 8428 7196 8484 7252
rect 8092 6188 8148 6244
rect 6860 5068 6916 5124
rect 6524 4956 6580 5012
rect 8764 6748 8820 6804
rect 7868 4284 7924 4340
rect 8428 4338 8484 4340
rect 8428 4286 8430 4338
rect 8430 4286 8482 4338
rect 8482 4286 8484 4338
rect 8428 4284 8484 4286
rect 10892 11170 10948 11172
rect 10892 11118 10894 11170
rect 10894 11118 10946 11170
rect 10946 11118 10948 11170
rect 10892 11116 10948 11118
rect 10668 10780 10724 10836
rect 9996 10444 10052 10500
rect 9660 9548 9716 9604
rect 9276 9434 9332 9436
rect 9276 9382 9278 9434
rect 9278 9382 9330 9434
rect 9330 9382 9332 9434
rect 9276 9380 9332 9382
rect 9380 9434 9436 9436
rect 9380 9382 9382 9434
rect 9382 9382 9434 9434
rect 9434 9382 9436 9434
rect 9380 9380 9436 9382
rect 9484 9434 9540 9436
rect 9484 9382 9486 9434
rect 9486 9382 9538 9434
rect 9538 9382 9540 9434
rect 9484 9380 9540 9382
rect 9772 8876 9828 8932
rect 9276 7866 9332 7868
rect 9276 7814 9278 7866
rect 9278 7814 9330 7866
rect 9330 7814 9332 7866
rect 9276 7812 9332 7814
rect 9380 7866 9436 7868
rect 9380 7814 9382 7866
rect 9382 7814 9434 7866
rect 9434 7814 9436 7866
rect 9380 7812 9436 7814
rect 9484 7866 9540 7868
rect 9484 7814 9486 7866
rect 9486 7814 9538 7866
rect 9538 7814 9540 7866
rect 9484 7812 9540 7814
rect 9100 6636 9156 6692
rect 9212 7644 9268 7700
rect 9436 6860 9492 6916
rect 9660 6860 9716 6916
rect 9660 6690 9716 6692
rect 9660 6638 9662 6690
rect 9662 6638 9714 6690
rect 9714 6638 9716 6690
rect 9660 6636 9716 6638
rect 9548 6524 9604 6580
rect 10444 9436 10500 9492
rect 11564 11564 11620 11620
rect 12124 12460 12180 12516
rect 12012 12236 12068 12292
rect 13308 14922 13364 14924
rect 13308 14870 13310 14922
rect 13310 14870 13362 14922
rect 13362 14870 13364 14922
rect 13308 14868 13364 14870
rect 13412 14922 13468 14924
rect 13412 14870 13414 14922
rect 13414 14870 13466 14922
rect 13466 14870 13468 14922
rect 13412 14868 13468 14870
rect 13516 14922 13572 14924
rect 13516 14870 13518 14922
rect 13518 14870 13570 14922
rect 13570 14870 13572 14922
rect 13516 14868 13572 14870
rect 14476 14588 14532 14644
rect 12460 13970 12516 13972
rect 12460 13918 12462 13970
rect 12462 13918 12514 13970
rect 12514 13918 12516 13970
rect 12460 13916 12516 13918
rect 12572 14252 12628 14308
rect 12908 13692 12964 13748
rect 13308 13354 13364 13356
rect 13308 13302 13310 13354
rect 13310 13302 13362 13354
rect 13362 13302 13364 13354
rect 13308 13300 13364 13302
rect 13412 13354 13468 13356
rect 13412 13302 13414 13354
rect 13414 13302 13466 13354
rect 13466 13302 13468 13354
rect 13412 13300 13468 13302
rect 13516 13354 13572 13356
rect 13516 13302 13518 13354
rect 13518 13302 13570 13354
rect 13570 13302 13572 13354
rect 13516 13300 13572 13302
rect 13356 13020 13412 13076
rect 12348 12236 12404 12292
rect 12236 11564 12292 11620
rect 12236 11340 12292 11396
rect 10780 10498 10836 10500
rect 10780 10446 10782 10498
rect 10782 10446 10834 10498
rect 10834 10446 10836 10498
rect 10780 10444 10836 10446
rect 10220 9154 10276 9156
rect 10220 9102 10222 9154
rect 10222 9102 10274 9154
rect 10274 9102 10276 9154
rect 10220 9100 10276 9102
rect 9996 7644 10052 7700
rect 10892 9436 10948 9492
rect 11900 9548 11956 9604
rect 11564 9100 11620 9156
rect 10892 9042 10948 9044
rect 10892 8990 10894 9042
rect 10894 8990 10946 9042
rect 10946 8990 10948 9042
rect 10892 8988 10948 8990
rect 11340 9042 11396 9044
rect 11340 8990 11342 9042
rect 11342 8990 11394 9042
rect 11394 8990 11396 9042
rect 11340 8988 11396 8990
rect 10780 8764 10836 8820
rect 11564 8428 11620 8484
rect 11788 8876 11844 8932
rect 11676 8258 11732 8260
rect 11676 8206 11678 8258
rect 11678 8206 11730 8258
rect 11730 8206 11732 8258
rect 11676 8204 11732 8206
rect 10780 7308 10836 7364
rect 9884 6412 9940 6468
rect 9276 6298 9332 6300
rect 9276 6246 9278 6298
rect 9278 6246 9330 6298
rect 9330 6246 9332 6298
rect 9276 6244 9332 6246
rect 9380 6298 9436 6300
rect 9380 6246 9382 6298
rect 9382 6246 9434 6298
rect 9434 6246 9436 6298
rect 9380 6244 9436 6246
rect 9484 6298 9540 6300
rect 9484 6246 9486 6298
rect 9486 6246 9538 6298
rect 9538 6246 9540 6298
rect 9484 6244 9540 6246
rect 9660 6300 9716 6356
rect 9772 6018 9828 6020
rect 9772 5966 9774 6018
rect 9774 5966 9826 6018
rect 9826 5966 9828 6018
rect 9772 5964 9828 5966
rect 9772 5682 9828 5684
rect 9772 5630 9774 5682
rect 9774 5630 9826 5682
rect 9826 5630 9828 5682
rect 9772 5628 9828 5630
rect 9772 5234 9828 5236
rect 9772 5182 9774 5234
rect 9774 5182 9826 5234
rect 9826 5182 9828 5234
rect 9772 5180 9828 5182
rect 9276 4730 9332 4732
rect 9276 4678 9278 4730
rect 9278 4678 9330 4730
rect 9330 4678 9332 4730
rect 9276 4676 9332 4678
rect 9380 4730 9436 4732
rect 9380 4678 9382 4730
rect 9382 4678 9434 4730
rect 9434 4678 9436 4730
rect 9380 4676 9436 4678
rect 9484 4730 9540 4732
rect 9484 4678 9486 4730
rect 9486 4678 9538 4730
rect 9538 4678 9540 4730
rect 9484 4676 9540 4678
rect 7868 3388 7924 3444
rect 10332 6578 10388 6580
rect 10332 6526 10334 6578
rect 10334 6526 10386 6578
rect 10386 6526 10388 6578
rect 10332 6524 10388 6526
rect 10220 6300 10276 6356
rect 12796 12236 12852 12292
rect 13356 12290 13412 12292
rect 13356 12238 13358 12290
rect 13358 12238 13410 12290
rect 13410 12238 13412 12290
rect 13356 12236 13412 12238
rect 14028 14364 14084 14420
rect 12572 11676 12628 11732
rect 13308 11786 13364 11788
rect 13132 11676 13188 11732
rect 13308 11734 13310 11786
rect 13310 11734 13362 11786
rect 13362 11734 13364 11786
rect 13308 11732 13364 11734
rect 13412 11786 13468 11788
rect 13412 11734 13414 11786
rect 13414 11734 13466 11786
rect 13466 11734 13468 11786
rect 13412 11732 13468 11734
rect 13516 11786 13572 11788
rect 13516 11734 13518 11786
rect 13518 11734 13570 11786
rect 13570 11734 13572 11786
rect 13516 11732 13572 11734
rect 12796 11564 12852 11620
rect 13020 9884 13076 9940
rect 13468 11394 13524 11396
rect 13468 11342 13470 11394
rect 13470 11342 13522 11394
rect 13522 11342 13524 11394
rect 13468 11340 13524 11342
rect 14476 14252 14532 14308
rect 13692 11340 13748 11396
rect 13308 10218 13364 10220
rect 13308 10166 13310 10218
rect 13310 10166 13362 10218
rect 13362 10166 13364 10218
rect 13308 10164 13364 10166
rect 13412 10218 13468 10220
rect 13412 10166 13414 10218
rect 13414 10166 13466 10218
rect 13466 10166 13468 10218
rect 13412 10164 13468 10166
rect 13516 10218 13572 10220
rect 13516 10166 13518 10218
rect 13518 10166 13570 10218
rect 13570 10166 13572 10218
rect 13516 10164 13572 10166
rect 13804 9996 13860 10052
rect 16604 15372 16660 15428
rect 16828 14924 16884 14980
rect 16380 14700 16436 14756
rect 16940 14476 16996 14532
rect 15148 14364 15204 14420
rect 16828 14306 16884 14308
rect 16828 14254 16830 14306
rect 16830 14254 16882 14306
rect 16882 14254 16884 14306
rect 16828 14252 16884 14254
rect 17612 15986 17668 15988
rect 17612 15934 17614 15986
rect 17614 15934 17666 15986
rect 17666 15934 17668 15986
rect 17612 15932 17668 15934
rect 17340 15706 17396 15708
rect 17340 15654 17342 15706
rect 17342 15654 17394 15706
rect 17394 15654 17396 15706
rect 17340 15652 17396 15654
rect 17444 15706 17500 15708
rect 17444 15654 17446 15706
rect 17446 15654 17498 15706
rect 17498 15654 17500 15706
rect 17444 15652 17500 15654
rect 17548 15706 17604 15708
rect 17548 15654 17550 15706
rect 17550 15654 17602 15706
rect 17602 15654 17604 15706
rect 17548 15652 17604 15654
rect 17164 15260 17220 15316
rect 18732 17612 18788 17668
rect 17948 17164 18004 17220
rect 17948 16828 18004 16884
rect 17836 16044 17892 16100
rect 18172 16604 18228 16660
rect 18620 17442 18676 17444
rect 18620 17390 18622 17442
rect 18622 17390 18674 17442
rect 18674 17390 18676 17442
rect 18620 17388 18676 17390
rect 18844 16716 18900 16772
rect 17836 15538 17892 15540
rect 17836 15486 17838 15538
rect 17838 15486 17890 15538
rect 17890 15486 17892 15538
rect 17836 15484 17892 15486
rect 18172 15874 18228 15876
rect 18172 15822 18174 15874
rect 18174 15822 18226 15874
rect 18226 15822 18228 15874
rect 18172 15820 18228 15822
rect 18060 15484 18116 15540
rect 17948 15372 18004 15428
rect 18732 16604 18788 16660
rect 18620 15820 18676 15876
rect 18508 15538 18564 15540
rect 18508 15486 18510 15538
rect 18510 15486 18562 15538
rect 18562 15486 18564 15538
rect 18508 15484 18564 15486
rect 17164 14754 17220 14756
rect 17164 14702 17166 14754
rect 17166 14702 17218 14754
rect 17218 14702 17220 14754
rect 17164 14700 17220 14702
rect 17836 14924 17892 14980
rect 18284 15314 18340 15316
rect 18284 15262 18286 15314
rect 18286 15262 18338 15314
rect 18338 15262 18340 15314
rect 18284 15260 18340 15262
rect 18508 15260 18564 15316
rect 20076 20076 20132 20132
rect 19964 18562 20020 18564
rect 19964 18510 19966 18562
rect 19966 18510 20018 18562
rect 20018 18510 20020 18562
rect 19964 18508 20020 18510
rect 19852 18450 19908 18452
rect 19852 18398 19854 18450
rect 19854 18398 19906 18450
rect 19906 18398 19908 18450
rect 19852 18396 19908 18398
rect 19964 17948 20020 18004
rect 19404 17442 19460 17444
rect 19404 17390 19406 17442
rect 19406 17390 19458 17442
rect 19458 17390 19460 17442
rect 19404 17388 19460 17390
rect 19404 16492 19460 16548
rect 19068 16098 19124 16100
rect 19068 16046 19070 16098
rect 19070 16046 19122 16098
rect 19122 16046 19124 16098
rect 19068 16044 19124 16046
rect 18844 15708 18900 15764
rect 19292 15820 19348 15876
rect 18844 15484 18900 15540
rect 18732 15426 18788 15428
rect 18732 15374 18734 15426
rect 18734 15374 18786 15426
rect 18786 15374 18788 15426
rect 18732 15372 18788 15374
rect 18172 14924 18228 14980
rect 17340 14138 17396 14140
rect 17340 14086 17342 14138
rect 17342 14086 17394 14138
rect 17394 14086 17396 14138
rect 17340 14084 17396 14086
rect 17444 14138 17500 14140
rect 17444 14086 17446 14138
rect 17446 14086 17498 14138
rect 17498 14086 17500 14138
rect 17444 14084 17500 14086
rect 17548 14138 17604 14140
rect 17548 14086 17550 14138
rect 17550 14086 17602 14138
rect 17602 14086 17604 14138
rect 17836 14140 17892 14196
rect 17548 14084 17604 14086
rect 17052 13916 17108 13972
rect 14812 13746 14868 13748
rect 14812 13694 14814 13746
rect 14814 13694 14866 13746
rect 14866 13694 14868 13746
rect 14812 13692 14868 13694
rect 15932 13634 15988 13636
rect 15932 13582 15934 13634
rect 15934 13582 15986 13634
rect 15986 13582 15988 13634
rect 15932 13580 15988 13582
rect 16380 13580 16436 13636
rect 14924 13468 14980 13524
rect 15596 13522 15652 13524
rect 15596 13470 15598 13522
rect 15598 13470 15650 13522
rect 15650 13470 15652 13522
rect 15596 13468 15652 13470
rect 16716 13804 16772 13860
rect 17612 13746 17668 13748
rect 17612 13694 17614 13746
rect 17614 13694 17666 13746
rect 17666 13694 17668 13746
rect 17612 13692 17668 13694
rect 17724 13468 17780 13524
rect 16604 12908 16660 12964
rect 17164 12962 17220 12964
rect 17164 12910 17166 12962
rect 17166 12910 17218 12962
rect 17218 12910 17220 12962
rect 17164 12908 17220 12910
rect 17340 12570 17396 12572
rect 17340 12518 17342 12570
rect 17342 12518 17394 12570
rect 17394 12518 17396 12570
rect 17340 12516 17396 12518
rect 17444 12570 17500 12572
rect 17444 12518 17446 12570
rect 17446 12518 17498 12570
rect 17498 12518 17500 12570
rect 17444 12516 17500 12518
rect 17548 12570 17604 12572
rect 17548 12518 17550 12570
rect 17550 12518 17602 12570
rect 17602 12518 17604 12570
rect 17548 12516 17604 12518
rect 16716 11900 16772 11956
rect 16716 11452 16772 11508
rect 18508 14642 18564 14644
rect 18508 14590 18510 14642
rect 18510 14590 18562 14642
rect 18562 14590 18564 14642
rect 18508 14588 18564 14590
rect 18620 14530 18676 14532
rect 18620 14478 18622 14530
rect 18622 14478 18674 14530
rect 18674 14478 18676 14530
rect 18620 14476 18676 14478
rect 18732 14252 18788 14308
rect 18508 13970 18564 13972
rect 18508 13918 18510 13970
rect 18510 13918 18562 13970
rect 18562 13918 18564 13970
rect 18508 13916 18564 13918
rect 19292 15538 19348 15540
rect 19292 15486 19294 15538
rect 19294 15486 19346 15538
rect 19346 15486 19348 15538
rect 19292 15484 19348 15486
rect 19404 15148 19460 15204
rect 19852 17388 19908 17444
rect 19628 17164 19684 17220
rect 20300 19346 20356 19348
rect 20300 19294 20302 19346
rect 20302 19294 20354 19346
rect 20354 19294 20356 19346
rect 20300 19292 20356 19294
rect 20972 20972 21028 21028
rect 20524 19964 20580 20020
rect 20412 19068 20468 19124
rect 19068 14476 19124 14532
rect 19292 14364 19348 14420
rect 19516 14418 19572 14420
rect 19516 14366 19518 14418
rect 19518 14366 19570 14418
rect 19570 14366 19572 14418
rect 19516 14364 19572 14366
rect 19404 14306 19460 14308
rect 19404 14254 19406 14306
rect 19406 14254 19458 14306
rect 19458 14254 19460 14306
rect 19404 14252 19460 14254
rect 19292 13970 19348 13972
rect 19292 13918 19294 13970
rect 19294 13918 19346 13970
rect 19346 13918 19348 13970
rect 19292 13916 19348 13918
rect 19180 13804 19236 13860
rect 18732 13468 18788 13524
rect 18396 13244 18452 13300
rect 20188 18396 20244 18452
rect 20748 18844 20804 18900
rect 20972 20130 21028 20132
rect 20972 20078 20974 20130
rect 20974 20078 21026 20130
rect 21026 20078 21028 20130
rect 20972 20076 21028 20078
rect 21308 23436 21364 23492
rect 21868 23660 21924 23716
rect 21980 23884 22036 23940
rect 21644 23324 21700 23380
rect 21532 23100 21588 23156
rect 21372 22762 21428 22764
rect 21372 22710 21374 22762
rect 21374 22710 21426 22762
rect 21426 22710 21428 22762
rect 21372 22708 21428 22710
rect 21476 22762 21532 22764
rect 21476 22710 21478 22762
rect 21478 22710 21530 22762
rect 21530 22710 21532 22762
rect 21476 22708 21532 22710
rect 21580 22762 21636 22764
rect 21580 22710 21582 22762
rect 21582 22710 21634 22762
rect 21634 22710 21636 22762
rect 21580 22708 21636 22710
rect 21420 22204 21476 22260
rect 21308 22146 21364 22148
rect 21308 22094 21310 22146
rect 21310 22094 21362 22146
rect 21362 22094 21364 22146
rect 21308 22092 21364 22094
rect 21644 22258 21700 22260
rect 21644 22206 21646 22258
rect 21646 22206 21698 22258
rect 21698 22206 21700 22258
rect 21644 22204 21700 22206
rect 21644 21644 21700 21700
rect 21372 21194 21428 21196
rect 21372 21142 21374 21194
rect 21374 21142 21426 21194
rect 21426 21142 21428 21194
rect 21372 21140 21428 21142
rect 21476 21194 21532 21196
rect 21476 21142 21478 21194
rect 21478 21142 21530 21194
rect 21530 21142 21532 21194
rect 21476 21140 21532 21142
rect 21580 21194 21636 21196
rect 21580 21142 21582 21194
rect 21582 21142 21634 21194
rect 21634 21142 21636 21194
rect 21580 21140 21636 21142
rect 21868 22764 21924 22820
rect 22092 23714 22148 23716
rect 22092 23662 22094 23714
rect 22094 23662 22146 23714
rect 22146 23662 22148 23714
rect 22092 23660 22148 23662
rect 21980 21532 22036 21588
rect 21868 21420 21924 21476
rect 21756 21084 21812 21140
rect 21868 21196 21924 21252
rect 21420 20188 21476 20244
rect 21756 19964 21812 20020
rect 21980 19964 22036 20020
rect 21532 19740 21588 19796
rect 21980 19740 22036 19796
rect 21372 19626 21428 19628
rect 21372 19574 21374 19626
rect 21374 19574 21426 19626
rect 21426 19574 21428 19626
rect 21372 19572 21428 19574
rect 21476 19626 21532 19628
rect 21476 19574 21478 19626
rect 21478 19574 21530 19626
rect 21530 19574 21532 19626
rect 21476 19572 21532 19574
rect 21580 19626 21636 19628
rect 21580 19574 21582 19626
rect 21582 19574 21634 19626
rect 21634 19574 21636 19626
rect 21580 19572 21636 19574
rect 21868 19404 21924 19460
rect 22652 24556 22708 24612
rect 22428 23996 22484 24052
rect 23436 26124 23492 26180
rect 23436 23938 23492 23940
rect 23436 23886 23438 23938
rect 23438 23886 23490 23938
rect 23490 23886 23492 23938
rect 23436 23884 23492 23886
rect 22876 23826 22932 23828
rect 22876 23774 22878 23826
rect 22878 23774 22930 23826
rect 22930 23774 22932 23826
rect 22876 23772 22932 23774
rect 24556 31276 24612 31332
rect 24892 31106 24948 31108
rect 24892 31054 24894 31106
rect 24894 31054 24946 31106
rect 24946 31054 24948 31106
rect 24892 31052 24948 31054
rect 24332 30156 24388 30212
rect 24332 29986 24388 29988
rect 24332 29934 24334 29986
rect 24334 29934 24386 29986
rect 24386 29934 24388 29986
rect 24332 29932 24388 29934
rect 24108 29596 24164 29652
rect 24668 29596 24724 29652
rect 23996 28812 24052 28868
rect 24556 28588 24612 28644
rect 24332 28252 24388 28308
rect 24668 28700 24724 28756
rect 24780 29260 24836 29316
rect 23996 27804 24052 27860
rect 24108 26908 24164 26964
rect 24892 29148 24948 29204
rect 25404 31386 25460 31388
rect 25404 31334 25406 31386
rect 25406 31334 25458 31386
rect 25458 31334 25460 31386
rect 25404 31332 25460 31334
rect 25508 31386 25564 31388
rect 25508 31334 25510 31386
rect 25510 31334 25562 31386
rect 25562 31334 25564 31386
rect 25508 31332 25564 31334
rect 25612 31386 25668 31388
rect 25612 31334 25614 31386
rect 25614 31334 25666 31386
rect 25666 31334 25668 31386
rect 25612 31332 25668 31334
rect 26236 31218 26292 31220
rect 26236 31166 26238 31218
rect 26238 31166 26290 31218
rect 26290 31166 26292 31218
rect 26236 31164 26292 31166
rect 25228 31052 25284 31108
rect 25228 30716 25284 30772
rect 25340 30156 25396 30212
rect 26572 30156 26628 30212
rect 25564 30098 25620 30100
rect 25564 30046 25566 30098
rect 25566 30046 25618 30098
rect 25618 30046 25620 30098
rect 25564 30044 25620 30046
rect 25404 29818 25460 29820
rect 25404 29766 25406 29818
rect 25406 29766 25458 29818
rect 25458 29766 25460 29818
rect 25404 29764 25460 29766
rect 25508 29818 25564 29820
rect 25508 29766 25510 29818
rect 25510 29766 25562 29818
rect 25562 29766 25564 29818
rect 25508 29764 25564 29766
rect 25612 29818 25668 29820
rect 25612 29766 25614 29818
rect 25614 29766 25666 29818
rect 25666 29766 25668 29818
rect 25612 29764 25668 29766
rect 25228 29148 25284 29204
rect 25564 28754 25620 28756
rect 25564 28702 25566 28754
rect 25566 28702 25618 28754
rect 25618 28702 25620 28754
rect 25564 28700 25620 28702
rect 25676 28364 25732 28420
rect 25404 28250 25460 28252
rect 25404 28198 25406 28250
rect 25406 28198 25458 28250
rect 25458 28198 25460 28250
rect 25404 28196 25460 28198
rect 25508 28250 25564 28252
rect 25508 28198 25510 28250
rect 25510 28198 25562 28250
rect 25562 28198 25564 28250
rect 25508 28196 25564 28198
rect 25612 28250 25668 28252
rect 25612 28198 25614 28250
rect 25614 28198 25666 28250
rect 25666 28198 25668 28250
rect 25788 28252 25844 28308
rect 25612 28196 25668 28198
rect 25116 27468 25172 27524
rect 25004 27356 25060 27412
rect 23996 26236 24052 26292
rect 24444 25564 24500 25620
rect 23996 25340 24052 25396
rect 22540 23154 22596 23156
rect 22540 23102 22542 23154
rect 22542 23102 22594 23154
rect 22594 23102 22596 23154
rect 22540 23100 22596 23102
rect 22988 22764 23044 22820
rect 22316 21644 22372 21700
rect 22316 21196 22372 21252
rect 22764 21756 22820 21812
rect 22764 21532 22820 21588
rect 22204 20076 22260 20132
rect 22540 21420 22596 21476
rect 20860 18508 20916 18564
rect 20748 18284 20804 18340
rect 20524 17948 20580 18004
rect 21644 18450 21700 18452
rect 21644 18398 21646 18450
rect 21646 18398 21698 18450
rect 21698 18398 21700 18450
rect 21644 18396 21700 18398
rect 22652 20860 22708 20916
rect 22652 20524 22708 20580
rect 22428 19964 22484 20020
rect 22876 21196 22932 21252
rect 22988 20972 23044 21028
rect 23884 23436 23940 23492
rect 23436 22876 23492 22932
rect 23212 22092 23268 22148
rect 22876 20130 22932 20132
rect 22876 20078 22878 20130
rect 22878 20078 22930 20130
rect 22930 20078 22932 20130
rect 22876 20076 22932 20078
rect 23100 19404 23156 19460
rect 23884 22540 23940 22596
rect 23884 22092 23940 22148
rect 23772 21810 23828 21812
rect 23772 21758 23774 21810
rect 23774 21758 23826 21810
rect 23826 21758 23828 21810
rect 23772 21756 23828 21758
rect 23660 21586 23716 21588
rect 23660 21534 23662 21586
rect 23662 21534 23714 21586
rect 23714 21534 23716 21586
rect 23660 21532 23716 21534
rect 23772 19852 23828 19908
rect 23884 20076 23940 20132
rect 21868 18732 21924 18788
rect 22316 18844 22372 18900
rect 22316 18508 22372 18564
rect 22092 18450 22148 18452
rect 22092 18398 22094 18450
rect 22094 18398 22146 18450
rect 22146 18398 22148 18450
rect 22092 18396 22148 18398
rect 21868 18172 21924 18228
rect 20636 17724 20692 17780
rect 20188 16492 20244 16548
rect 20300 17612 20356 17668
rect 19740 15874 19796 15876
rect 19740 15822 19742 15874
rect 19742 15822 19794 15874
rect 19794 15822 19796 15874
rect 19740 15820 19796 15822
rect 19964 15372 20020 15428
rect 20076 15708 20132 15764
rect 20188 15596 20244 15652
rect 21372 18058 21428 18060
rect 21372 18006 21374 18058
rect 21374 18006 21426 18058
rect 21426 18006 21428 18058
rect 21372 18004 21428 18006
rect 21476 18058 21532 18060
rect 21476 18006 21478 18058
rect 21478 18006 21530 18058
rect 21530 18006 21532 18058
rect 21476 18004 21532 18006
rect 21580 18058 21636 18060
rect 21580 18006 21582 18058
rect 21582 18006 21634 18058
rect 21634 18006 21636 18058
rect 21580 18004 21636 18006
rect 21980 17948 22036 18004
rect 21980 17778 22036 17780
rect 21980 17726 21982 17778
rect 21982 17726 22034 17778
rect 22034 17726 22036 17778
rect 21980 17724 22036 17726
rect 20524 17388 20580 17444
rect 20412 16716 20468 16772
rect 20636 16940 20692 16996
rect 21308 17612 21364 17668
rect 21084 17164 21140 17220
rect 22204 17778 22260 17780
rect 22204 17726 22206 17778
rect 22206 17726 22258 17778
rect 22258 17726 22260 17778
rect 22204 17724 22260 17726
rect 22204 17388 22260 17444
rect 21980 17276 22036 17332
rect 21644 16940 21700 16996
rect 21372 16490 21428 16492
rect 21372 16438 21374 16490
rect 21374 16438 21426 16490
rect 21426 16438 21428 16490
rect 21372 16436 21428 16438
rect 21476 16490 21532 16492
rect 21476 16438 21478 16490
rect 21478 16438 21530 16490
rect 21530 16438 21532 16490
rect 21476 16436 21532 16438
rect 21580 16490 21636 16492
rect 21580 16438 21582 16490
rect 21582 16438 21634 16490
rect 21634 16438 21636 16490
rect 21580 16436 21636 16438
rect 21532 15986 21588 15988
rect 21532 15934 21534 15986
rect 21534 15934 21586 15986
rect 21586 15934 21588 15986
rect 21532 15932 21588 15934
rect 20524 15426 20580 15428
rect 20524 15374 20526 15426
rect 20526 15374 20578 15426
rect 20578 15374 20580 15426
rect 20524 15372 20580 15374
rect 20412 15260 20468 15316
rect 19740 14700 19796 14756
rect 19068 12962 19124 12964
rect 19068 12910 19070 12962
rect 19070 12910 19122 12962
rect 19122 12910 19124 12962
rect 19068 12908 19124 12910
rect 19852 14364 19908 14420
rect 20076 14530 20132 14532
rect 20076 14478 20078 14530
rect 20078 14478 20130 14530
rect 20130 14478 20132 14530
rect 20076 14476 20132 14478
rect 20524 14530 20580 14532
rect 20524 14478 20526 14530
rect 20526 14478 20578 14530
rect 20578 14478 20580 14530
rect 20524 14476 20580 14478
rect 21196 15538 21252 15540
rect 21196 15486 21198 15538
rect 21198 15486 21250 15538
rect 21250 15486 21252 15538
rect 21196 15484 21252 15486
rect 20636 14306 20692 14308
rect 20636 14254 20638 14306
rect 20638 14254 20690 14306
rect 20690 14254 20692 14306
rect 20636 14252 20692 14254
rect 20188 13916 20244 13972
rect 20412 13916 20468 13972
rect 20524 13746 20580 13748
rect 20524 13694 20526 13746
rect 20526 13694 20578 13746
rect 20578 13694 20580 13746
rect 20524 13692 20580 13694
rect 19852 13468 19908 13524
rect 20300 13580 20356 13636
rect 20636 13580 20692 13636
rect 21644 15820 21700 15876
rect 21644 15426 21700 15428
rect 21644 15374 21646 15426
rect 21646 15374 21698 15426
rect 21698 15374 21700 15426
rect 21644 15372 21700 15374
rect 21980 15314 22036 15316
rect 21980 15262 21982 15314
rect 21982 15262 22034 15314
rect 22034 15262 22036 15314
rect 21980 15260 22036 15262
rect 21308 15036 21364 15092
rect 21980 15036 22036 15092
rect 21372 14922 21428 14924
rect 21372 14870 21374 14922
rect 21374 14870 21426 14922
rect 21426 14870 21428 14922
rect 21372 14868 21428 14870
rect 21476 14922 21532 14924
rect 21476 14870 21478 14922
rect 21478 14870 21530 14922
rect 21530 14870 21532 14922
rect 21476 14868 21532 14870
rect 21580 14922 21636 14924
rect 21580 14870 21582 14922
rect 21582 14870 21634 14922
rect 21634 14870 21636 14922
rect 21580 14868 21636 14870
rect 21196 14476 21252 14532
rect 21084 14364 21140 14420
rect 19628 13132 19684 13188
rect 17052 11394 17108 11396
rect 17052 11342 17054 11394
rect 17054 11342 17106 11394
rect 17106 11342 17108 11394
rect 17052 11340 17108 11342
rect 13916 9938 13972 9940
rect 13916 9886 13918 9938
rect 13918 9886 13970 9938
rect 13970 9886 13972 9938
rect 13916 9884 13972 9886
rect 13132 9772 13188 9828
rect 13804 9714 13860 9716
rect 13804 9662 13806 9714
rect 13806 9662 13858 9714
rect 13858 9662 13860 9714
rect 13804 9660 13860 9662
rect 12236 9100 12292 9156
rect 12012 8428 12068 8484
rect 11004 6636 11060 6692
rect 11340 6690 11396 6692
rect 11340 6638 11342 6690
rect 11342 6638 11394 6690
rect 11394 6638 11396 6690
rect 11340 6636 11396 6638
rect 11788 6578 11844 6580
rect 11788 6526 11790 6578
rect 11790 6526 11842 6578
rect 11842 6526 11844 6578
rect 11788 6524 11844 6526
rect 11900 6300 11956 6356
rect 11900 5964 11956 6020
rect 10556 5180 10612 5236
rect 11676 5068 11732 5124
rect 9276 3162 9332 3164
rect 9276 3110 9278 3162
rect 9278 3110 9330 3162
rect 9330 3110 9332 3162
rect 9276 3108 9332 3110
rect 9380 3162 9436 3164
rect 9380 3110 9382 3162
rect 9382 3110 9434 3162
rect 9434 3110 9436 3162
rect 9380 3108 9436 3110
rect 9484 3162 9540 3164
rect 9484 3110 9486 3162
rect 9486 3110 9538 3162
rect 9538 3110 9540 3162
rect 9484 3108 9540 3110
rect 12460 8876 12516 8932
rect 12572 8988 12628 9044
rect 12348 7644 12404 7700
rect 12460 8204 12516 8260
rect 12124 7308 12180 7364
rect 12124 6860 12180 6916
rect 12348 6636 12404 6692
rect 12908 8988 12964 9044
rect 13692 9100 13748 9156
rect 13308 8650 13364 8652
rect 13308 8598 13310 8650
rect 13310 8598 13362 8650
rect 13362 8598 13364 8650
rect 13308 8596 13364 8598
rect 13412 8650 13468 8652
rect 13412 8598 13414 8650
rect 13414 8598 13466 8650
rect 13466 8598 13468 8650
rect 13412 8596 13468 8598
rect 13516 8650 13572 8652
rect 13516 8598 13518 8650
rect 13518 8598 13570 8650
rect 13570 8598 13572 8650
rect 13516 8596 13572 8598
rect 12572 6748 12628 6804
rect 12572 6466 12628 6468
rect 12572 6414 12574 6466
rect 12574 6414 12626 6466
rect 12626 6414 12628 6466
rect 12572 6412 12628 6414
rect 12124 5628 12180 5684
rect 12460 5628 12516 5684
rect 12348 5122 12404 5124
rect 12348 5070 12350 5122
rect 12350 5070 12402 5122
rect 12402 5070 12404 5122
rect 12348 5068 12404 5070
rect 13356 7308 13412 7364
rect 13692 7644 13748 7700
rect 13020 6748 13076 6804
rect 12796 6578 12852 6580
rect 12796 6526 12798 6578
rect 12798 6526 12850 6578
rect 12850 6526 12852 6578
rect 12796 6524 12852 6526
rect 12796 6188 12852 6244
rect 13308 7082 13364 7084
rect 13308 7030 13310 7082
rect 13310 7030 13362 7082
rect 13362 7030 13364 7082
rect 13308 7028 13364 7030
rect 13412 7082 13468 7084
rect 13412 7030 13414 7082
rect 13414 7030 13466 7082
rect 13466 7030 13468 7082
rect 13412 7028 13468 7030
rect 13516 7082 13572 7084
rect 13516 7030 13518 7082
rect 13518 7030 13570 7082
rect 13570 7030 13572 7082
rect 13516 7028 13572 7030
rect 13244 6076 13300 6132
rect 13580 6690 13636 6692
rect 13580 6638 13582 6690
rect 13582 6638 13634 6690
rect 13634 6638 13636 6690
rect 13580 6636 13636 6638
rect 13132 5964 13188 6020
rect 14140 10556 14196 10612
rect 17340 11002 17396 11004
rect 17340 10950 17342 11002
rect 17342 10950 17394 11002
rect 17394 10950 17396 11002
rect 17340 10948 17396 10950
rect 17444 11002 17500 11004
rect 17444 10950 17446 11002
rect 17446 10950 17498 11002
rect 17498 10950 17500 11002
rect 17444 10948 17500 10950
rect 17548 11002 17604 11004
rect 17548 10950 17550 11002
rect 17550 10950 17602 11002
rect 17602 10950 17604 11002
rect 17548 10948 17604 10950
rect 14252 10444 14308 10500
rect 14364 10108 14420 10164
rect 14028 6524 14084 6580
rect 13580 5628 13636 5684
rect 13692 6300 13748 6356
rect 13308 5514 13364 5516
rect 13308 5462 13310 5514
rect 13310 5462 13362 5514
rect 13362 5462 13364 5514
rect 13308 5460 13364 5462
rect 13412 5514 13468 5516
rect 13412 5462 13414 5514
rect 13414 5462 13466 5514
rect 13466 5462 13468 5514
rect 13412 5460 13468 5462
rect 13516 5514 13572 5516
rect 13516 5462 13518 5514
rect 13518 5462 13570 5514
rect 13570 5462 13572 5514
rect 13516 5460 13572 5462
rect 14140 6412 14196 6468
rect 14252 6188 14308 6244
rect 14364 5852 14420 5908
rect 14812 9602 14868 9604
rect 14812 9550 14814 9602
rect 14814 9550 14866 9602
rect 14866 9550 14868 9602
rect 14812 9548 14868 9550
rect 15148 10108 15204 10164
rect 15708 10610 15764 10612
rect 15708 10558 15710 10610
rect 15710 10558 15762 10610
rect 15762 10558 15764 10610
rect 15708 10556 15764 10558
rect 15932 10498 15988 10500
rect 15932 10446 15934 10498
rect 15934 10446 15986 10498
rect 15986 10446 15988 10498
rect 15932 10444 15988 10446
rect 14924 8258 14980 8260
rect 14924 8206 14926 8258
rect 14926 8206 14978 8258
rect 14978 8206 14980 8258
rect 14924 8204 14980 8206
rect 14588 5068 14644 5124
rect 14812 5180 14868 5236
rect 13308 3946 13364 3948
rect 13308 3894 13310 3946
rect 13310 3894 13362 3946
rect 13362 3894 13364 3946
rect 13308 3892 13364 3894
rect 13412 3946 13468 3948
rect 13412 3894 13414 3946
rect 13414 3894 13466 3946
rect 13466 3894 13468 3946
rect 13412 3892 13468 3894
rect 13516 3946 13572 3948
rect 13516 3894 13518 3946
rect 13518 3894 13570 3946
rect 13570 3894 13572 3946
rect 13516 3892 13572 3894
rect 12684 3388 12740 3444
rect 13356 3442 13412 3444
rect 13356 3390 13358 3442
rect 13358 3390 13410 3442
rect 13410 3390 13412 3442
rect 13356 3388 13412 3390
rect 13804 3388 13860 3444
rect 15596 9602 15652 9604
rect 15596 9550 15598 9602
rect 15598 9550 15650 9602
rect 15650 9550 15652 9602
rect 15596 9548 15652 9550
rect 16268 9212 16324 9268
rect 16156 9100 16212 9156
rect 16716 8988 16772 9044
rect 15820 8876 15876 8932
rect 16604 8930 16660 8932
rect 16604 8878 16606 8930
rect 16606 8878 16658 8930
rect 16658 8878 16660 8930
rect 16604 8876 16660 8878
rect 16716 8428 16772 8484
rect 16828 9100 16884 9156
rect 16604 7644 16660 7700
rect 16492 7532 16548 7588
rect 16716 7586 16772 7588
rect 16716 7534 16718 7586
rect 16718 7534 16770 7586
rect 16770 7534 16772 7586
rect 16716 7532 16772 7534
rect 15036 6636 15092 6692
rect 17612 10610 17668 10612
rect 17612 10558 17614 10610
rect 17614 10558 17666 10610
rect 17666 10558 17668 10610
rect 17612 10556 17668 10558
rect 17340 9434 17396 9436
rect 17340 9382 17342 9434
rect 17342 9382 17394 9434
rect 17394 9382 17396 9434
rect 17340 9380 17396 9382
rect 17444 9434 17500 9436
rect 17444 9382 17446 9434
rect 17446 9382 17498 9434
rect 17498 9382 17500 9434
rect 17444 9380 17500 9382
rect 17548 9434 17604 9436
rect 17548 9382 17550 9434
rect 17550 9382 17602 9434
rect 17602 9382 17604 9434
rect 17548 9380 17604 9382
rect 17500 9266 17556 9268
rect 17500 9214 17502 9266
rect 17502 9214 17554 9266
rect 17554 9214 17556 9266
rect 17500 9212 17556 9214
rect 17948 9772 18004 9828
rect 17948 9548 18004 9604
rect 18172 9660 18228 9716
rect 19068 9212 19124 9268
rect 17724 9042 17780 9044
rect 17724 8990 17726 9042
rect 17726 8990 17778 9042
rect 17778 8990 17780 9042
rect 17724 8988 17780 8990
rect 17836 8428 17892 8484
rect 17340 7866 17396 7868
rect 17340 7814 17342 7866
rect 17342 7814 17394 7866
rect 17394 7814 17396 7866
rect 17340 7812 17396 7814
rect 17444 7866 17500 7868
rect 17444 7814 17446 7866
rect 17446 7814 17498 7866
rect 17498 7814 17500 7866
rect 17444 7812 17500 7814
rect 17548 7866 17604 7868
rect 17548 7814 17550 7866
rect 17550 7814 17602 7866
rect 17602 7814 17604 7866
rect 17548 7812 17604 7814
rect 17612 7698 17668 7700
rect 17612 7646 17614 7698
rect 17614 7646 17666 7698
rect 17666 7646 17668 7698
rect 17612 7644 17668 7646
rect 17388 7474 17444 7476
rect 17388 7422 17390 7474
rect 17390 7422 17442 7474
rect 17442 7422 17444 7474
rect 17388 7420 17444 7422
rect 16940 7196 16996 7252
rect 17052 6690 17108 6692
rect 17052 6638 17054 6690
rect 17054 6638 17106 6690
rect 17106 6638 17108 6690
rect 17052 6636 17108 6638
rect 16604 6524 16660 6580
rect 15820 5628 15876 5684
rect 15148 5180 15204 5236
rect 17612 7196 17668 7252
rect 17276 6466 17332 6468
rect 17276 6414 17278 6466
rect 17278 6414 17330 6466
rect 17330 6414 17332 6466
rect 17276 6412 17332 6414
rect 17340 6298 17396 6300
rect 17340 6246 17342 6298
rect 17342 6246 17394 6298
rect 17394 6246 17396 6298
rect 17340 6244 17396 6246
rect 17444 6298 17500 6300
rect 17444 6246 17446 6298
rect 17446 6246 17498 6298
rect 17498 6246 17500 6298
rect 17444 6244 17500 6246
rect 17548 6298 17604 6300
rect 17548 6246 17550 6298
rect 17550 6246 17602 6298
rect 17602 6246 17604 6298
rect 17548 6244 17604 6246
rect 17276 5964 17332 6020
rect 18060 8428 18116 8484
rect 18396 7756 18452 7812
rect 18508 7420 18564 7476
rect 18620 6412 18676 6468
rect 17500 5906 17556 5908
rect 17500 5854 17502 5906
rect 17502 5854 17554 5906
rect 17554 5854 17556 5906
rect 17500 5852 17556 5854
rect 16604 5628 16660 5684
rect 16940 5740 16996 5796
rect 15372 5122 15428 5124
rect 15372 5070 15374 5122
rect 15374 5070 15426 5122
rect 15426 5070 15428 5122
rect 15372 5068 15428 5070
rect 16380 5516 16436 5572
rect 16380 5180 16436 5236
rect 15596 4338 15652 4340
rect 15596 4286 15598 4338
rect 15598 4286 15650 4338
rect 15650 4286 15652 4338
rect 15596 4284 15652 4286
rect 17724 5628 17780 5684
rect 17164 4844 17220 4900
rect 17340 4730 17396 4732
rect 17340 4678 17342 4730
rect 17342 4678 17394 4730
rect 17394 4678 17396 4730
rect 17340 4676 17396 4678
rect 17444 4730 17500 4732
rect 17444 4678 17446 4730
rect 17446 4678 17498 4730
rect 17498 4678 17500 4730
rect 17444 4676 17500 4678
rect 17548 4730 17604 4732
rect 17548 4678 17550 4730
rect 17550 4678 17602 4730
rect 17602 4678 17604 4730
rect 17548 4676 17604 4678
rect 17948 5516 18004 5572
rect 18396 5628 18452 5684
rect 18844 5404 18900 5460
rect 18396 5068 18452 5124
rect 20076 13132 20132 13188
rect 19964 12012 20020 12068
rect 19740 10834 19796 10836
rect 19740 10782 19742 10834
rect 19742 10782 19794 10834
rect 19794 10782 19796 10834
rect 19740 10780 19796 10782
rect 19292 9772 19348 9828
rect 19180 8204 19236 8260
rect 20300 10610 20356 10612
rect 20300 10558 20302 10610
rect 20302 10558 20354 10610
rect 20354 10558 20356 10610
rect 20300 10556 20356 10558
rect 20860 13356 20916 13412
rect 21084 13244 21140 13300
rect 21308 14364 21364 14420
rect 21420 14306 21476 14308
rect 21420 14254 21422 14306
rect 21422 14254 21474 14306
rect 21474 14254 21476 14306
rect 21420 14252 21476 14254
rect 21868 14028 21924 14084
rect 21644 13692 21700 13748
rect 21756 13804 21812 13860
rect 21308 13580 21364 13636
rect 21372 13354 21428 13356
rect 21372 13302 21374 13354
rect 21374 13302 21426 13354
rect 21426 13302 21428 13354
rect 21372 13300 21428 13302
rect 21476 13354 21532 13356
rect 21476 13302 21478 13354
rect 21478 13302 21530 13354
rect 21530 13302 21532 13354
rect 21476 13300 21532 13302
rect 21580 13354 21636 13356
rect 21580 13302 21582 13354
rect 21582 13302 21634 13354
rect 21634 13302 21636 13354
rect 21580 13300 21636 13302
rect 22988 19234 23044 19236
rect 22988 19182 22990 19234
rect 22990 19182 23042 19234
rect 23042 19182 23044 19234
rect 22988 19180 23044 19182
rect 22764 18562 22820 18564
rect 22764 18510 22766 18562
rect 22766 18510 22818 18562
rect 22818 18510 22820 18562
rect 22764 18508 22820 18510
rect 22988 18732 23044 18788
rect 23548 19068 23604 19124
rect 24220 23826 24276 23828
rect 24220 23774 24222 23826
rect 24222 23774 24274 23826
rect 24274 23774 24276 23826
rect 24220 23772 24276 23774
rect 24668 25340 24724 25396
rect 24444 22316 24500 22372
rect 24220 21698 24276 21700
rect 24220 21646 24222 21698
rect 24222 21646 24274 21698
rect 24274 21646 24276 21698
rect 24220 21644 24276 21646
rect 24444 21698 24500 21700
rect 24444 21646 24446 21698
rect 24446 21646 24498 21698
rect 24498 21646 24500 21698
rect 24444 21644 24500 21646
rect 24108 19628 24164 19684
rect 24108 19292 24164 19348
rect 24220 19964 24276 20020
rect 24332 19458 24388 19460
rect 24332 19406 24334 19458
rect 24334 19406 24386 19458
rect 24386 19406 24388 19458
rect 24332 19404 24388 19406
rect 22540 17554 22596 17556
rect 22540 17502 22542 17554
rect 22542 17502 22594 17554
rect 22594 17502 22596 17554
rect 22540 17500 22596 17502
rect 22652 16098 22708 16100
rect 22652 16046 22654 16098
rect 22654 16046 22706 16098
rect 22706 16046 22708 16098
rect 22652 16044 22708 16046
rect 22540 15986 22596 15988
rect 22540 15934 22542 15986
rect 22542 15934 22594 15986
rect 22594 15934 22596 15986
rect 22540 15932 22596 15934
rect 22428 15202 22484 15204
rect 22428 15150 22430 15202
rect 22430 15150 22482 15202
rect 22482 15150 22484 15202
rect 22428 15148 22484 15150
rect 22204 15036 22260 15092
rect 22204 14028 22260 14084
rect 22092 13916 22148 13972
rect 22092 13580 22148 13636
rect 22428 13186 22484 13188
rect 22428 13134 22430 13186
rect 22430 13134 22482 13186
rect 22482 13134 22484 13186
rect 22428 13132 22484 13134
rect 21868 11900 21924 11956
rect 21372 11786 21428 11788
rect 21372 11734 21374 11786
rect 21374 11734 21426 11786
rect 21426 11734 21428 11786
rect 21372 11732 21428 11734
rect 21476 11786 21532 11788
rect 21476 11734 21478 11786
rect 21478 11734 21530 11786
rect 21530 11734 21532 11786
rect 21476 11732 21532 11734
rect 21580 11786 21636 11788
rect 21580 11734 21582 11786
rect 21582 11734 21634 11786
rect 21634 11734 21636 11786
rect 21580 11732 21636 11734
rect 21532 11394 21588 11396
rect 21532 11342 21534 11394
rect 21534 11342 21586 11394
rect 21586 11342 21588 11394
rect 21532 11340 21588 11342
rect 21308 10834 21364 10836
rect 21308 10782 21310 10834
rect 21310 10782 21362 10834
rect 21362 10782 21364 10834
rect 21308 10780 21364 10782
rect 20972 10556 21028 10612
rect 20636 9996 20692 10052
rect 19628 8988 19684 9044
rect 19740 8204 19796 8260
rect 19964 9826 20020 9828
rect 19964 9774 19966 9826
rect 19966 9774 20018 9826
rect 20018 9774 20020 9826
rect 19964 9772 20020 9774
rect 20300 9772 20356 9828
rect 20636 9548 20692 9604
rect 21372 10218 21428 10220
rect 21372 10166 21374 10218
rect 21374 10166 21426 10218
rect 21426 10166 21428 10218
rect 21372 10164 21428 10166
rect 21476 10218 21532 10220
rect 21476 10166 21478 10218
rect 21478 10166 21530 10218
rect 21530 10166 21532 10218
rect 21476 10164 21532 10166
rect 21580 10218 21636 10220
rect 21580 10166 21582 10218
rect 21582 10166 21634 10218
rect 21634 10166 21636 10218
rect 21868 10220 21924 10276
rect 21580 10164 21636 10166
rect 21868 9772 21924 9828
rect 21372 8650 21428 8652
rect 21372 8598 21374 8650
rect 21374 8598 21426 8650
rect 21426 8598 21428 8650
rect 21372 8596 21428 8598
rect 21476 8650 21532 8652
rect 21476 8598 21478 8650
rect 21478 8598 21530 8650
rect 21530 8598 21532 8650
rect 21476 8596 21532 8598
rect 21580 8650 21636 8652
rect 21580 8598 21582 8650
rect 21582 8598 21634 8650
rect 21634 8598 21636 8650
rect 21580 8596 21636 8598
rect 19292 8092 19348 8148
rect 19516 7868 19572 7924
rect 19852 8034 19908 8036
rect 19852 7982 19854 8034
rect 19854 7982 19906 8034
rect 19906 7982 19908 8034
rect 19852 7980 19908 7982
rect 20300 8146 20356 8148
rect 20300 8094 20302 8146
rect 20302 8094 20354 8146
rect 20354 8094 20356 8146
rect 20300 8092 20356 8094
rect 19964 7868 20020 7924
rect 21868 8146 21924 8148
rect 21868 8094 21870 8146
rect 21870 8094 21922 8146
rect 21922 8094 21924 8146
rect 21868 8092 21924 8094
rect 20636 7644 20692 7700
rect 19292 7586 19348 7588
rect 19292 7534 19294 7586
rect 19294 7534 19346 7586
rect 19346 7534 19348 7586
rect 19292 7532 19348 7534
rect 20076 7532 20132 7588
rect 19180 7420 19236 7476
rect 19404 7308 19460 7364
rect 19068 5906 19124 5908
rect 19068 5854 19070 5906
rect 19070 5854 19122 5906
rect 19122 5854 19124 5906
rect 19068 5852 19124 5854
rect 19292 5740 19348 5796
rect 19292 5010 19348 5012
rect 19292 4958 19294 5010
rect 19294 4958 19346 5010
rect 19346 4958 19348 5010
rect 19292 4956 19348 4958
rect 19740 6018 19796 6020
rect 19740 5966 19742 6018
rect 19742 5966 19794 6018
rect 19794 5966 19796 6018
rect 19740 5964 19796 5966
rect 19740 5404 19796 5460
rect 18732 4844 18788 4900
rect 17388 4338 17444 4340
rect 17388 4286 17390 4338
rect 17390 4286 17442 4338
rect 17442 4286 17444 4338
rect 17388 4284 17444 4286
rect 19180 4172 19236 4228
rect 19740 4898 19796 4900
rect 19740 4846 19742 4898
rect 19742 4846 19794 4898
rect 19794 4846 19796 4898
rect 19740 4844 19796 4846
rect 19740 4060 19796 4116
rect 17340 3162 17396 3164
rect 17340 3110 17342 3162
rect 17342 3110 17394 3162
rect 17394 3110 17396 3162
rect 17340 3108 17396 3110
rect 17444 3162 17500 3164
rect 17444 3110 17446 3162
rect 17446 3110 17498 3162
rect 17498 3110 17500 3162
rect 17444 3108 17500 3110
rect 17548 3162 17604 3164
rect 17548 3110 17550 3162
rect 17550 3110 17602 3162
rect 17602 3110 17604 3162
rect 17548 3108 17604 3110
rect 19852 3612 19908 3668
rect 21644 7756 21700 7812
rect 21756 7586 21812 7588
rect 21756 7534 21758 7586
rect 21758 7534 21810 7586
rect 21810 7534 21812 7586
rect 21756 7532 21812 7534
rect 20748 6802 20804 6804
rect 20748 6750 20750 6802
rect 20750 6750 20802 6802
rect 20802 6750 20804 6802
rect 20748 6748 20804 6750
rect 20300 5068 20356 5124
rect 20748 5852 20804 5908
rect 20860 4338 20916 4340
rect 20860 4286 20862 4338
rect 20862 4286 20914 4338
rect 20914 4286 20916 4338
rect 20860 4284 20916 4286
rect 20300 4226 20356 4228
rect 20300 4174 20302 4226
rect 20302 4174 20354 4226
rect 20354 4174 20356 4226
rect 20300 4172 20356 4174
rect 20748 4060 20804 4116
rect 21372 7082 21428 7084
rect 21372 7030 21374 7082
rect 21374 7030 21426 7082
rect 21426 7030 21428 7082
rect 21372 7028 21428 7030
rect 21476 7082 21532 7084
rect 21476 7030 21478 7082
rect 21478 7030 21530 7082
rect 21530 7030 21532 7082
rect 21476 7028 21532 7030
rect 21580 7082 21636 7084
rect 21580 7030 21582 7082
rect 21582 7030 21634 7082
rect 21634 7030 21636 7082
rect 21580 7028 21636 7030
rect 22540 10498 22596 10500
rect 22540 10446 22542 10498
rect 22542 10446 22594 10498
rect 22594 10446 22596 10498
rect 22540 10444 22596 10446
rect 22316 10220 22372 10276
rect 22204 9938 22260 9940
rect 22204 9886 22206 9938
rect 22206 9886 22258 9938
rect 22258 9886 22260 9938
rect 22204 9884 22260 9886
rect 22988 17276 23044 17332
rect 23324 18732 23380 18788
rect 23772 18844 23828 18900
rect 24892 24444 24948 24500
rect 24892 21420 24948 21476
rect 24780 21362 24836 21364
rect 24780 21310 24782 21362
rect 24782 21310 24834 21362
rect 24834 21310 24836 21362
rect 24780 21308 24836 21310
rect 24668 20578 24724 20580
rect 24668 20526 24670 20578
rect 24670 20526 24722 20578
rect 24722 20526 24724 20578
rect 24668 20524 24724 20526
rect 24892 20076 24948 20132
rect 24780 19740 24836 19796
rect 25788 28082 25844 28084
rect 25788 28030 25790 28082
rect 25790 28030 25842 28082
rect 25842 28030 25844 28082
rect 25788 28028 25844 28030
rect 25452 27916 25508 27972
rect 25900 27804 25956 27860
rect 26124 28252 26180 28308
rect 25228 26908 25284 26964
rect 25404 26682 25460 26684
rect 25404 26630 25406 26682
rect 25406 26630 25458 26682
rect 25458 26630 25460 26682
rect 25404 26628 25460 26630
rect 25508 26682 25564 26684
rect 25508 26630 25510 26682
rect 25510 26630 25562 26682
rect 25562 26630 25564 26682
rect 25508 26628 25564 26630
rect 25612 26682 25668 26684
rect 25612 26630 25614 26682
rect 25614 26630 25666 26682
rect 25666 26630 25668 26682
rect 25612 26628 25668 26630
rect 25788 26684 25844 26740
rect 25340 26290 25396 26292
rect 25340 26238 25342 26290
rect 25342 26238 25394 26290
rect 25394 26238 25396 26290
rect 25340 26236 25396 26238
rect 25228 25228 25284 25284
rect 25404 25114 25460 25116
rect 25404 25062 25406 25114
rect 25406 25062 25458 25114
rect 25458 25062 25460 25114
rect 25404 25060 25460 25062
rect 25508 25114 25564 25116
rect 25508 25062 25510 25114
rect 25510 25062 25562 25114
rect 25562 25062 25564 25114
rect 25508 25060 25564 25062
rect 25612 25114 25668 25116
rect 25612 25062 25614 25114
rect 25614 25062 25666 25114
rect 25666 25062 25668 25114
rect 25612 25060 25668 25062
rect 25564 24946 25620 24948
rect 25564 24894 25566 24946
rect 25566 24894 25618 24946
rect 25618 24894 25620 24946
rect 25564 24892 25620 24894
rect 25228 23436 25284 23492
rect 25404 23546 25460 23548
rect 25404 23494 25406 23546
rect 25406 23494 25458 23546
rect 25458 23494 25460 23546
rect 25404 23492 25460 23494
rect 25508 23546 25564 23548
rect 25508 23494 25510 23546
rect 25510 23494 25562 23546
rect 25562 23494 25564 23546
rect 25508 23492 25564 23494
rect 25612 23546 25668 23548
rect 25612 23494 25614 23546
rect 25614 23494 25666 23546
rect 25666 23494 25668 23546
rect 25612 23492 25668 23494
rect 25228 23212 25284 23268
rect 25452 23100 25508 23156
rect 26348 29148 26404 29204
rect 26572 29036 26628 29092
rect 26908 28866 26964 28868
rect 26908 28814 26910 28866
rect 26910 28814 26962 28866
rect 26962 28814 26964 28866
rect 26908 28812 26964 28814
rect 26460 28476 26516 28532
rect 26348 28364 26404 28420
rect 26460 27970 26516 27972
rect 26460 27918 26462 27970
rect 26462 27918 26514 27970
rect 26514 27918 26516 27970
rect 26460 27916 26516 27918
rect 26796 28364 26852 28420
rect 26124 25452 26180 25508
rect 26572 25676 26628 25732
rect 26124 25116 26180 25172
rect 25900 23884 25956 23940
rect 25900 23548 25956 23604
rect 25452 22428 25508 22484
rect 25564 22540 25620 22596
rect 25228 22204 25284 22260
rect 25116 22146 25172 22148
rect 25116 22094 25118 22146
rect 25118 22094 25170 22146
rect 25170 22094 25172 22146
rect 25116 22092 25172 22094
rect 25564 22092 25620 22148
rect 25788 22428 25844 22484
rect 25404 21978 25460 21980
rect 25404 21926 25406 21978
rect 25406 21926 25458 21978
rect 25458 21926 25460 21978
rect 25404 21924 25460 21926
rect 25508 21978 25564 21980
rect 25508 21926 25510 21978
rect 25510 21926 25562 21978
rect 25562 21926 25564 21978
rect 25508 21924 25564 21926
rect 25612 21978 25668 21980
rect 25612 21926 25614 21978
rect 25614 21926 25666 21978
rect 25666 21926 25668 21978
rect 25612 21924 25668 21926
rect 25340 21698 25396 21700
rect 25340 21646 25342 21698
rect 25342 21646 25394 21698
rect 25394 21646 25396 21698
rect 25340 21644 25396 21646
rect 25340 21420 25396 21476
rect 25788 21586 25844 21588
rect 25788 21534 25790 21586
rect 25790 21534 25842 21586
rect 25842 21534 25844 21586
rect 25788 21532 25844 21534
rect 26124 22092 26180 22148
rect 26236 24332 26292 24388
rect 26124 20914 26180 20916
rect 26124 20862 26126 20914
rect 26126 20862 26178 20914
rect 26178 20862 26180 20914
rect 26124 20860 26180 20862
rect 25404 20410 25460 20412
rect 25404 20358 25406 20410
rect 25406 20358 25458 20410
rect 25458 20358 25460 20410
rect 25404 20356 25460 20358
rect 25508 20410 25564 20412
rect 25508 20358 25510 20410
rect 25510 20358 25562 20410
rect 25562 20358 25564 20410
rect 25508 20356 25564 20358
rect 25612 20410 25668 20412
rect 25612 20358 25614 20410
rect 25614 20358 25666 20410
rect 25666 20358 25668 20410
rect 25612 20356 25668 20358
rect 25340 20242 25396 20244
rect 25340 20190 25342 20242
rect 25342 20190 25394 20242
rect 25394 20190 25396 20242
rect 25340 20188 25396 20190
rect 25676 20242 25732 20244
rect 25676 20190 25678 20242
rect 25678 20190 25730 20242
rect 25730 20190 25732 20242
rect 25676 20188 25732 20190
rect 25452 19292 25508 19348
rect 25004 19068 25060 19124
rect 26908 28140 26964 28196
rect 26908 27858 26964 27860
rect 26908 27806 26910 27858
rect 26910 27806 26962 27858
rect 26962 27806 26964 27858
rect 26908 27804 26964 27806
rect 26908 27468 26964 27524
rect 27356 27020 27412 27076
rect 27132 25900 27188 25956
rect 27356 25676 27412 25732
rect 27020 25340 27076 25396
rect 26348 21756 26404 21812
rect 26572 23548 26628 23604
rect 27020 24050 27076 24052
rect 27020 23998 27022 24050
rect 27022 23998 27074 24050
rect 27074 23998 27076 24050
rect 27020 23996 27076 23998
rect 26796 22258 26852 22260
rect 26796 22206 26798 22258
rect 26798 22206 26850 22258
rect 26850 22206 26852 22258
rect 26796 22204 26852 22206
rect 26908 23884 26964 23940
rect 26572 21420 26628 21476
rect 26796 21980 26852 22036
rect 26908 21084 26964 21140
rect 27020 23660 27076 23716
rect 27244 25506 27300 25508
rect 27244 25454 27246 25506
rect 27246 25454 27298 25506
rect 27298 25454 27300 25506
rect 27244 25452 27300 25454
rect 27244 24892 27300 24948
rect 28364 30156 28420 30212
rect 28476 30044 28532 30100
rect 28700 31164 28756 31220
rect 27692 28588 27748 28644
rect 27580 28364 27636 28420
rect 27804 26908 27860 26964
rect 27580 25228 27636 25284
rect 27468 25004 27524 25060
rect 27244 23826 27300 23828
rect 27244 23774 27246 23826
rect 27246 23774 27298 23826
rect 27298 23774 27300 23826
rect 27244 23772 27300 23774
rect 27356 23324 27412 23380
rect 27132 22764 27188 22820
rect 27244 22876 27300 22932
rect 27692 24668 27748 24724
rect 28140 27804 28196 27860
rect 28252 27580 28308 27636
rect 28588 28588 28644 28644
rect 28364 27356 28420 27412
rect 28476 27692 28532 27748
rect 28252 26684 28308 26740
rect 27692 23324 27748 23380
rect 27132 21980 27188 22036
rect 27244 21868 27300 21924
rect 27132 21420 27188 21476
rect 26796 20524 26852 20580
rect 26572 20300 26628 20356
rect 27020 20860 27076 20916
rect 27916 22764 27972 22820
rect 28364 25282 28420 25284
rect 28364 25230 28366 25282
rect 28366 25230 28418 25282
rect 28418 25230 28420 25282
rect 28364 25228 28420 25230
rect 29148 31106 29204 31108
rect 29148 31054 29150 31106
rect 29150 31054 29202 31106
rect 29202 31054 29204 31106
rect 29148 31052 29204 31054
rect 29260 30940 29316 30996
rect 30492 31052 30548 31108
rect 29436 30602 29492 30604
rect 29436 30550 29438 30602
rect 29438 30550 29490 30602
rect 29490 30550 29492 30602
rect 29436 30548 29492 30550
rect 29540 30602 29596 30604
rect 29540 30550 29542 30602
rect 29542 30550 29594 30602
rect 29594 30550 29596 30602
rect 29540 30548 29596 30550
rect 29644 30602 29700 30604
rect 29644 30550 29646 30602
rect 29646 30550 29698 30602
rect 29698 30550 29700 30602
rect 29644 30548 29700 30550
rect 29596 30210 29652 30212
rect 29596 30158 29598 30210
rect 29598 30158 29650 30210
rect 29650 30158 29652 30210
rect 29596 30156 29652 30158
rect 29436 29034 29492 29036
rect 29436 28982 29438 29034
rect 29438 28982 29490 29034
rect 29490 28982 29492 29034
rect 29436 28980 29492 28982
rect 29540 29034 29596 29036
rect 29540 28982 29542 29034
rect 29542 28982 29594 29034
rect 29594 28982 29596 29034
rect 29540 28980 29596 28982
rect 29644 29034 29700 29036
rect 29644 28982 29646 29034
rect 29646 28982 29698 29034
rect 29698 28982 29700 29034
rect 29644 28980 29700 28982
rect 29148 28700 29204 28756
rect 28700 25676 28756 25732
rect 29372 28530 29428 28532
rect 29372 28478 29374 28530
rect 29374 28478 29426 28530
rect 29426 28478 29428 28530
rect 29372 28476 29428 28478
rect 29596 28812 29652 28868
rect 28588 25394 28644 25396
rect 28588 25342 28590 25394
rect 28590 25342 28642 25394
rect 28642 25342 28644 25394
rect 28588 25340 28644 25342
rect 28700 25452 28756 25508
rect 28476 25116 28532 25172
rect 28476 23548 28532 23604
rect 28252 23154 28308 23156
rect 28252 23102 28254 23154
rect 28254 23102 28306 23154
rect 28306 23102 28308 23154
rect 28252 23100 28308 23102
rect 28140 22930 28196 22932
rect 28140 22878 28142 22930
rect 28142 22878 28194 22930
rect 28194 22878 28196 22930
rect 28140 22876 28196 22878
rect 28476 23324 28532 23380
rect 29484 28252 29540 28308
rect 29484 27916 29540 27972
rect 29436 27466 29492 27468
rect 29436 27414 29438 27466
rect 29438 27414 29490 27466
rect 29490 27414 29492 27466
rect 29436 27412 29492 27414
rect 29540 27466 29596 27468
rect 29540 27414 29542 27466
rect 29542 27414 29594 27466
rect 29594 27414 29596 27466
rect 29540 27412 29596 27414
rect 29644 27466 29700 27468
rect 29644 27414 29646 27466
rect 29646 27414 29698 27466
rect 29698 27414 29700 27466
rect 29644 27412 29700 27414
rect 29596 27074 29652 27076
rect 29596 27022 29598 27074
rect 29598 27022 29650 27074
rect 29650 27022 29652 27074
rect 29596 27020 29652 27022
rect 29260 26962 29316 26964
rect 29260 26910 29262 26962
rect 29262 26910 29314 26962
rect 29314 26910 29316 26962
rect 29260 26908 29316 26910
rect 29372 26684 29428 26740
rect 30156 28476 30212 28532
rect 30268 30156 30324 30212
rect 30380 29484 30436 29540
rect 30156 28252 30212 28308
rect 29148 26348 29204 26404
rect 29036 26290 29092 26292
rect 29036 26238 29038 26290
rect 29038 26238 29090 26290
rect 29090 26238 29092 26290
rect 29036 26236 29092 26238
rect 29036 26012 29092 26068
rect 29036 25788 29092 25844
rect 29484 26572 29540 26628
rect 29820 26572 29876 26628
rect 29484 26066 29540 26068
rect 29484 26014 29486 26066
rect 29486 26014 29538 26066
rect 29538 26014 29540 26066
rect 29484 26012 29540 26014
rect 29260 25788 29316 25844
rect 29436 25898 29492 25900
rect 29436 25846 29438 25898
rect 29438 25846 29490 25898
rect 29490 25846 29492 25898
rect 29436 25844 29492 25846
rect 29540 25898 29596 25900
rect 29540 25846 29542 25898
rect 29542 25846 29594 25898
rect 29594 25846 29596 25898
rect 29540 25844 29596 25846
rect 29644 25898 29700 25900
rect 29644 25846 29646 25898
rect 29646 25846 29698 25898
rect 29698 25846 29700 25898
rect 29644 25844 29700 25846
rect 29260 25564 29316 25620
rect 29036 25452 29092 25508
rect 29372 25228 29428 25284
rect 29596 24892 29652 24948
rect 28812 23996 28868 24052
rect 29148 23938 29204 23940
rect 29148 23886 29150 23938
rect 29150 23886 29202 23938
rect 29202 23886 29204 23938
rect 29148 23884 29204 23886
rect 29708 24668 29764 24724
rect 29436 24330 29492 24332
rect 29436 24278 29438 24330
rect 29438 24278 29490 24330
rect 29490 24278 29492 24330
rect 29436 24276 29492 24278
rect 29540 24330 29596 24332
rect 29540 24278 29542 24330
rect 29542 24278 29594 24330
rect 29594 24278 29596 24330
rect 29540 24276 29596 24278
rect 29644 24330 29700 24332
rect 29644 24278 29646 24330
rect 29646 24278 29698 24330
rect 29698 24278 29700 24330
rect 29644 24276 29700 24278
rect 29708 24108 29764 24164
rect 29372 23266 29428 23268
rect 29372 23214 29374 23266
rect 29374 23214 29426 23266
rect 29426 23214 29428 23266
rect 29372 23212 29428 23214
rect 29484 23100 29540 23156
rect 28364 22764 28420 22820
rect 27804 22428 27860 22484
rect 27468 21532 27524 21588
rect 27356 21196 27412 21252
rect 27244 20300 27300 20356
rect 26012 19794 26068 19796
rect 26012 19742 26014 19794
rect 26014 19742 26066 19794
rect 26066 19742 26068 19794
rect 26012 19740 26068 19742
rect 25788 19292 25844 19348
rect 26460 19516 26516 19572
rect 26236 19292 26292 19348
rect 24108 18620 24164 18676
rect 23436 18508 23492 18564
rect 23772 18508 23828 18564
rect 23212 17724 23268 17780
rect 23212 16828 23268 16884
rect 24780 17778 24836 17780
rect 24780 17726 24782 17778
rect 24782 17726 24834 17778
rect 24834 17726 24836 17778
rect 24780 17724 24836 17726
rect 24668 17612 24724 17668
rect 23884 17500 23940 17556
rect 23436 16828 23492 16884
rect 23548 16940 23604 16996
rect 23548 16770 23604 16772
rect 23548 16718 23550 16770
rect 23550 16718 23602 16770
rect 23602 16718 23604 16770
rect 23548 16716 23604 16718
rect 23212 15820 23268 15876
rect 22876 15538 22932 15540
rect 22876 15486 22878 15538
rect 22878 15486 22930 15538
rect 22930 15486 22932 15538
rect 22876 15484 22932 15486
rect 23548 16322 23604 16324
rect 23548 16270 23550 16322
rect 23550 16270 23602 16322
rect 23602 16270 23604 16322
rect 23548 16268 23604 16270
rect 23548 15426 23604 15428
rect 23548 15374 23550 15426
rect 23550 15374 23602 15426
rect 23602 15374 23604 15426
rect 23548 15372 23604 15374
rect 23884 15484 23940 15540
rect 22988 14924 23044 14980
rect 23884 15314 23940 15316
rect 23884 15262 23886 15314
rect 23886 15262 23938 15314
rect 23938 15262 23940 15314
rect 23884 15260 23940 15262
rect 24556 17442 24612 17444
rect 24556 17390 24558 17442
rect 24558 17390 24610 17442
rect 24610 17390 24612 17442
rect 24556 17388 24612 17390
rect 24444 16716 24500 16772
rect 24556 15932 24612 15988
rect 24108 15708 24164 15764
rect 24444 15372 24500 15428
rect 22876 14476 22932 14532
rect 23324 13916 23380 13972
rect 23100 13692 23156 13748
rect 23436 13804 23492 13860
rect 23772 14530 23828 14532
rect 23772 14478 23774 14530
rect 23774 14478 23826 14530
rect 23826 14478 23828 14530
rect 23772 14476 23828 14478
rect 23996 13916 24052 13972
rect 23772 13858 23828 13860
rect 23772 13806 23774 13858
rect 23774 13806 23826 13858
rect 23826 13806 23828 13858
rect 23772 13804 23828 13806
rect 23660 13692 23716 13748
rect 24668 15820 24724 15876
rect 24780 15260 24836 15316
rect 25404 18842 25460 18844
rect 25404 18790 25406 18842
rect 25406 18790 25458 18842
rect 25458 18790 25460 18842
rect 25404 18788 25460 18790
rect 25508 18842 25564 18844
rect 25508 18790 25510 18842
rect 25510 18790 25562 18842
rect 25562 18790 25564 18842
rect 25508 18788 25564 18790
rect 25612 18842 25668 18844
rect 25612 18790 25614 18842
rect 25614 18790 25666 18842
rect 25666 18790 25668 18842
rect 25612 18788 25668 18790
rect 25788 18844 25844 18900
rect 25004 18396 25060 18452
rect 25900 18450 25956 18452
rect 25900 18398 25902 18450
rect 25902 18398 25954 18450
rect 25954 18398 25956 18450
rect 25900 18396 25956 18398
rect 25452 18284 25508 18340
rect 25900 17612 25956 17668
rect 25340 17554 25396 17556
rect 25340 17502 25342 17554
rect 25342 17502 25394 17554
rect 25394 17502 25396 17554
rect 25340 17500 25396 17502
rect 25404 17274 25460 17276
rect 25404 17222 25406 17274
rect 25406 17222 25458 17274
rect 25458 17222 25460 17274
rect 25404 17220 25460 17222
rect 25508 17274 25564 17276
rect 25508 17222 25510 17274
rect 25510 17222 25562 17274
rect 25562 17222 25564 17274
rect 25508 17220 25564 17222
rect 25612 17274 25668 17276
rect 25612 17222 25614 17274
rect 25614 17222 25666 17274
rect 25666 17222 25668 17274
rect 25612 17220 25668 17222
rect 25116 16716 25172 16772
rect 25564 16658 25620 16660
rect 25564 16606 25566 16658
rect 25566 16606 25618 16658
rect 25618 16606 25620 16658
rect 25564 16604 25620 16606
rect 25116 16156 25172 16212
rect 24220 13916 24276 13972
rect 23772 13244 23828 13300
rect 23324 12962 23380 12964
rect 23324 12910 23326 12962
rect 23326 12910 23378 12962
rect 23378 12910 23380 12962
rect 23324 12908 23380 12910
rect 24220 13132 24276 13188
rect 23996 12962 24052 12964
rect 23996 12910 23998 12962
rect 23998 12910 24050 12962
rect 24050 12910 24052 12962
rect 23996 12908 24052 12910
rect 24556 12962 24612 12964
rect 24556 12910 24558 12962
rect 24558 12910 24610 12962
rect 24610 12910 24612 12962
rect 24556 12908 24612 12910
rect 23212 12402 23268 12404
rect 23212 12350 23214 12402
rect 23214 12350 23266 12402
rect 23266 12350 23268 12402
rect 23212 12348 23268 12350
rect 23884 12402 23940 12404
rect 23884 12350 23886 12402
rect 23886 12350 23938 12402
rect 23938 12350 23940 12402
rect 23884 12348 23940 12350
rect 22876 10780 22932 10836
rect 23324 10444 23380 10500
rect 22764 10108 22820 10164
rect 22988 10332 23044 10388
rect 22316 9266 22372 9268
rect 22316 9214 22318 9266
rect 22318 9214 22370 9266
rect 22370 9214 22372 9266
rect 22316 9212 22372 9214
rect 22540 9884 22596 9940
rect 24220 12290 24276 12292
rect 24220 12238 24222 12290
rect 24222 12238 24274 12290
rect 24274 12238 24276 12290
rect 24220 12236 24276 12238
rect 25004 15932 25060 15988
rect 26124 18508 26180 18564
rect 26460 18620 26516 18676
rect 26348 17724 26404 17780
rect 26236 17612 26292 17668
rect 26124 17500 26180 17556
rect 26124 17164 26180 17220
rect 26012 16994 26068 16996
rect 26012 16942 26014 16994
rect 26014 16942 26066 16994
rect 26066 16942 26068 16994
rect 26012 16940 26068 16942
rect 26124 16604 26180 16660
rect 25564 15874 25620 15876
rect 25564 15822 25566 15874
rect 25566 15822 25618 15874
rect 25618 15822 25620 15874
rect 25564 15820 25620 15822
rect 25116 15708 25172 15764
rect 25404 15706 25460 15708
rect 25404 15654 25406 15706
rect 25406 15654 25458 15706
rect 25458 15654 25460 15706
rect 25404 15652 25460 15654
rect 25508 15706 25564 15708
rect 25508 15654 25510 15706
rect 25510 15654 25562 15706
rect 25562 15654 25564 15706
rect 25508 15652 25564 15654
rect 25612 15706 25668 15708
rect 25612 15654 25614 15706
rect 25614 15654 25666 15706
rect 25666 15654 25668 15706
rect 25612 15652 25668 15654
rect 25116 15484 25172 15540
rect 25564 15484 25620 15540
rect 25788 15426 25844 15428
rect 25788 15374 25790 15426
rect 25790 15374 25842 15426
rect 25842 15374 25844 15426
rect 25788 15372 25844 15374
rect 25564 15260 25620 15316
rect 25676 14642 25732 14644
rect 25676 14590 25678 14642
rect 25678 14590 25730 14642
rect 25730 14590 25732 14642
rect 25676 14588 25732 14590
rect 25404 14138 25460 14140
rect 25404 14086 25406 14138
rect 25406 14086 25458 14138
rect 25458 14086 25460 14138
rect 25404 14084 25460 14086
rect 25508 14138 25564 14140
rect 25508 14086 25510 14138
rect 25510 14086 25562 14138
rect 25562 14086 25564 14138
rect 25508 14084 25564 14086
rect 25612 14138 25668 14140
rect 25612 14086 25614 14138
rect 25614 14086 25666 14138
rect 25666 14086 25668 14138
rect 25612 14084 25668 14086
rect 26012 15932 26068 15988
rect 26012 15596 26068 15652
rect 26124 15372 26180 15428
rect 25900 14364 25956 14420
rect 25452 13970 25508 13972
rect 25452 13918 25454 13970
rect 25454 13918 25506 13970
rect 25506 13918 25508 13970
rect 25452 13916 25508 13918
rect 25228 13580 25284 13636
rect 24892 13132 24948 13188
rect 26124 13020 26180 13076
rect 25228 12908 25284 12964
rect 24780 12460 24836 12516
rect 25404 12570 25460 12572
rect 25404 12518 25406 12570
rect 25406 12518 25458 12570
rect 25458 12518 25460 12570
rect 25404 12516 25460 12518
rect 25508 12570 25564 12572
rect 25508 12518 25510 12570
rect 25510 12518 25562 12570
rect 25562 12518 25564 12570
rect 25508 12516 25564 12518
rect 25612 12570 25668 12572
rect 25612 12518 25614 12570
rect 25614 12518 25666 12570
rect 25666 12518 25668 12570
rect 25612 12516 25668 12518
rect 25228 12236 25284 12292
rect 24556 10668 24612 10724
rect 25004 11282 25060 11284
rect 25004 11230 25006 11282
rect 25006 11230 25058 11282
rect 25058 11230 25060 11282
rect 25004 11228 25060 11230
rect 24668 10556 24724 10612
rect 23548 9884 23604 9940
rect 23884 10444 23940 10500
rect 25004 10220 25060 10276
rect 24892 10108 24948 10164
rect 24444 9826 24500 9828
rect 24444 9774 24446 9826
rect 24446 9774 24498 9826
rect 24498 9774 24500 9826
rect 24444 9772 24500 9774
rect 23324 9714 23380 9716
rect 23324 9662 23326 9714
rect 23326 9662 23378 9714
rect 23378 9662 23380 9714
rect 23324 9660 23380 9662
rect 24332 9714 24388 9716
rect 24332 9662 24334 9714
rect 24334 9662 24386 9714
rect 24386 9662 24388 9714
rect 24332 9660 24388 9662
rect 22540 8876 22596 8932
rect 22316 8370 22372 8372
rect 22316 8318 22318 8370
rect 22318 8318 22370 8370
rect 22370 8318 22372 8370
rect 22316 8316 22372 8318
rect 22092 8204 22148 8260
rect 22092 7586 22148 7588
rect 22092 7534 22094 7586
rect 22094 7534 22146 7586
rect 22146 7534 22148 7586
rect 22092 7532 22148 7534
rect 21756 6466 21812 6468
rect 21756 6414 21758 6466
rect 21758 6414 21810 6466
rect 21810 6414 21812 6466
rect 21756 6412 21812 6414
rect 21980 6412 22036 6468
rect 21868 5794 21924 5796
rect 21868 5742 21870 5794
rect 21870 5742 21922 5794
rect 21922 5742 21924 5794
rect 21868 5740 21924 5742
rect 21372 5514 21428 5516
rect 21372 5462 21374 5514
rect 21374 5462 21426 5514
rect 21426 5462 21428 5514
rect 21372 5460 21428 5462
rect 21476 5514 21532 5516
rect 21476 5462 21478 5514
rect 21478 5462 21530 5514
rect 21530 5462 21532 5514
rect 21476 5460 21532 5462
rect 21580 5514 21636 5516
rect 21580 5462 21582 5514
rect 21582 5462 21634 5514
rect 21634 5462 21636 5514
rect 21580 5460 21636 5462
rect 21084 3724 21140 3780
rect 21308 5180 21364 5236
rect 21644 5068 21700 5124
rect 21532 4172 21588 4228
rect 21372 3946 21428 3948
rect 21372 3894 21374 3946
rect 21374 3894 21426 3946
rect 21426 3894 21428 3946
rect 21372 3892 21428 3894
rect 21476 3946 21532 3948
rect 21476 3894 21478 3946
rect 21478 3894 21530 3946
rect 21530 3894 21532 3946
rect 21476 3892 21532 3894
rect 21580 3946 21636 3948
rect 21580 3894 21582 3946
rect 21582 3894 21634 3946
rect 21634 3894 21636 3946
rect 21580 3892 21636 3894
rect 22540 6748 22596 6804
rect 22204 6130 22260 6132
rect 22204 6078 22206 6130
rect 22206 6078 22258 6130
rect 22258 6078 22260 6130
rect 22204 6076 22260 6078
rect 22764 7474 22820 7476
rect 22764 7422 22766 7474
rect 22766 7422 22818 7474
rect 22818 7422 22820 7474
rect 22764 7420 22820 7422
rect 22652 6636 22708 6692
rect 22764 6412 22820 6468
rect 23772 9212 23828 9268
rect 23212 8764 23268 8820
rect 24332 9212 24388 9268
rect 24556 9154 24612 9156
rect 24556 9102 24558 9154
rect 24558 9102 24610 9154
rect 24610 9102 24612 9154
rect 24556 9100 24612 9102
rect 24444 8876 24500 8932
rect 23436 8428 23492 8484
rect 23324 7756 23380 7812
rect 23100 7474 23156 7476
rect 23100 7422 23102 7474
rect 23102 7422 23154 7474
rect 23154 7422 23156 7474
rect 23100 7420 23156 7422
rect 23436 7474 23492 7476
rect 23436 7422 23438 7474
rect 23438 7422 23490 7474
rect 23490 7422 23492 7474
rect 23436 7420 23492 7422
rect 23996 8034 24052 8036
rect 23996 7982 23998 8034
rect 23998 7982 24050 8034
rect 24050 7982 24052 8034
rect 23996 7980 24052 7982
rect 23660 7308 23716 7364
rect 24332 7980 24388 8036
rect 24668 7980 24724 8036
rect 24556 7420 24612 7476
rect 24332 7084 24388 7140
rect 24444 7308 24500 7364
rect 24220 6860 24276 6916
rect 22876 6300 22932 6356
rect 22652 5964 22708 6020
rect 22764 6188 22820 6244
rect 23436 6076 23492 6132
rect 23548 6300 23604 6356
rect 23100 5906 23156 5908
rect 23100 5854 23102 5906
rect 23102 5854 23154 5906
rect 23154 5854 23156 5906
rect 23100 5852 23156 5854
rect 24780 7420 24836 7476
rect 24668 7308 24724 7364
rect 24556 6748 24612 6804
rect 24220 6300 24276 6356
rect 24444 6300 24500 6356
rect 24780 6412 24836 6468
rect 24108 6188 24164 6244
rect 24332 6076 24388 6132
rect 22540 5234 22596 5236
rect 22540 5182 22542 5234
rect 22542 5182 22594 5234
rect 22594 5182 22596 5234
rect 22540 5180 22596 5182
rect 23324 5740 23380 5796
rect 23212 5068 23268 5124
rect 23660 5628 23716 5684
rect 22092 3836 22148 3892
rect 21868 3666 21924 3668
rect 21868 3614 21870 3666
rect 21870 3614 21922 3666
rect 21922 3614 21924 3666
rect 21868 3612 21924 3614
rect 22876 3388 22932 3444
rect 23996 4956 24052 5012
rect 24108 5516 24164 5572
rect 24556 5234 24612 5236
rect 24556 5182 24558 5234
rect 24558 5182 24610 5234
rect 24610 5182 24612 5234
rect 24556 5180 24612 5182
rect 24332 5122 24388 5124
rect 24332 5070 24334 5122
rect 24334 5070 24386 5122
rect 24386 5070 24388 5122
rect 24332 5068 24388 5070
rect 25340 12178 25396 12180
rect 25340 12126 25342 12178
rect 25342 12126 25394 12178
rect 25394 12126 25396 12178
rect 25340 12124 25396 12126
rect 25900 12738 25956 12740
rect 25900 12686 25902 12738
rect 25902 12686 25954 12738
rect 25954 12686 25956 12738
rect 25900 12684 25956 12686
rect 26908 19964 26964 20020
rect 26684 18956 26740 19012
rect 26796 18620 26852 18676
rect 27020 19906 27076 19908
rect 27020 19854 27022 19906
rect 27022 19854 27074 19906
rect 27074 19854 27076 19906
rect 27020 19852 27076 19854
rect 27132 19516 27188 19572
rect 27804 22204 27860 22260
rect 27692 21308 27748 21364
rect 27916 21868 27972 21924
rect 28140 22370 28196 22372
rect 28140 22318 28142 22370
rect 28142 22318 28194 22370
rect 28194 22318 28196 22370
rect 28140 22316 28196 22318
rect 28476 22258 28532 22260
rect 28476 22206 28478 22258
rect 28478 22206 28530 22258
rect 28530 22206 28532 22258
rect 28476 22204 28532 22206
rect 28252 21698 28308 21700
rect 28252 21646 28254 21698
rect 28254 21646 28306 21698
rect 28306 21646 28308 21698
rect 28252 21644 28308 21646
rect 28140 21420 28196 21476
rect 27580 20076 27636 20132
rect 27580 19516 27636 19572
rect 29932 23212 29988 23268
rect 30044 25452 30100 25508
rect 29708 22988 29764 23044
rect 29436 22762 29492 22764
rect 29436 22710 29438 22762
rect 29438 22710 29490 22762
rect 29490 22710 29492 22762
rect 29436 22708 29492 22710
rect 29540 22762 29596 22764
rect 29540 22710 29542 22762
rect 29542 22710 29594 22762
rect 29594 22710 29596 22762
rect 29540 22708 29596 22710
rect 29644 22762 29700 22764
rect 29644 22710 29646 22762
rect 29646 22710 29698 22762
rect 29698 22710 29700 22762
rect 29644 22708 29700 22710
rect 29484 22204 29540 22260
rect 28924 21196 28980 21252
rect 29148 20802 29204 20804
rect 29148 20750 29150 20802
rect 29150 20750 29202 20802
rect 29202 20750 29204 20802
rect 29148 20748 29204 20750
rect 28588 20636 28644 20692
rect 27916 19852 27972 19908
rect 27468 18844 27524 18900
rect 26908 18508 26964 18564
rect 26796 17666 26852 17668
rect 26796 17614 26798 17666
rect 26798 17614 26850 17666
rect 26850 17614 26852 17666
rect 26796 17612 26852 17614
rect 26572 17106 26628 17108
rect 26572 17054 26574 17106
rect 26574 17054 26626 17106
rect 26626 17054 26628 17106
rect 26572 17052 26628 17054
rect 27020 17276 27076 17332
rect 26684 16940 26740 16996
rect 26796 17052 26852 17108
rect 27692 18562 27748 18564
rect 27692 18510 27694 18562
rect 27694 18510 27746 18562
rect 27746 18510 27748 18562
rect 27692 18508 27748 18510
rect 27468 18172 27524 18228
rect 27244 17612 27300 17668
rect 27356 17388 27412 17444
rect 27132 17052 27188 17108
rect 27244 17276 27300 17332
rect 27020 16828 27076 16884
rect 26796 15372 26852 15428
rect 26460 15260 26516 15316
rect 26572 14700 26628 14756
rect 27356 16882 27412 16884
rect 27356 16830 27358 16882
rect 27358 16830 27410 16882
rect 27410 16830 27412 16882
rect 27356 16828 27412 16830
rect 27692 17388 27748 17444
rect 28028 19404 28084 19460
rect 27916 18674 27972 18676
rect 27916 18622 27918 18674
rect 27918 18622 27970 18674
rect 27970 18622 27972 18674
rect 27916 18620 27972 18622
rect 28364 19852 28420 19908
rect 28476 19180 28532 19236
rect 29820 21586 29876 21588
rect 29820 21534 29822 21586
rect 29822 21534 29874 21586
rect 29874 21534 29876 21586
rect 29820 21532 29876 21534
rect 29436 21194 29492 21196
rect 29436 21142 29438 21194
rect 29438 21142 29490 21194
rect 29490 21142 29492 21194
rect 29436 21140 29492 21142
rect 29540 21194 29596 21196
rect 29540 21142 29542 21194
rect 29542 21142 29594 21194
rect 29594 21142 29596 21194
rect 29540 21140 29596 21142
rect 29644 21194 29700 21196
rect 29644 21142 29646 21194
rect 29646 21142 29698 21194
rect 29698 21142 29700 21194
rect 29644 21140 29700 21142
rect 29260 20300 29316 20356
rect 29372 20972 29428 21028
rect 29372 19964 29428 20020
rect 29436 19626 29492 19628
rect 29436 19574 29438 19626
rect 29438 19574 29490 19626
rect 29490 19574 29492 19626
rect 29436 19572 29492 19574
rect 29540 19626 29596 19628
rect 29540 19574 29542 19626
rect 29542 19574 29594 19626
rect 29594 19574 29596 19626
rect 29540 19572 29596 19574
rect 29644 19626 29700 19628
rect 29644 19574 29646 19626
rect 29646 19574 29698 19626
rect 29698 19574 29700 19626
rect 29644 19572 29700 19574
rect 29148 19458 29204 19460
rect 29148 19406 29150 19458
rect 29150 19406 29202 19458
rect 29202 19406 29204 19458
rect 29148 19404 29204 19406
rect 29484 19404 29540 19460
rect 28700 19180 28756 19236
rect 28476 18844 28532 18900
rect 29932 20076 29988 20132
rect 29932 19628 29988 19684
rect 29148 18956 29204 19012
rect 28700 18620 28756 18676
rect 29596 18620 29652 18676
rect 28364 18508 28420 18564
rect 28252 18284 28308 18340
rect 26908 14700 26964 14756
rect 27916 17612 27972 17668
rect 26908 14028 26964 14084
rect 26572 13746 26628 13748
rect 26572 13694 26574 13746
rect 26574 13694 26626 13746
rect 26626 13694 26628 13746
rect 26572 13692 26628 13694
rect 26684 13244 26740 13300
rect 26460 13074 26516 13076
rect 26460 13022 26462 13074
rect 26462 13022 26514 13074
rect 26514 13022 26516 13074
rect 26460 13020 26516 13022
rect 26684 13020 26740 13076
rect 26572 12850 26628 12852
rect 26572 12798 26574 12850
rect 26574 12798 26626 12850
rect 26626 12798 26628 12850
rect 26572 12796 26628 12798
rect 26348 12738 26404 12740
rect 26348 12686 26350 12738
rect 26350 12686 26402 12738
rect 26402 12686 26404 12738
rect 26348 12684 26404 12686
rect 27244 12572 27300 12628
rect 25900 11788 25956 11844
rect 27468 15708 27524 15764
rect 27804 16770 27860 16772
rect 27804 16718 27806 16770
rect 27806 16718 27858 16770
rect 27858 16718 27860 16770
rect 27804 16716 27860 16718
rect 27580 14812 27636 14868
rect 27468 13746 27524 13748
rect 27468 13694 27470 13746
rect 27470 13694 27522 13746
rect 27522 13694 27524 13746
rect 27468 13692 27524 13694
rect 26012 11564 26068 11620
rect 25452 11228 25508 11284
rect 25404 11002 25460 11004
rect 25404 10950 25406 11002
rect 25406 10950 25458 11002
rect 25458 10950 25460 11002
rect 25404 10948 25460 10950
rect 25508 11002 25564 11004
rect 25508 10950 25510 11002
rect 25510 10950 25562 11002
rect 25562 10950 25564 11002
rect 25508 10948 25564 10950
rect 25612 11002 25668 11004
rect 25612 10950 25614 11002
rect 25614 10950 25666 11002
rect 25666 10950 25668 11002
rect 25612 10948 25668 10950
rect 27356 11788 27412 11844
rect 25564 10668 25620 10724
rect 25452 10610 25508 10612
rect 25452 10558 25454 10610
rect 25454 10558 25506 10610
rect 25506 10558 25508 10610
rect 25452 10556 25508 10558
rect 25340 10498 25396 10500
rect 25340 10446 25342 10498
rect 25342 10446 25394 10498
rect 25394 10446 25396 10498
rect 25340 10444 25396 10446
rect 25228 9996 25284 10052
rect 25452 9884 25508 9940
rect 26460 10722 26516 10724
rect 26460 10670 26462 10722
rect 26462 10670 26514 10722
rect 26514 10670 26516 10722
rect 26460 10668 26516 10670
rect 26012 10444 26068 10500
rect 25228 9714 25284 9716
rect 25228 9662 25230 9714
rect 25230 9662 25282 9714
rect 25282 9662 25284 9714
rect 25228 9660 25284 9662
rect 25340 9548 25396 9604
rect 25676 9602 25732 9604
rect 25676 9550 25678 9602
rect 25678 9550 25730 9602
rect 25730 9550 25732 9602
rect 25676 9548 25732 9550
rect 25404 9434 25460 9436
rect 25404 9382 25406 9434
rect 25406 9382 25458 9434
rect 25458 9382 25460 9434
rect 25404 9380 25460 9382
rect 25508 9434 25564 9436
rect 25508 9382 25510 9434
rect 25510 9382 25562 9434
rect 25562 9382 25564 9434
rect 25508 9380 25564 9382
rect 25612 9434 25668 9436
rect 25612 9382 25614 9434
rect 25614 9382 25666 9434
rect 25666 9382 25668 9434
rect 25612 9380 25668 9382
rect 25564 9266 25620 9268
rect 25564 9214 25566 9266
rect 25566 9214 25618 9266
rect 25618 9214 25620 9266
rect 25564 9212 25620 9214
rect 25116 8652 25172 8708
rect 25340 8652 25396 8708
rect 25900 9436 25956 9492
rect 25788 8316 25844 8372
rect 26348 10556 26404 10612
rect 26572 10556 26628 10612
rect 26124 9100 26180 9156
rect 25404 7866 25460 7868
rect 25404 7814 25406 7866
rect 25406 7814 25458 7866
rect 25458 7814 25460 7866
rect 25404 7812 25460 7814
rect 25508 7866 25564 7868
rect 25508 7814 25510 7866
rect 25510 7814 25562 7866
rect 25562 7814 25564 7866
rect 25508 7812 25564 7814
rect 25612 7866 25668 7868
rect 25612 7814 25614 7866
rect 25614 7814 25666 7866
rect 25666 7814 25668 7866
rect 25612 7812 25668 7814
rect 25116 7644 25172 7700
rect 25228 7308 25284 7364
rect 24892 6188 24948 6244
rect 24444 4508 24500 4564
rect 25340 6466 25396 6468
rect 25340 6414 25342 6466
rect 25342 6414 25394 6466
rect 25394 6414 25396 6466
rect 25340 6412 25396 6414
rect 25004 4396 25060 4452
rect 25116 6188 25172 6244
rect 23996 3442 24052 3444
rect 23996 3390 23998 3442
rect 23998 3390 24050 3442
rect 24050 3390 24052 3442
rect 23996 3388 24052 3390
rect 24668 4226 24724 4228
rect 24668 4174 24670 4226
rect 24670 4174 24722 4226
rect 24722 4174 24724 4226
rect 24668 4172 24724 4174
rect 24780 3500 24836 3556
rect 25900 6860 25956 6916
rect 26684 9884 26740 9940
rect 26572 9548 26628 9604
rect 27244 11452 27300 11508
rect 27132 10610 27188 10612
rect 27132 10558 27134 10610
rect 27134 10558 27186 10610
rect 27186 10558 27188 10610
rect 27132 10556 27188 10558
rect 27020 9996 27076 10052
rect 27132 9938 27188 9940
rect 27132 9886 27134 9938
rect 27134 9886 27186 9938
rect 27186 9886 27188 9938
rect 27132 9884 27188 9886
rect 28140 17666 28196 17668
rect 28140 17614 28142 17666
rect 28142 17614 28194 17666
rect 28194 17614 28196 17666
rect 28140 17612 28196 17614
rect 28140 17276 28196 17332
rect 28588 18396 28644 18452
rect 28700 18060 28756 18116
rect 28812 18172 28868 18228
rect 28588 17948 28644 18004
rect 28476 17612 28532 17668
rect 28252 17164 28308 17220
rect 28476 17388 28532 17444
rect 28364 17106 28420 17108
rect 28364 17054 28366 17106
rect 28366 17054 28418 17106
rect 28418 17054 28420 17106
rect 28364 17052 28420 17054
rect 27916 15148 27972 15204
rect 27916 13858 27972 13860
rect 27916 13806 27918 13858
rect 27918 13806 27970 13858
rect 27970 13806 27972 13858
rect 27916 13804 27972 13806
rect 27804 13468 27860 13524
rect 28252 16098 28308 16100
rect 28252 16046 28254 16098
rect 28254 16046 28306 16098
rect 28306 16046 28308 16098
rect 28252 16044 28308 16046
rect 28252 15708 28308 15764
rect 28700 16156 28756 16212
rect 29484 18396 29540 18452
rect 29260 18338 29316 18340
rect 29260 18286 29262 18338
rect 29262 18286 29314 18338
rect 29314 18286 29316 18338
rect 29260 18284 29316 18286
rect 30380 28364 30436 28420
rect 30268 24108 30324 24164
rect 30268 23938 30324 23940
rect 30268 23886 30270 23938
rect 30270 23886 30322 23938
rect 30322 23886 30324 23938
rect 30268 23884 30324 23886
rect 30268 22370 30324 22372
rect 30268 22318 30270 22370
rect 30270 22318 30322 22370
rect 30322 22318 30324 22370
rect 30268 22316 30324 22318
rect 30268 21586 30324 21588
rect 30268 21534 30270 21586
rect 30270 21534 30322 21586
rect 30322 21534 30324 21586
rect 30268 21532 30324 21534
rect 30604 30044 30660 30100
rect 30492 23324 30548 23380
rect 30604 28140 30660 28196
rect 30828 28476 30884 28532
rect 30716 24892 30772 24948
rect 31052 30268 31108 30324
rect 32172 30882 32228 30884
rect 32172 30830 32174 30882
rect 32174 30830 32226 30882
rect 32226 30830 32228 30882
rect 32172 30828 32228 30830
rect 31276 30268 31332 30324
rect 32172 30268 32228 30324
rect 31388 29596 31444 29652
rect 31276 28812 31332 28868
rect 31276 28588 31332 28644
rect 31052 26012 31108 26068
rect 31276 24892 31332 24948
rect 31948 29426 32004 29428
rect 31948 29374 31950 29426
rect 31950 29374 32002 29426
rect 32002 29374 32004 29426
rect 31948 29372 32004 29374
rect 32732 30994 32788 30996
rect 32732 30942 32734 30994
rect 32734 30942 32786 30994
rect 32786 30942 32788 30994
rect 32732 30940 32788 30942
rect 33468 31386 33524 31388
rect 33468 31334 33470 31386
rect 33470 31334 33522 31386
rect 33522 31334 33524 31386
rect 33468 31332 33524 31334
rect 33572 31386 33628 31388
rect 33572 31334 33574 31386
rect 33574 31334 33626 31386
rect 33626 31334 33628 31386
rect 33572 31332 33628 31334
rect 33676 31386 33732 31388
rect 33676 31334 33678 31386
rect 33678 31334 33730 31386
rect 33730 31334 33732 31386
rect 33676 31332 33732 31334
rect 32956 30770 33012 30772
rect 32956 30718 32958 30770
rect 32958 30718 33010 30770
rect 33010 30718 33012 30770
rect 32956 30716 33012 30718
rect 32844 30380 32900 30436
rect 32508 29596 32564 29652
rect 32396 29036 32452 29092
rect 33180 29314 33236 29316
rect 33180 29262 33182 29314
rect 33182 29262 33234 29314
rect 33234 29262 33236 29314
rect 33180 29260 33236 29262
rect 33068 28924 33124 28980
rect 32284 28812 32340 28868
rect 33180 28754 33236 28756
rect 33180 28702 33182 28754
rect 33182 28702 33234 28754
rect 33234 28702 33236 28754
rect 33180 28700 33236 28702
rect 33180 27580 33236 27636
rect 31948 24610 32004 24612
rect 31948 24558 31950 24610
rect 31950 24558 32002 24610
rect 32002 24558 32004 24610
rect 31948 24556 32004 24558
rect 30268 20076 30324 20132
rect 30268 19068 30324 19124
rect 30156 18844 30212 18900
rect 29932 18508 29988 18564
rect 30492 18732 30548 18788
rect 30604 19180 30660 19236
rect 29708 18284 29764 18340
rect 29820 18226 29876 18228
rect 29820 18174 29822 18226
rect 29822 18174 29874 18226
rect 29874 18174 29876 18226
rect 29820 18172 29876 18174
rect 29436 18058 29492 18060
rect 29436 18006 29438 18058
rect 29438 18006 29490 18058
rect 29490 18006 29492 18058
rect 29436 18004 29492 18006
rect 29540 18058 29596 18060
rect 29540 18006 29542 18058
rect 29542 18006 29594 18058
rect 29594 18006 29596 18058
rect 29540 18004 29596 18006
rect 29644 18058 29700 18060
rect 29644 18006 29646 18058
rect 29646 18006 29698 18058
rect 29698 18006 29700 18058
rect 29644 18004 29700 18006
rect 29260 17612 29316 17668
rect 29372 17836 29428 17892
rect 29372 16994 29428 16996
rect 29372 16942 29374 16994
rect 29374 16942 29426 16994
rect 29426 16942 29428 16994
rect 29372 16940 29428 16942
rect 29820 17052 29876 17108
rect 28924 16044 28980 16100
rect 28476 15596 28532 15652
rect 28476 15314 28532 15316
rect 28476 15262 28478 15314
rect 28478 15262 28530 15314
rect 28530 15262 28532 15314
rect 28476 15260 28532 15262
rect 28364 14924 28420 14980
rect 28252 14588 28308 14644
rect 28588 14924 28644 14980
rect 28700 15426 28756 15428
rect 28700 15374 28702 15426
rect 28702 15374 28754 15426
rect 28754 15374 28756 15426
rect 28700 15372 28756 15374
rect 28364 13580 28420 13636
rect 28476 14812 28532 14868
rect 28588 14700 28644 14756
rect 28588 13692 28644 13748
rect 27468 10556 27524 10612
rect 26908 9212 26964 9268
rect 27468 9602 27524 9604
rect 27468 9550 27470 9602
rect 27470 9550 27522 9602
rect 27522 9550 27524 9602
rect 27468 9548 27524 9550
rect 26236 8258 26292 8260
rect 26236 8206 26238 8258
rect 26238 8206 26290 8258
rect 26290 8206 26292 8258
rect 26236 8204 26292 8206
rect 26796 8034 26852 8036
rect 26796 7982 26798 8034
rect 26798 7982 26850 8034
rect 26850 7982 26852 8034
rect 26796 7980 26852 7982
rect 27692 12738 27748 12740
rect 27692 12686 27694 12738
rect 27694 12686 27746 12738
rect 27746 12686 27748 12738
rect 27692 12684 27748 12686
rect 28028 12012 28084 12068
rect 28476 13132 28532 13188
rect 29436 16490 29492 16492
rect 29436 16438 29438 16490
rect 29438 16438 29490 16490
rect 29490 16438 29492 16490
rect 29436 16436 29492 16438
rect 29540 16490 29596 16492
rect 29540 16438 29542 16490
rect 29542 16438 29594 16490
rect 29594 16438 29596 16490
rect 29540 16436 29596 16438
rect 29644 16490 29700 16492
rect 29644 16438 29646 16490
rect 29646 16438 29698 16490
rect 29698 16438 29700 16490
rect 29644 16436 29700 16438
rect 29372 16098 29428 16100
rect 29372 16046 29374 16098
rect 29374 16046 29426 16098
rect 29426 16046 29428 16098
rect 29372 16044 29428 16046
rect 29260 15708 29316 15764
rect 29036 14252 29092 14308
rect 28924 13468 28980 13524
rect 29436 14922 29492 14924
rect 29436 14870 29438 14922
rect 29438 14870 29490 14922
rect 29490 14870 29492 14922
rect 29436 14868 29492 14870
rect 29540 14922 29596 14924
rect 29540 14870 29542 14922
rect 29542 14870 29594 14922
rect 29594 14870 29596 14922
rect 29540 14868 29596 14870
rect 29644 14922 29700 14924
rect 29644 14870 29646 14922
rect 29646 14870 29698 14922
rect 29698 14870 29700 14922
rect 29644 14868 29700 14870
rect 30268 18060 30324 18116
rect 30044 17612 30100 17668
rect 30940 22316 30996 22372
rect 31948 23884 32004 23940
rect 31052 20300 31108 20356
rect 31052 20018 31108 20020
rect 31052 19966 31054 20018
rect 31054 19966 31106 20018
rect 31106 19966 31108 20018
rect 31052 19964 31108 19966
rect 30492 17164 30548 17220
rect 30268 16770 30324 16772
rect 30268 16718 30270 16770
rect 30270 16718 30322 16770
rect 30322 16718 30324 16770
rect 30268 16716 30324 16718
rect 29932 15484 29988 15540
rect 29708 14306 29764 14308
rect 29708 14254 29710 14306
rect 29710 14254 29762 14306
rect 29762 14254 29764 14306
rect 29708 14252 29764 14254
rect 29820 14140 29876 14196
rect 30268 15596 30324 15652
rect 30940 18450 30996 18452
rect 30940 18398 30942 18450
rect 30942 18398 30994 18450
rect 30994 18398 30996 18450
rect 30940 18396 30996 18398
rect 31052 18284 31108 18340
rect 30380 15202 30436 15204
rect 30380 15150 30382 15202
rect 30382 15150 30434 15202
rect 30434 15150 30436 15202
rect 30380 15148 30436 15150
rect 30044 14140 30100 14196
rect 29596 13634 29652 13636
rect 29596 13582 29598 13634
rect 29598 13582 29650 13634
rect 29650 13582 29652 13634
rect 29596 13580 29652 13582
rect 29820 13468 29876 13524
rect 29436 13354 29492 13356
rect 29436 13302 29438 13354
rect 29438 13302 29490 13354
rect 29490 13302 29492 13354
rect 29436 13300 29492 13302
rect 29540 13354 29596 13356
rect 29540 13302 29542 13354
rect 29542 13302 29594 13354
rect 29594 13302 29596 13354
rect 29540 13300 29596 13302
rect 29644 13354 29700 13356
rect 29644 13302 29646 13354
rect 29646 13302 29698 13354
rect 29698 13302 29700 13354
rect 29644 13300 29700 13302
rect 28700 12684 28756 12740
rect 28700 12460 28756 12516
rect 29148 12684 29204 12740
rect 28588 11900 28644 11956
rect 28252 11452 28308 11508
rect 28364 11228 28420 11284
rect 28252 11170 28308 11172
rect 28252 11118 28254 11170
rect 28254 11118 28306 11170
rect 28306 11118 28308 11170
rect 28252 11116 28308 11118
rect 28140 9826 28196 9828
rect 28140 9774 28142 9826
rect 28142 9774 28194 9826
rect 28194 9774 28196 9826
rect 28140 9772 28196 9774
rect 28028 9100 28084 9156
rect 26796 7644 26852 7700
rect 26684 7586 26740 7588
rect 26684 7534 26686 7586
rect 26686 7534 26738 7586
rect 26738 7534 26740 7586
rect 26684 7532 26740 7534
rect 26908 7420 26964 7476
rect 26460 6860 26516 6916
rect 25676 6690 25732 6692
rect 25676 6638 25678 6690
rect 25678 6638 25730 6690
rect 25730 6638 25732 6690
rect 25676 6636 25732 6638
rect 25564 6412 25620 6468
rect 25404 6298 25460 6300
rect 25404 6246 25406 6298
rect 25406 6246 25458 6298
rect 25458 6246 25460 6298
rect 25404 6244 25460 6246
rect 25508 6298 25564 6300
rect 25508 6246 25510 6298
rect 25510 6246 25562 6298
rect 25562 6246 25564 6298
rect 25508 6244 25564 6246
rect 25612 6298 25668 6300
rect 25612 6246 25614 6298
rect 25614 6246 25666 6298
rect 25666 6246 25668 6298
rect 25612 6244 25668 6246
rect 26348 6690 26404 6692
rect 26348 6638 26350 6690
rect 26350 6638 26402 6690
rect 26402 6638 26404 6690
rect 26348 6636 26404 6638
rect 26012 6076 26068 6132
rect 26348 6076 26404 6132
rect 25340 5906 25396 5908
rect 25340 5854 25342 5906
rect 25342 5854 25394 5906
rect 25394 5854 25396 5906
rect 25340 5852 25396 5854
rect 25676 5852 25732 5908
rect 25340 5122 25396 5124
rect 25340 5070 25342 5122
rect 25342 5070 25394 5122
rect 25394 5070 25396 5122
rect 25340 5068 25396 5070
rect 26348 5906 26404 5908
rect 26348 5854 26350 5906
rect 26350 5854 26402 5906
rect 26402 5854 26404 5906
rect 26348 5852 26404 5854
rect 25564 4898 25620 4900
rect 25564 4846 25566 4898
rect 25566 4846 25618 4898
rect 25618 4846 25620 4898
rect 25564 4844 25620 4846
rect 25404 4730 25460 4732
rect 25404 4678 25406 4730
rect 25406 4678 25458 4730
rect 25458 4678 25460 4730
rect 25404 4676 25460 4678
rect 25508 4730 25564 4732
rect 25508 4678 25510 4730
rect 25510 4678 25562 4730
rect 25562 4678 25564 4730
rect 25508 4676 25564 4678
rect 25612 4730 25668 4732
rect 25612 4678 25614 4730
rect 25614 4678 25666 4730
rect 25666 4678 25668 4730
rect 25612 4676 25668 4678
rect 25340 4508 25396 4564
rect 26460 5404 26516 5460
rect 26348 5292 26404 5348
rect 25564 4284 25620 4340
rect 26348 4284 26404 4340
rect 26236 4172 26292 4228
rect 25900 3442 25956 3444
rect 25900 3390 25902 3442
rect 25902 3390 25954 3442
rect 25954 3390 25956 3442
rect 25900 3388 25956 3390
rect 26796 6748 26852 6804
rect 27132 7420 27188 7476
rect 28140 8258 28196 8260
rect 28140 8206 28142 8258
rect 28142 8206 28194 8258
rect 28194 8206 28196 8258
rect 28140 8204 28196 8206
rect 27020 6972 27076 7028
rect 26684 6412 26740 6468
rect 26796 6076 26852 6132
rect 28700 10332 28756 10388
rect 29596 12908 29652 12964
rect 28924 12178 28980 12180
rect 28924 12126 28926 12178
rect 28926 12126 28978 12178
rect 28978 12126 28980 12178
rect 28924 12124 28980 12126
rect 29036 12066 29092 12068
rect 29036 12014 29038 12066
rect 29038 12014 29090 12066
rect 29090 12014 29092 12066
rect 29036 12012 29092 12014
rect 28812 10780 28868 10836
rect 28588 9212 28644 9268
rect 29436 11786 29492 11788
rect 29436 11734 29438 11786
rect 29438 11734 29490 11786
rect 29490 11734 29492 11786
rect 29436 11732 29492 11734
rect 29540 11786 29596 11788
rect 29540 11734 29542 11786
rect 29542 11734 29594 11786
rect 29594 11734 29596 11786
rect 29540 11732 29596 11734
rect 29644 11786 29700 11788
rect 29644 11734 29646 11786
rect 29646 11734 29698 11786
rect 29698 11734 29700 11786
rect 29644 11732 29700 11734
rect 29372 11116 29428 11172
rect 29260 10444 29316 10500
rect 29436 10218 29492 10220
rect 29436 10166 29438 10218
rect 29438 10166 29490 10218
rect 29490 10166 29492 10218
rect 29436 10164 29492 10166
rect 29540 10218 29596 10220
rect 29540 10166 29542 10218
rect 29542 10166 29594 10218
rect 29594 10166 29596 10218
rect 29540 10164 29596 10166
rect 29644 10218 29700 10220
rect 29644 10166 29646 10218
rect 29646 10166 29698 10218
rect 29698 10166 29700 10218
rect 29644 10164 29700 10166
rect 30156 13132 30212 13188
rect 30156 12796 30212 12852
rect 29932 11452 29988 11508
rect 30044 12460 30100 12516
rect 29932 11282 29988 11284
rect 29932 11230 29934 11282
rect 29934 11230 29986 11282
rect 29986 11230 29988 11282
rect 29932 11228 29988 11230
rect 29148 9996 29204 10052
rect 29260 9714 29316 9716
rect 29260 9662 29262 9714
rect 29262 9662 29314 9714
rect 29314 9662 29316 9714
rect 29260 9660 29316 9662
rect 29260 9266 29316 9268
rect 29260 9214 29262 9266
rect 29262 9214 29314 9266
rect 29314 9214 29316 9266
rect 29260 9212 29316 9214
rect 29596 9602 29652 9604
rect 29596 9550 29598 9602
rect 29598 9550 29650 9602
rect 29650 9550 29652 9602
rect 29596 9548 29652 9550
rect 29148 9154 29204 9156
rect 29148 9102 29150 9154
rect 29150 9102 29202 9154
rect 29202 9102 29204 9154
rect 29148 9100 29204 9102
rect 29436 8650 29492 8652
rect 29436 8598 29438 8650
rect 29438 8598 29490 8650
rect 29490 8598 29492 8650
rect 29436 8596 29492 8598
rect 29540 8650 29596 8652
rect 29540 8598 29542 8650
rect 29542 8598 29594 8650
rect 29594 8598 29596 8650
rect 29540 8596 29596 8598
rect 29644 8650 29700 8652
rect 29644 8598 29646 8650
rect 29646 8598 29698 8650
rect 29698 8598 29700 8650
rect 29644 8596 29700 8598
rect 29484 8428 29540 8484
rect 28588 7980 28644 8036
rect 29148 7644 29204 7700
rect 27692 7420 27748 7476
rect 28588 7586 28644 7588
rect 28588 7534 28590 7586
rect 28590 7534 28642 7586
rect 28642 7534 28644 7586
rect 28588 7532 28644 7534
rect 28924 7586 28980 7588
rect 28924 7534 28926 7586
rect 28926 7534 28978 7586
rect 28978 7534 28980 7586
rect 28924 7532 28980 7534
rect 27692 6972 27748 7028
rect 27580 6300 27636 6356
rect 26908 5404 26964 5460
rect 26796 5346 26852 5348
rect 26796 5294 26798 5346
rect 26798 5294 26850 5346
rect 26850 5294 26852 5346
rect 26796 5292 26852 5294
rect 28252 6972 28308 7028
rect 28140 6748 28196 6804
rect 27356 5292 27412 5348
rect 27692 5852 27748 5908
rect 26684 4508 26740 4564
rect 28028 5628 28084 5684
rect 28028 5122 28084 5124
rect 28028 5070 28030 5122
rect 28030 5070 28082 5122
rect 28082 5070 28084 5122
rect 28028 5068 28084 5070
rect 28252 6130 28308 6132
rect 28252 6078 28254 6130
rect 28254 6078 28306 6130
rect 28306 6078 28308 6130
rect 28252 6076 28308 6078
rect 28700 6860 28756 6916
rect 28476 6188 28532 6244
rect 28588 6300 28644 6356
rect 28812 5906 28868 5908
rect 28812 5854 28814 5906
rect 28814 5854 28866 5906
rect 28866 5854 28868 5906
rect 28812 5852 28868 5854
rect 28364 5292 28420 5348
rect 28588 5292 28644 5348
rect 29148 7420 29204 7476
rect 29148 6188 29204 6244
rect 29436 7082 29492 7084
rect 29436 7030 29438 7082
rect 29438 7030 29490 7082
rect 29490 7030 29492 7082
rect 29436 7028 29492 7030
rect 29540 7082 29596 7084
rect 29540 7030 29542 7082
rect 29542 7030 29594 7082
rect 29594 7030 29596 7082
rect 29540 7028 29596 7030
rect 29644 7082 29700 7084
rect 29644 7030 29646 7082
rect 29646 7030 29698 7082
rect 29698 7030 29700 7082
rect 29644 7028 29700 7030
rect 30156 11900 30212 11956
rect 30156 11116 30212 11172
rect 31500 20076 31556 20132
rect 31612 19404 31668 19460
rect 31276 18732 31332 18788
rect 31164 17164 31220 17220
rect 31500 17836 31556 17892
rect 31500 16828 31556 16884
rect 30828 15148 30884 15204
rect 30604 14252 30660 14308
rect 31164 14028 31220 14084
rect 33068 27244 33124 27300
rect 33180 26178 33236 26180
rect 33180 26126 33182 26178
rect 33182 26126 33234 26178
rect 33234 26126 33236 26178
rect 33180 26124 33236 26126
rect 33180 25618 33236 25620
rect 33180 25566 33182 25618
rect 33182 25566 33234 25618
rect 33234 25566 33236 25618
rect 33180 25564 33236 25566
rect 32508 24722 32564 24724
rect 32508 24670 32510 24722
rect 32510 24670 32562 24722
rect 32562 24670 32564 24722
rect 32508 24668 32564 24670
rect 32172 20524 32228 20580
rect 32060 20188 32116 20244
rect 32172 19852 32228 19908
rect 32060 18844 32116 18900
rect 31724 18060 31780 18116
rect 31724 14476 31780 14532
rect 31724 13970 31780 13972
rect 31724 13918 31726 13970
rect 31726 13918 31778 13970
rect 31778 13918 31780 13970
rect 31724 13916 31780 13918
rect 30828 13692 30884 13748
rect 30492 10108 30548 10164
rect 30604 13580 30660 13636
rect 30716 13074 30772 13076
rect 30716 13022 30718 13074
rect 30718 13022 30770 13074
rect 30770 13022 30772 13074
rect 30716 13020 30772 13022
rect 30716 12572 30772 12628
rect 32172 18620 32228 18676
rect 33180 24444 33236 24500
rect 32732 23884 32788 23940
rect 32396 21420 32452 21476
rect 32620 22876 32676 22932
rect 32396 20690 32452 20692
rect 32396 20638 32398 20690
rect 32398 20638 32450 20690
rect 32450 20638 32452 20690
rect 32396 20636 32452 20638
rect 32620 21868 32676 21924
rect 32508 18396 32564 18452
rect 32060 17500 32116 17556
rect 31948 16940 32004 16996
rect 33180 23266 33236 23268
rect 33180 23214 33182 23266
rect 33182 23214 33234 23266
rect 33234 23214 33236 23266
rect 33180 23212 33236 23214
rect 33068 22930 33124 22932
rect 33068 22878 33070 22930
rect 33070 22878 33122 22930
rect 33122 22878 33124 22930
rect 33068 22876 33124 22878
rect 32732 20076 32788 20132
rect 33468 29818 33524 29820
rect 33468 29766 33470 29818
rect 33470 29766 33522 29818
rect 33522 29766 33524 29818
rect 33468 29764 33524 29766
rect 33572 29818 33628 29820
rect 33572 29766 33574 29818
rect 33574 29766 33626 29818
rect 33626 29766 33628 29818
rect 33572 29764 33628 29766
rect 33676 29818 33732 29820
rect 33676 29766 33678 29818
rect 33678 29766 33730 29818
rect 33730 29766 33732 29818
rect 33676 29764 33732 29766
rect 34076 28588 34132 28644
rect 33468 28250 33524 28252
rect 33468 28198 33470 28250
rect 33470 28198 33522 28250
rect 33522 28198 33524 28250
rect 33468 28196 33524 28198
rect 33572 28250 33628 28252
rect 33572 28198 33574 28250
rect 33574 28198 33626 28250
rect 33626 28198 33628 28250
rect 33572 28196 33628 28198
rect 33676 28250 33732 28252
rect 33676 28198 33678 28250
rect 33678 28198 33730 28250
rect 33730 28198 33732 28250
rect 33676 28196 33732 28198
rect 33468 26682 33524 26684
rect 33468 26630 33470 26682
rect 33470 26630 33522 26682
rect 33522 26630 33524 26682
rect 33468 26628 33524 26630
rect 33572 26682 33628 26684
rect 33572 26630 33574 26682
rect 33574 26630 33626 26682
rect 33626 26630 33628 26682
rect 33572 26628 33628 26630
rect 33676 26682 33732 26684
rect 33676 26630 33678 26682
rect 33678 26630 33730 26682
rect 33730 26630 33732 26682
rect 33676 26628 33732 26630
rect 33852 26124 33908 26180
rect 33468 25114 33524 25116
rect 33468 25062 33470 25114
rect 33470 25062 33522 25114
rect 33522 25062 33524 25114
rect 33468 25060 33524 25062
rect 33572 25114 33628 25116
rect 33572 25062 33574 25114
rect 33574 25062 33626 25114
rect 33626 25062 33628 25114
rect 33572 25060 33628 25062
rect 33676 25114 33732 25116
rect 33676 25062 33678 25114
rect 33678 25062 33730 25114
rect 33730 25062 33732 25114
rect 33676 25060 33732 25062
rect 33468 23546 33524 23548
rect 33468 23494 33470 23546
rect 33470 23494 33522 23546
rect 33522 23494 33524 23546
rect 33468 23492 33524 23494
rect 33572 23546 33628 23548
rect 33572 23494 33574 23546
rect 33574 23494 33626 23546
rect 33626 23494 33628 23546
rect 33572 23492 33628 23494
rect 33676 23546 33732 23548
rect 33676 23494 33678 23546
rect 33678 23494 33730 23546
rect 33730 23494 33732 23546
rect 33676 23492 33732 23494
rect 33964 24668 34020 24724
rect 32732 19852 32788 19908
rect 32956 20524 33012 20580
rect 33468 21978 33524 21980
rect 33468 21926 33470 21978
rect 33470 21926 33522 21978
rect 33522 21926 33524 21978
rect 33468 21924 33524 21926
rect 33572 21978 33628 21980
rect 33572 21926 33574 21978
rect 33574 21926 33626 21978
rect 33626 21926 33628 21978
rect 33572 21924 33628 21926
rect 33676 21978 33732 21980
rect 33676 21926 33678 21978
rect 33678 21926 33730 21978
rect 33730 21926 33732 21978
rect 33676 21924 33732 21926
rect 33180 20412 33236 20468
rect 33468 20410 33524 20412
rect 33468 20358 33470 20410
rect 33470 20358 33522 20410
rect 33522 20358 33524 20410
rect 33468 20356 33524 20358
rect 33572 20410 33628 20412
rect 33572 20358 33574 20410
rect 33574 20358 33626 20410
rect 33626 20358 33628 20410
rect 33572 20356 33628 20358
rect 33676 20410 33732 20412
rect 33676 20358 33678 20410
rect 33678 20358 33730 20410
rect 33730 20358 33732 20410
rect 33676 20356 33732 20358
rect 33180 19628 33236 19684
rect 33068 19404 33124 19460
rect 33068 19180 33124 19236
rect 33852 19180 33908 19236
rect 33468 18842 33524 18844
rect 33468 18790 33470 18842
rect 33470 18790 33522 18842
rect 33522 18790 33524 18842
rect 33468 18788 33524 18790
rect 33572 18842 33628 18844
rect 33572 18790 33574 18842
rect 33574 18790 33626 18842
rect 33626 18790 33628 18842
rect 33572 18788 33628 18790
rect 33676 18842 33732 18844
rect 33676 18790 33678 18842
rect 33678 18790 33730 18842
rect 33730 18790 33732 18842
rect 33676 18788 33732 18790
rect 33292 18396 33348 18452
rect 32956 17500 33012 17556
rect 33468 17274 33524 17276
rect 33468 17222 33470 17274
rect 33470 17222 33522 17274
rect 33522 17222 33524 17274
rect 33468 17220 33524 17222
rect 33572 17274 33628 17276
rect 33572 17222 33574 17274
rect 33574 17222 33626 17274
rect 33626 17222 33628 17274
rect 33572 17220 33628 17222
rect 33676 17274 33732 17276
rect 33676 17222 33678 17274
rect 33678 17222 33730 17274
rect 33730 17222 33732 17274
rect 33676 17220 33732 17222
rect 33180 16994 33236 16996
rect 33180 16942 33182 16994
rect 33182 16942 33234 16994
rect 33234 16942 33236 16994
rect 33180 16940 33236 16942
rect 32956 16098 33012 16100
rect 32956 16046 32958 16098
rect 32958 16046 33010 16098
rect 33010 16046 33012 16098
rect 32956 16044 33012 16046
rect 31052 12962 31108 12964
rect 31052 12910 31054 12962
rect 31054 12910 31106 12962
rect 31106 12910 31108 12962
rect 31052 12908 31108 12910
rect 31276 12850 31332 12852
rect 31276 12798 31278 12850
rect 31278 12798 31330 12850
rect 31330 12798 31332 12850
rect 31276 12796 31332 12798
rect 32508 15596 32564 15652
rect 33180 15426 33236 15428
rect 33180 15374 33182 15426
rect 33182 15374 33234 15426
rect 33234 15374 33236 15426
rect 33180 15372 33236 15374
rect 32396 14028 32452 14084
rect 32396 13356 32452 13412
rect 32284 12572 32340 12628
rect 32396 12796 32452 12852
rect 32060 12124 32116 12180
rect 31836 10556 31892 10612
rect 31724 10498 31780 10500
rect 31724 10446 31726 10498
rect 31726 10446 31778 10498
rect 31778 10446 31780 10498
rect 31724 10444 31780 10446
rect 31052 10108 31108 10164
rect 31836 9436 31892 9492
rect 32508 12684 32564 12740
rect 32956 12796 33012 12852
rect 33068 14140 33124 14196
rect 32732 12684 32788 12740
rect 33468 15706 33524 15708
rect 33468 15654 33470 15706
rect 33470 15654 33522 15706
rect 33522 15654 33524 15706
rect 33468 15652 33524 15654
rect 33572 15706 33628 15708
rect 33572 15654 33574 15706
rect 33574 15654 33626 15706
rect 33626 15654 33628 15706
rect 33572 15652 33628 15654
rect 33676 15706 33732 15708
rect 33676 15654 33678 15706
rect 33678 15654 33730 15706
rect 33730 15654 33732 15706
rect 33676 15652 33732 15654
rect 33468 14138 33524 14140
rect 33468 14086 33470 14138
rect 33470 14086 33522 14138
rect 33522 14086 33524 14138
rect 33468 14084 33524 14086
rect 33572 14138 33628 14140
rect 33572 14086 33574 14138
rect 33574 14086 33626 14138
rect 33626 14086 33628 14138
rect 33572 14084 33628 14086
rect 33676 14138 33732 14140
rect 33676 14086 33678 14138
rect 33678 14086 33730 14138
rect 33730 14086 33732 14138
rect 33676 14084 33732 14086
rect 33180 12178 33236 12180
rect 33180 12126 33182 12178
rect 33182 12126 33234 12178
rect 33234 12126 33236 12178
rect 33180 12124 33236 12126
rect 32620 11394 32676 11396
rect 32620 11342 32622 11394
rect 32622 11342 32674 11394
rect 32674 11342 32676 11394
rect 32620 11340 32676 11342
rect 30940 9042 30996 9044
rect 30940 8990 30942 9042
rect 30942 8990 30994 9042
rect 30994 8990 30996 9042
rect 30940 8988 30996 8990
rect 30268 7644 30324 7700
rect 31612 8540 31668 8596
rect 31052 7698 31108 7700
rect 31052 7646 31054 7698
rect 31054 7646 31106 7698
rect 31106 7646 31108 7698
rect 31052 7644 31108 7646
rect 30492 7420 30548 7476
rect 29820 6578 29876 6580
rect 29820 6526 29822 6578
rect 29822 6526 29874 6578
rect 29874 6526 29876 6578
rect 29820 6524 29876 6526
rect 29596 6300 29652 6356
rect 31164 7362 31220 7364
rect 31164 7310 31166 7362
rect 31166 7310 31218 7362
rect 31218 7310 31220 7362
rect 31164 7308 31220 7310
rect 30604 6860 30660 6916
rect 30716 6748 30772 6804
rect 31724 8428 31780 8484
rect 31500 7308 31556 7364
rect 30044 6076 30100 6132
rect 30156 6412 30212 6468
rect 29820 6018 29876 6020
rect 29820 5966 29822 6018
rect 29822 5966 29874 6018
rect 29874 5966 29876 6018
rect 29820 5964 29876 5966
rect 30492 6076 30548 6132
rect 30380 5906 30436 5908
rect 30380 5854 30382 5906
rect 30382 5854 30434 5906
rect 30434 5854 30436 5906
rect 30380 5852 30436 5854
rect 29372 5628 29428 5684
rect 29436 5514 29492 5516
rect 29436 5462 29438 5514
rect 29438 5462 29490 5514
rect 29490 5462 29492 5514
rect 29436 5460 29492 5462
rect 29540 5514 29596 5516
rect 29540 5462 29542 5514
rect 29542 5462 29594 5514
rect 29594 5462 29596 5514
rect 29540 5460 29596 5462
rect 29644 5514 29700 5516
rect 29644 5462 29646 5514
rect 29646 5462 29698 5514
rect 29698 5462 29700 5514
rect 29644 5460 29700 5462
rect 29036 5122 29092 5124
rect 29036 5070 29038 5122
rect 29038 5070 29090 5122
rect 29090 5070 29092 5122
rect 29036 5068 29092 5070
rect 30828 5964 30884 6020
rect 32060 7868 32116 7924
rect 32732 9436 32788 9492
rect 32508 9100 32564 9156
rect 32396 8540 32452 8596
rect 32396 7868 32452 7924
rect 32508 8092 32564 8148
rect 31948 7532 32004 7588
rect 31164 6466 31220 6468
rect 31164 6414 31166 6466
rect 31166 6414 31218 6466
rect 31218 6414 31220 6466
rect 31164 6412 31220 6414
rect 30604 5740 30660 5796
rect 28588 4338 28644 4340
rect 28588 4286 28590 4338
rect 28590 4286 28642 4338
rect 28642 4286 28644 4338
rect 28588 4284 28644 4286
rect 27580 3724 27636 3780
rect 26572 3612 26628 3668
rect 27020 3554 27076 3556
rect 27020 3502 27022 3554
rect 27022 3502 27074 3554
rect 27074 3502 27076 3554
rect 27020 3500 27076 3502
rect 26348 3388 26404 3444
rect 27468 3442 27524 3444
rect 27468 3390 27470 3442
rect 27470 3390 27522 3442
rect 27522 3390 27524 3442
rect 27468 3388 27524 3390
rect 25404 3162 25460 3164
rect 25404 3110 25406 3162
rect 25406 3110 25458 3162
rect 25458 3110 25460 3162
rect 25404 3108 25460 3110
rect 25508 3162 25564 3164
rect 25508 3110 25510 3162
rect 25510 3110 25562 3162
rect 25562 3110 25564 3162
rect 25508 3108 25564 3110
rect 25612 3162 25668 3164
rect 25612 3110 25614 3162
rect 25614 3110 25666 3162
rect 25666 3110 25668 3162
rect 25612 3108 25668 3110
rect 25116 1148 25172 1204
rect 28588 3724 28644 3780
rect 30268 4172 30324 4228
rect 29436 3946 29492 3948
rect 29436 3894 29438 3946
rect 29438 3894 29490 3946
rect 29490 3894 29492 3946
rect 29436 3892 29492 3894
rect 29540 3946 29596 3948
rect 29540 3894 29542 3946
rect 29542 3894 29594 3946
rect 29594 3894 29596 3946
rect 29540 3892 29596 3894
rect 29644 3946 29700 3948
rect 29644 3894 29646 3946
rect 29646 3894 29698 3946
rect 29698 3894 29700 3946
rect 29644 3892 29700 3894
rect 28700 3388 28756 3444
rect 29148 3500 29204 3556
rect 29596 3554 29652 3556
rect 29596 3502 29598 3554
rect 29598 3502 29650 3554
rect 29650 3502 29652 3554
rect 29596 3500 29652 3502
rect 30268 3554 30324 3556
rect 30268 3502 30270 3554
rect 30270 3502 30322 3554
rect 30322 3502 30324 3554
rect 30268 3500 30324 3502
rect 29372 3442 29428 3444
rect 29372 3390 29374 3442
rect 29374 3390 29426 3442
rect 29426 3390 29428 3442
rect 29372 3388 29428 3390
rect 31948 6300 32004 6356
rect 31724 6130 31780 6132
rect 31724 6078 31726 6130
rect 31726 6078 31778 6130
rect 31778 6078 31780 6130
rect 31724 6076 31780 6078
rect 31276 4172 31332 4228
rect 30716 3612 30772 3668
rect 31948 5068 32004 5124
rect 31724 4396 31780 4452
rect 32172 7474 32228 7476
rect 32172 7422 32174 7474
rect 32174 7422 32226 7474
rect 32226 7422 32228 7474
rect 32172 7420 32228 7422
rect 32284 5682 32340 5684
rect 32284 5630 32286 5682
rect 32286 5630 32338 5682
rect 32338 5630 32340 5682
rect 32284 5628 32340 5630
rect 32396 5122 32452 5124
rect 32396 5070 32398 5122
rect 32398 5070 32450 5122
rect 32450 5070 32452 5122
rect 32396 5068 32452 5070
rect 32172 4396 32228 4452
rect 32284 3724 32340 3780
rect 33180 11506 33236 11508
rect 33180 11454 33182 11506
rect 33182 11454 33234 11506
rect 33234 11454 33236 11506
rect 33180 11452 33236 11454
rect 32956 10780 33012 10836
rect 33068 10444 33124 10500
rect 33468 12570 33524 12572
rect 33468 12518 33470 12570
rect 33470 12518 33522 12570
rect 33522 12518 33524 12570
rect 33468 12516 33524 12518
rect 33572 12570 33628 12572
rect 33572 12518 33574 12570
rect 33574 12518 33626 12570
rect 33626 12518 33628 12570
rect 33572 12516 33628 12518
rect 33676 12570 33732 12572
rect 33676 12518 33678 12570
rect 33678 12518 33730 12570
rect 33730 12518 33732 12570
rect 33676 12516 33732 12518
rect 33852 11900 33908 11956
rect 33468 11002 33524 11004
rect 33468 10950 33470 11002
rect 33470 10950 33522 11002
rect 33522 10950 33524 11002
rect 33468 10948 33524 10950
rect 33572 11002 33628 11004
rect 33572 10950 33574 11002
rect 33574 10950 33626 11002
rect 33626 10950 33628 11002
rect 33572 10948 33628 10950
rect 33676 11002 33732 11004
rect 33676 10950 33678 11002
rect 33678 10950 33730 11002
rect 33730 10950 33732 11002
rect 33676 10948 33732 10950
rect 32844 5292 32900 5348
rect 33468 9434 33524 9436
rect 33468 9382 33470 9434
rect 33470 9382 33522 9434
rect 33522 9382 33524 9434
rect 33468 9380 33524 9382
rect 33572 9434 33628 9436
rect 33572 9382 33574 9434
rect 33574 9382 33626 9434
rect 33626 9382 33628 9434
rect 33572 9380 33628 9382
rect 33676 9434 33732 9436
rect 33676 9382 33678 9434
rect 33678 9382 33730 9434
rect 33730 9382 33732 9434
rect 33676 9380 33732 9382
rect 33292 9266 33348 9268
rect 33292 9214 33294 9266
rect 33294 9214 33346 9266
rect 33346 9214 33348 9266
rect 33292 9212 33348 9214
rect 33852 8316 33908 8372
rect 33468 7866 33524 7868
rect 33468 7814 33470 7866
rect 33470 7814 33522 7866
rect 33522 7814 33524 7866
rect 33468 7812 33524 7814
rect 33572 7866 33628 7868
rect 33572 7814 33574 7866
rect 33574 7814 33626 7866
rect 33626 7814 33628 7866
rect 33572 7812 33628 7814
rect 33676 7866 33732 7868
rect 33676 7814 33678 7866
rect 33678 7814 33730 7866
rect 33730 7814 33732 7866
rect 33676 7812 33732 7814
rect 33180 7420 33236 7476
rect 33852 7420 33908 7476
rect 33468 6298 33524 6300
rect 33068 6188 33124 6244
rect 33468 6246 33470 6298
rect 33470 6246 33522 6298
rect 33522 6246 33524 6298
rect 33468 6244 33524 6246
rect 33572 6298 33628 6300
rect 33572 6246 33574 6298
rect 33574 6246 33626 6298
rect 33626 6246 33628 6298
rect 33572 6244 33628 6246
rect 33676 6298 33732 6300
rect 33676 6246 33678 6298
rect 33678 6246 33730 6298
rect 33730 6246 33732 6298
rect 33676 6244 33732 6246
rect 33180 5794 33236 5796
rect 33180 5742 33182 5794
rect 33182 5742 33234 5794
rect 33234 5742 33236 5794
rect 33180 5740 33236 5742
rect 33468 4730 33524 4732
rect 33468 4678 33470 4730
rect 33470 4678 33522 4730
rect 33522 4678 33524 4730
rect 33468 4676 33524 4678
rect 33572 4730 33628 4732
rect 33572 4678 33574 4730
rect 33574 4678 33626 4730
rect 33626 4678 33628 4730
rect 33572 4676 33628 4678
rect 33676 4730 33732 4732
rect 33676 4678 33678 4730
rect 33678 4678 33730 4730
rect 33730 4678 33732 4730
rect 33676 4676 33732 4678
rect 33180 4226 33236 4228
rect 33180 4174 33182 4226
rect 33182 4174 33234 4226
rect 33234 4174 33236 4226
rect 33180 4172 33236 4174
rect 33180 3948 33236 4004
rect 33852 3500 33908 3556
rect 33468 3162 33524 3164
rect 33468 3110 33470 3162
rect 33470 3110 33522 3162
rect 33522 3110 33524 3162
rect 33468 3108 33524 3110
rect 33572 3162 33628 3164
rect 33572 3110 33574 3162
rect 33574 3110 33626 3162
rect 33626 3110 33628 3162
rect 33572 3108 33628 3110
rect 33676 3162 33732 3164
rect 33676 3110 33678 3162
rect 33678 3110 33730 3162
rect 33730 3110 33732 3162
rect 33676 3108 33732 3110
<< metal3 >>
rect 34200 33460 35000 33488
rect 23874 33404 23884 33460
rect 23940 33404 35000 33460
rect 34200 33376 35000 33404
rect 20626 33068 20636 33124
rect 20692 33068 27468 33124
rect 27524 33068 27534 33124
rect 8754 32060 8764 32116
rect 8820 32060 20748 32116
rect 20804 32060 20814 32116
rect 19618 31948 19628 32004
rect 19684 31948 28924 32004
rect 28980 31948 28990 32004
rect 4946 31836 4956 31892
rect 5012 31836 6076 31892
rect 6132 31836 6142 31892
rect 7970 31836 7980 31892
rect 8036 31836 9436 31892
rect 9492 31836 9502 31892
rect 6850 31724 6860 31780
rect 6916 31724 26236 31780
rect 26292 31724 26302 31780
rect 10434 31612 10444 31668
rect 10500 31612 23884 31668
rect 23940 31612 23950 31668
rect 5058 31500 5068 31556
rect 5124 31500 19628 31556
rect 19684 31500 19694 31556
rect 9266 31332 9276 31388
rect 9332 31332 9380 31388
rect 9436 31332 9484 31388
rect 9540 31332 9550 31388
rect 17330 31332 17340 31388
rect 17396 31332 17444 31388
rect 17500 31332 17548 31388
rect 17604 31332 17614 31388
rect 25394 31332 25404 31388
rect 25460 31332 25508 31388
rect 25564 31332 25612 31388
rect 25668 31332 25678 31388
rect 33458 31332 33468 31388
rect 33524 31332 33572 31388
rect 33628 31332 33676 31388
rect 33732 31332 33742 31388
rect 20850 31276 20860 31332
rect 20916 31276 24556 31332
rect 24612 31276 24622 31332
rect 5842 31164 5852 31220
rect 5908 31164 7196 31220
rect 7252 31164 7262 31220
rect 19506 31164 19516 31220
rect 19572 31164 21756 31220
rect 21812 31164 21822 31220
rect 22866 31164 22876 31220
rect 22932 31164 26236 31220
rect 26292 31164 26302 31220
rect 28690 31164 28700 31220
rect 28756 31164 33236 31220
rect 3714 31052 3724 31108
rect 3780 31052 20972 31108
rect 21028 31052 21038 31108
rect 23650 31052 23660 31108
rect 23716 31052 23726 31108
rect 24882 31052 24892 31108
rect 24948 31052 25228 31108
rect 25284 31052 25294 31108
rect 29138 31052 29148 31108
rect 29204 31052 30492 31108
rect 30548 31052 30558 31108
rect 12226 30940 12236 30996
rect 12292 30940 13804 30996
rect 13860 30940 13870 30996
rect 18610 30940 18620 30996
rect 18676 30940 20748 30996
rect 20804 30940 20814 30996
rect 23660 30884 23716 31052
rect 29250 30940 29260 30996
rect 29316 30940 32732 30996
rect 32788 30940 32798 30996
rect 13346 30828 13356 30884
rect 13412 30828 23716 30884
rect 24332 30828 32172 30884
rect 32228 30828 32238 30884
rect 24332 30772 24388 30828
rect 33180 30772 33236 31164
rect 34200 30772 35000 30800
rect 13458 30716 13468 30772
rect 13524 30716 15260 30772
rect 15316 30716 15326 30772
rect 21858 30716 21868 30772
rect 21924 30716 24388 30772
rect 25218 30716 25228 30772
rect 25284 30716 32956 30772
rect 33012 30716 33022 30772
rect 33180 30716 35000 30772
rect 34200 30688 35000 30716
rect 5234 30548 5244 30604
rect 5300 30548 5348 30604
rect 5404 30548 5452 30604
rect 5508 30548 5518 30604
rect 13298 30548 13308 30604
rect 13364 30548 13412 30604
rect 13468 30548 13516 30604
rect 13572 30548 13582 30604
rect 21362 30548 21372 30604
rect 21428 30548 21476 30604
rect 21532 30548 21580 30604
rect 21636 30548 21646 30604
rect 29426 30548 29436 30604
rect 29492 30548 29540 30604
rect 29596 30548 29644 30604
rect 29700 30548 29710 30604
rect 14802 30492 14812 30548
rect 14868 30492 15372 30548
rect 15428 30492 15438 30548
rect 22764 30492 28700 30548
rect 28756 30492 28766 30548
rect 22764 30436 22820 30492
rect 14018 30380 14028 30436
rect 14084 30380 16492 30436
rect 16548 30380 16558 30436
rect 20402 30380 20412 30436
rect 20468 30380 22820 30436
rect 23426 30380 23436 30436
rect 23492 30380 32844 30436
rect 32900 30380 32910 30436
rect 7186 30268 7196 30324
rect 7252 30268 20076 30324
rect 20132 30268 20142 30324
rect 20626 30268 20636 30324
rect 20692 30268 31052 30324
rect 31108 30268 31118 30324
rect 31266 30268 31276 30324
rect 31332 30268 32172 30324
rect 32228 30268 32238 30324
rect 14886 30156 14924 30212
rect 14980 30156 14990 30212
rect 17826 30156 17836 30212
rect 17892 30156 18508 30212
rect 18564 30156 20300 30212
rect 20356 30156 23436 30212
rect 23492 30156 23502 30212
rect 24322 30156 24332 30212
rect 24388 30156 25340 30212
rect 25396 30156 25406 30212
rect 26562 30156 26572 30212
rect 26628 30156 28364 30212
rect 28420 30156 29596 30212
rect 29652 30156 30268 30212
rect 30324 30156 30334 30212
rect 2930 30044 2940 30100
rect 2996 30044 3948 30100
rect 4004 30044 4014 30100
rect 6402 30044 6412 30100
rect 6468 30044 7644 30100
rect 7700 30044 7710 30100
rect 12338 30044 12348 30100
rect 12404 30044 15036 30100
rect 15092 30044 15102 30100
rect 18722 30044 18732 30100
rect 18788 30044 25564 30100
rect 25620 30044 25630 30100
rect 28466 30044 28476 30100
rect 28532 30044 30604 30100
rect 30660 30044 30670 30100
rect 8306 29932 8316 29988
rect 8372 29932 8876 29988
rect 8932 29932 8942 29988
rect 9426 29932 9436 29988
rect 9492 29932 12684 29988
rect 12740 29932 12750 29988
rect 16930 29932 16940 29988
rect 16996 29932 17276 29988
rect 17332 29932 17342 29988
rect 20066 29932 20076 29988
rect 20132 29932 24332 29988
rect 24388 29932 24398 29988
rect 9266 29764 9276 29820
rect 9332 29764 9380 29820
rect 9436 29764 9484 29820
rect 9540 29764 9550 29820
rect 17330 29764 17340 29820
rect 17396 29764 17444 29820
rect 17500 29764 17548 29820
rect 17604 29764 17614 29820
rect 25394 29764 25404 29820
rect 25460 29764 25508 29820
rect 25564 29764 25612 29820
rect 25668 29764 25678 29820
rect 33458 29764 33468 29820
rect 33524 29764 33572 29820
rect 33628 29764 33676 29820
rect 33732 29764 33742 29820
rect 17724 29708 22316 29764
rect 22372 29708 24948 29764
rect 17724 29652 17780 29708
rect 24892 29652 24948 29708
rect 5506 29596 5516 29652
rect 5572 29596 6860 29652
rect 6916 29596 6926 29652
rect 9090 29596 9100 29652
rect 9156 29596 11676 29652
rect 11732 29596 15932 29652
rect 15988 29596 15998 29652
rect 16482 29596 16492 29652
rect 16548 29596 17780 29652
rect 18386 29596 18396 29652
rect 18452 29596 24108 29652
rect 24164 29596 24668 29652
rect 24724 29596 24734 29652
rect 24892 29596 31388 29652
rect 31444 29596 32508 29652
rect 32564 29596 32574 29652
rect 6626 29484 6636 29540
rect 6692 29484 8652 29540
rect 8708 29484 8718 29540
rect 9650 29484 9660 29540
rect 9716 29484 10556 29540
rect 10612 29484 10622 29540
rect 14998 29484 15036 29540
rect 15092 29484 15102 29540
rect 15698 29484 15708 29540
rect 15764 29484 18620 29540
rect 18676 29484 18686 29540
rect 22876 29484 30380 29540
rect 30436 29484 30446 29540
rect 22876 29428 22932 29484
rect 7746 29372 7756 29428
rect 7812 29372 8540 29428
rect 8596 29372 10332 29428
rect 10388 29372 10398 29428
rect 10556 29372 12124 29428
rect 12180 29372 12190 29428
rect 12562 29372 12572 29428
rect 12628 29372 14364 29428
rect 14420 29372 16156 29428
rect 16212 29372 16222 29428
rect 18834 29372 18844 29428
rect 18900 29372 20972 29428
rect 21028 29372 21308 29428
rect 21364 29372 22652 29428
rect 22708 29372 22718 29428
rect 22866 29372 22876 29428
rect 22932 29372 22942 29428
rect 26226 29372 26236 29428
rect 26292 29372 31948 29428
rect 32004 29372 32014 29428
rect 10556 29316 10612 29372
rect 1698 29260 1708 29316
rect 1764 29260 2268 29316
rect 2324 29260 4508 29316
rect 4564 29260 4574 29316
rect 5282 29260 5292 29316
rect 5348 29260 6524 29316
rect 6580 29260 6590 29316
rect 6738 29260 6748 29316
rect 6804 29260 9324 29316
rect 9380 29260 9660 29316
rect 9716 29260 10612 29316
rect 10882 29260 10892 29316
rect 10948 29260 15148 29316
rect 17826 29260 17836 29316
rect 17892 29260 19516 29316
rect 19572 29260 19582 29316
rect 20514 29260 20524 29316
rect 20580 29260 22988 29316
rect 23044 29260 24780 29316
rect 24836 29260 33180 29316
rect 33236 29260 33246 29316
rect 15092 29204 15148 29260
rect 4620 29148 5852 29204
rect 5908 29148 14140 29204
rect 14196 29148 14206 29204
rect 15092 29148 15708 29204
rect 15764 29148 15774 29204
rect 18274 29148 18284 29204
rect 18340 29148 23436 29204
rect 23492 29148 23502 29204
rect 24882 29148 24892 29204
rect 24948 29148 25228 29204
rect 25284 29148 25294 29204
rect 26338 29148 26348 29204
rect 26404 29148 29876 29204
rect 4620 29092 4676 29148
rect 25228 29092 25284 29148
rect 29820 29092 29876 29148
rect 4610 29036 4620 29092
rect 4676 29036 4686 29092
rect 9090 29036 9100 29092
rect 9156 29036 9772 29092
rect 9828 29036 9838 29092
rect 13692 29036 16044 29092
rect 16100 29036 16492 29092
rect 16548 29036 16558 29092
rect 17378 29036 17388 29092
rect 17444 29036 20076 29092
rect 20132 29036 20142 29092
rect 25228 29036 26572 29092
rect 26628 29036 26638 29092
rect 29810 29036 29820 29092
rect 29876 29036 32396 29092
rect 32452 29036 32462 29092
rect 5234 28980 5244 29036
rect 5300 28980 5348 29036
rect 5404 28980 5452 29036
rect 5508 28980 5518 29036
rect 13298 28980 13308 29036
rect 13364 28980 13412 29036
rect 13468 28980 13516 29036
rect 13572 28980 13582 29036
rect 6514 28924 6524 28980
rect 6580 28924 8092 28980
rect 8148 28924 12796 28980
rect 12852 28924 12862 28980
rect 13692 28868 13748 29036
rect 21362 28980 21372 29036
rect 21428 28980 21476 29036
rect 21532 28980 21580 29036
rect 21636 28980 21646 29036
rect 29426 28980 29436 29036
rect 29492 28980 29540 29036
rect 29596 28980 29644 29036
rect 29700 28980 29710 29036
rect 4834 28812 4844 28868
rect 4900 28812 6636 28868
rect 6692 28812 6702 28868
rect 9202 28812 9212 28868
rect 9268 28812 13748 28868
rect 13804 28924 17724 28980
rect 17780 28924 17790 28980
rect 29820 28924 33068 28980
rect 33124 28924 33134 28980
rect 13804 28756 13860 28924
rect 29820 28868 29876 28924
rect 14690 28812 14700 28868
rect 14756 28812 15820 28868
rect 15876 28812 15886 28868
rect 20850 28812 20860 28868
rect 20916 28812 20972 28868
rect 21028 28812 21308 28868
rect 21364 28812 21374 28868
rect 23986 28812 23996 28868
rect 24052 28812 26908 28868
rect 26964 28812 26974 28868
rect 29586 28812 29596 28868
rect 29652 28812 29876 28868
rect 31266 28812 31276 28868
rect 31332 28812 32284 28868
rect 32340 28812 32350 28868
rect 4050 28700 4060 28756
rect 4116 28700 6076 28756
rect 6132 28700 6142 28756
rect 10994 28700 11004 28756
rect 11060 28700 12908 28756
rect 12964 28700 13468 28756
rect 13524 28700 13860 28756
rect 15026 28700 15036 28756
rect 15092 28700 17948 28756
rect 18004 28700 18284 28756
rect 18340 28700 18350 28756
rect 19292 28700 19964 28756
rect 20020 28700 20030 28756
rect 20402 28700 20412 28756
rect 20468 28700 21644 28756
rect 21700 28700 21710 28756
rect 24658 28700 24668 28756
rect 24724 28700 25564 28756
rect 25620 28700 25630 28756
rect 29138 28700 29148 28756
rect 29204 28700 33180 28756
rect 33236 28700 33246 28756
rect 19292 28644 19348 28700
rect 5170 28588 5180 28644
rect 5236 28588 6300 28644
rect 6356 28588 6366 28644
rect 11554 28588 11564 28644
rect 11620 28588 12124 28644
rect 12180 28588 15484 28644
rect 15540 28588 15550 28644
rect 18386 28588 18396 28644
rect 18452 28588 19292 28644
rect 19348 28588 19358 28644
rect 19618 28588 19628 28644
rect 19684 28588 20300 28644
rect 20356 28588 20366 28644
rect 24546 28588 24556 28644
rect 24612 28588 27692 28644
rect 27748 28588 28588 28644
rect 28644 28588 28654 28644
rect 31266 28588 31276 28644
rect 31332 28588 34076 28644
rect 34132 28588 34142 28644
rect 9986 28476 9996 28532
rect 10052 28476 10892 28532
rect 10948 28476 10958 28532
rect 13122 28476 13132 28532
rect 13188 28476 14028 28532
rect 14084 28476 14094 28532
rect 15026 28476 15036 28532
rect 15092 28476 16828 28532
rect 16884 28476 16894 28532
rect 18834 28476 18844 28532
rect 18900 28476 20468 28532
rect 20626 28476 20636 28532
rect 20692 28476 20860 28532
rect 20916 28476 20926 28532
rect 21074 28476 21084 28532
rect 21140 28476 21644 28532
rect 21700 28476 21710 28532
rect 21858 28476 21868 28532
rect 21924 28476 26460 28532
rect 26516 28476 26526 28532
rect 29026 28476 29036 28532
rect 29092 28476 29372 28532
rect 29428 28476 29438 28532
rect 30146 28476 30156 28532
rect 30212 28476 30828 28532
rect 30884 28476 30894 28532
rect 7858 28364 7868 28420
rect 7924 28364 9772 28420
rect 9828 28364 10220 28420
rect 10276 28364 10332 28420
rect 10388 28364 10398 28420
rect 13570 28364 13580 28420
rect 13636 28364 14196 28420
rect 17490 28364 17500 28420
rect 17556 28364 18620 28420
rect 18676 28364 19404 28420
rect 19460 28364 19470 28420
rect 14140 28308 14196 28364
rect 20412 28308 20468 28476
rect 21186 28364 21196 28420
rect 21252 28364 22316 28420
rect 22372 28364 22382 28420
rect 25666 28364 25676 28420
rect 25732 28364 26348 28420
rect 26404 28364 26796 28420
rect 26852 28364 26862 28420
rect 27570 28364 27580 28420
rect 27636 28364 30380 28420
rect 30436 28364 30446 28420
rect 10770 28252 10780 28308
rect 10836 28252 12236 28308
rect 12292 28252 13692 28308
rect 13748 28252 13758 28308
rect 14140 28252 15148 28308
rect 18498 28252 18508 28308
rect 18564 28252 18574 28308
rect 20412 28252 24332 28308
rect 24388 28252 24398 28308
rect 25778 28252 25788 28308
rect 25844 28252 26124 28308
rect 26180 28252 26190 28308
rect 29474 28252 29484 28308
rect 29540 28252 30156 28308
rect 30212 28252 30222 28308
rect 9266 28196 9276 28252
rect 9332 28196 9380 28252
rect 9436 28196 9484 28252
rect 9540 28196 9550 28252
rect 9650 28140 9660 28196
rect 9716 28140 13804 28196
rect 13860 28140 13870 28196
rect 6290 28028 6300 28084
rect 6356 28028 8092 28084
rect 8148 28028 8540 28084
rect 8596 28028 8606 28084
rect 15092 28028 15148 28252
rect 17330 28196 17340 28252
rect 17396 28196 17444 28252
rect 17500 28196 17548 28252
rect 17604 28196 17614 28252
rect 18508 28196 18564 28252
rect 25394 28196 25404 28252
rect 25460 28196 25508 28252
rect 25564 28196 25612 28252
rect 25668 28196 25678 28252
rect 33458 28196 33468 28252
rect 33524 28196 33572 28252
rect 33628 28196 33676 28252
rect 33732 28196 33742 28252
rect 18508 28140 22540 28196
rect 22596 28140 22606 28196
rect 26898 28140 26908 28196
rect 26964 28140 30604 28196
rect 30660 28140 30670 28196
rect 34200 28084 35000 28112
rect 15204 28028 15214 28084
rect 17266 28028 17276 28084
rect 17332 28028 18508 28084
rect 18564 28028 18574 28084
rect 20514 28028 20524 28084
rect 20580 28028 25788 28084
rect 25844 28028 25854 28084
rect 30258 28028 30268 28084
rect 30324 28028 35000 28084
rect 34200 28000 35000 28028
rect 7746 27916 7756 27972
rect 7812 27916 8764 27972
rect 8820 27916 9212 27972
rect 9268 27916 9278 27972
rect 9538 27916 9548 27972
rect 9604 27916 10780 27972
rect 10836 27916 10846 27972
rect 13682 27916 13692 27972
rect 13748 27916 25452 27972
rect 25508 27916 25518 27972
rect 26450 27916 26460 27972
rect 26516 27916 29484 27972
rect 29540 27916 29550 27972
rect 6290 27804 6300 27860
rect 6356 27804 6636 27860
rect 6692 27804 6702 27860
rect 11778 27804 11788 27860
rect 11844 27804 13132 27860
rect 13188 27804 17052 27860
rect 17108 27804 20412 27860
rect 20468 27804 20478 27860
rect 20850 27804 20860 27860
rect 20916 27804 23996 27860
rect 24052 27804 25900 27860
rect 25956 27804 25966 27860
rect 26898 27804 26908 27860
rect 26964 27804 28140 27860
rect 28196 27804 28206 27860
rect 6738 27692 6748 27748
rect 6804 27692 8988 27748
rect 9044 27692 11508 27748
rect 18946 27692 18956 27748
rect 19012 27692 21756 27748
rect 21812 27692 21822 27748
rect 22530 27692 22540 27748
rect 22596 27692 28476 27748
rect 28532 27692 28542 27748
rect 11452 27636 11508 27692
rect 4610 27580 4620 27636
rect 4676 27580 7812 27636
rect 8642 27580 8652 27636
rect 8708 27580 9772 27636
rect 9828 27580 9838 27636
rect 11442 27580 11452 27636
rect 11508 27580 12348 27636
rect 12404 27580 12414 27636
rect 19170 27580 19180 27636
rect 19236 27580 20524 27636
rect 20580 27580 20590 27636
rect 28242 27580 28252 27636
rect 28308 27580 33180 27636
rect 33236 27580 33246 27636
rect 7756 27524 7812 27580
rect 6178 27468 6188 27524
rect 6244 27468 6748 27524
rect 6804 27468 6814 27524
rect 7746 27468 7756 27524
rect 7812 27468 11228 27524
rect 11284 27468 11294 27524
rect 25106 27468 25116 27524
rect 25172 27468 26908 27524
rect 26964 27468 26974 27524
rect 5234 27412 5244 27468
rect 5300 27412 5348 27468
rect 5404 27412 5452 27468
rect 5508 27412 5518 27468
rect 13298 27412 13308 27468
rect 13364 27412 13412 27468
rect 13468 27412 13516 27468
rect 13572 27412 13582 27468
rect 21362 27412 21372 27468
rect 21428 27412 21476 27468
rect 21532 27412 21580 27468
rect 21636 27412 21646 27468
rect 29426 27412 29436 27468
rect 29492 27412 29540 27468
rect 29596 27412 29644 27468
rect 29700 27412 29710 27468
rect 8418 27356 8428 27412
rect 8484 27356 9660 27412
rect 9716 27356 9726 27412
rect 14102 27356 14140 27412
rect 14196 27356 14206 27412
rect 14774 27356 14812 27412
rect 14868 27356 14878 27412
rect 24994 27356 25004 27412
rect 25060 27356 28364 27412
rect 28420 27356 28430 27412
rect 8530 27244 8540 27300
rect 8596 27244 12012 27300
rect 12068 27244 12078 27300
rect 12898 27244 12908 27300
rect 12964 27244 14252 27300
rect 14308 27244 14318 27300
rect 18722 27244 18732 27300
rect 18788 27244 20188 27300
rect 20244 27244 20254 27300
rect 22194 27244 22204 27300
rect 22260 27244 33068 27300
rect 33124 27244 33134 27300
rect 2930 27132 2940 27188
rect 2996 27132 7980 27188
rect 8036 27132 8046 27188
rect 9090 27132 9100 27188
rect 9156 27132 22428 27188
rect 22484 27132 23436 27188
rect 23492 27132 23502 27188
rect 7074 27020 7084 27076
rect 7140 27020 8204 27076
rect 8260 27020 8270 27076
rect 8866 27020 8876 27076
rect 8932 27020 8942 27076
rect 14242 27020 14252 27076
rect 14308 27020 14318 27076
rect 17042 27020 17052 27076
rect 17108 27020 19292 27076
rect 19348 27020 19358 27076
rect 20514 27020 20524 27076
rect 20580 27020 20860 27076
rect 20916 27020 20926 27076
rect 27346 27020 27356 27076
rect 27412 27020 29596 27076
rect 29652 27020 29662 27076
rect 5954 26908 5964 26964
rect 6020 26908 6972 26964
rect 7028 26908 7038 26964
rect 7158 26908 7196 26964
rect 7252 26908 7262 26964
rect 7298 26796 7308 26852
rect 7364 26796 7980 26852
rect 8036 26796 8046 26852
rect 6626 26684 6636 26740
rect 6692 26684 8540 26740
rect 8596 26684 8606 26740
rect 4946 26572 4956 26628
rect 5012 26572 7308 26628
rect 7364 26572 7374 26628
rect 8876 26516 8932 27020
rect 14252 26964 14308 27020
rect 9762 26908 9772 26964
rect 9828 26908 10668 26964
rect 10724 26908 10734 26964
rect 10892 26908 11228 26964
rect 11284 26908 11294 26964
rect 11890 26908 11900 26964
rect 11956 26908 12460 26964
rect 12516 26908 12572 26964
rect 12628 26908 13468 26964
rect 13524 26908 13534 26964
rect 14252 26908 14812 26964
rect 14868 26908 15820 26964
rect 15876 26908 15886 26964
rect 20402 26908 20412 26964
rect 20468 26908 24108 26964
rect 24164 26908 25228 26964
rect 25284 26908 25294 26964
rect 27794 26908 27804 26964
rect 27860 26908 29260 26964
rect 29316 26908 29326 26964
rect 10892 26852 10948 26908
rect 9986 26796 9996 26852
rect 10052 26796 10948 26852
rect 11106 26796 11116 26852
rect 11172 26796 14420 26852
rect 14690 26796 14700 26852
rect 14756 26796 15988 26852
rect 14364 26740 14420 26796
rect 15932 26740 15988 26796
rect 16156 26796 25844 26852
rect 10294 26684 10332 26740
rect 10388 26684 10398 26740
rect 12114 26684 12124 26740
rect 12180 26684 14140 26740
rect 14196 26684 14206 26740
rect 14364 26684 14812 26740
rect 14868 26684 14878 26740
rect 15922 26684 15932 26740
rect 15988 26684 15998 26740
rect 9266 26628 9276 26684
rect 9332 26628 9380 26684
rect 9436 26628 9484 26684
rect 9540 26628 9550 26684
rect 16156 26628 16212 26796
rect 25788 26740 25844 26796
rect 21074 26684 21084 26740
rect 21140 26684 21644 26740
rect 21700 26684 21710 26740
rect 25778 26684 25788 26740
rect 25844 26684 25854 26740
rect 28242 26684 28252 26740
rect 28308 26684 29372 26740
rect 29428 26684 29438 26740
rect 17330 26628 17340 26684
rect 17396 26628 17444 26684
rect 17500 26628 17548 26684
rect 17604 26628 17614 26684
rect 25394 26628 25404 26684
rect 25460 26628 25508 26684
rect 25564 26628 25612 26684
rect 25668 26628 25678 26684
rect 33458 26628 33468 26684
rect 33524 26628 33572 26684
rect 33628 26628 33676 26684
rect 33732 26628 33742 26684
rect 13794 26572 13804 26628
rect 13860 26572 14812 26628
rect 14868 26572 16212 26628
rect 18498 26572 18508 26628
rect 18564 26572 18844 26628
rect 18900 26572 18910 26628
rect 20934 26572 20972 26628
rect 21028 26572 21038 26628
rect 29474 26572 29484 26628
rect 29540 26572 29820 26628
rect 29876 26572 29886 26628
rect 6402 26460 6412 26516
rect 6468 26460 6748 26516
rect 6804 26460 6814 26516
rect 7858 26460 7868 26516
rect 7924 26460 8372 26516
rect 8876 26460 12572 26516
rect 12628 26460 12638 26516
rect 15222 26460 15260 26516
rect 15316 26460 15326 26516
rect 17042 26460 17052 26516
rect 17108 26460 17724 26516
rect 17780 26460 18732 26516
rect 18788 26460 19740 26516
rect 19796 26460 19806 26516
rect 19954 26460 19964 26516
rect 20020 26460 22092 26516
rect 22148 26460 22158 26516
rect 8316 26404 8372 26460
rect 5058 26348 5068 26404
rect 5124 26348 7196 26404
rect 7252 26348 7420 26404
rect 7476 26348 8092 26404
rect 8148 26348 8158 26404
rect 8316 26348 9772 26404
rect 9828 26348 17388 26404
rect 17444 26348 18508 26404
rect 18564 26348 18574 26404
rect 19282 26348 19292 26404
rect 19348 26348 19628 26404
rect 19684 26348 19694 26404
rect 23090 26348 23100 26404
rect 23156 26348 29148 26404
rect 29204 26348 29214 26404
rect 4946 26236 4956 26292
rect 5012 26236 6748 26292
rect 6804 26236 6814 26292
rect 8978 26236 8988 26292
rect 9044 26236 9212 26292
rect 9268 26236 9278 26292
rect 9986 26236 9996 26292
rect 10052 26236 12572 26292
rect 12628 26236 14028 26292
rect 14084 26236 18172 26292
rect 18228 26236 18238 26292
rect 18722 26236 18732 26292
rect 18788 26236 20748 26292
rect 20804 26236 20814 26292
rect 23986 26236 23996 26292
rect 24052 26236 25340 26292
rect 25396 26236 25406 26292
rect 28998 26236 29036 26292
rect 29092 26236 29102 26292
rect 5506 26124 5516 26180
rect 5572 26124 6300 26180
rect 6356 26124 6366 26180
rect 7970 26124 7980 26180
rect 8036 26124 10668 26180
rect 10724 26124 12348 26180
rect 12404 26124 12414 26180
rect 16118 26124 16156 26180
rect 16212 26124 16222 26180
rect 16594 26124 16604 26180
rect 16660 26124 18620 26180
rect 18676 26124 19180 26180
rect 19236 26124 19246 26180
rect 19618 26124 19628 26180
rect 19684 26124 20412 26180
rect 20468 26124 20478 26180
rect 21858 26124 21868 26180
rect 21924 26124 22204 26180
rect 22260 26124 22596 26180
rect 23426 26124 23436 26180
rect 23492 26124 33180 26180
rect 33236 26124 33852 26180
rect 33908 26124 33918 26180
rect 22540 26068 22596 26124
rect 3378 26012 3388 26068
rect 3444 26012 6188 26068
rect 6244 26012 6254 26068
rect 6738 26012 6748 26068
rect 6804 26012 7868 26068
rect 7924 26012 7934 26068
rect 9874 26012 9884 26068
rect 9940 26012 10892 26068
rect 10948 26012 10958 26068
rect 11890 26012 11900 26068
rect 11956 26012 12236 26068
rect 12292 26012 12302 26068
rect 15362 26012 15372 26068
rect 15428 26012 17500 26068
rect 17556 26012 17566 26068
rect 18050 26012 18060 26068
rect 18116 26012 22316 26068
rect 22372 26012 22382 26068
rect 22540 26012 29036 26068
rect 29092 26012 29102 26068
rect 29474 26012 29484 26068
rect 29540 26012 31052 26068
rect 31108 26012 31118 26068
rect 11900 25956 11956 26012
rect 6290 25900 6300 25956
rect 6356 25900 11956 25956
rect 15138 25900 15148 25956
rect 15204 25900 16156 25956
rect 16212 25900 16940 25956
rect 16996 25900 17006 25956
rect 26908 25900 27132 25956
rect 27188 25900 27198 25956
rect 5234 25844 5244 25900
rect 5300 25844 5348 25900
rect 5404 25844 5452 25900
rect 5508 25844 5518 25900
rect 13298 25844 13308 25900
rect 13364 25844 13412 25900
rect 13468 25844 13516 25900
rect 13572 25844 13582 25900
rect 21362 25844 21372 25900
rect 21428 25844 21476 25900
rect 21532 25844 21580 25900
rect 21636 25844 21646 25900
rect 6038 25788 6076 25844
rect 6132 25788 6142 25844
rect 6514 25788 6524 25844
rect 6580 25788 10276 25844
rect 12646 25788 12684 25844
rect 12740 25788 12750 25844
rect 13906 25788 13916 25844
rect 13972 25788 15372 25844
rect 15428 25788 20524 25844
rect 20580 25788 20590 25844
rect 10220 25732 10276 25788
rect 26908 25732 26964 25900
rect 29426 25844 29436 25900
rect 29492 25844 29540 25900
rect 29596 25844 29644 25900
rect 29700 25844 29710 25900
rect 4722 25676 4732 25732
rect 4788 25676 5068 25732
rect 5124 25676 8428 25732
rect 8484 25676 8494 25732
rect 8866 25676 8876 25732
rect 8932 25676 9996 25732
rect 10052 25676 10062 25732
rect 10220 25676 14140 25732
rect 14196 25676 14206 25732
rect 14578 25676 14588 25732
rect 14644 25676 15932 25732
rect 15988 25676 15998 25732
rect 22082 25676 22092 25732
rect 22148 25676 26572 25732
rect 26628 25676 26964 25732
rect 27132 25788 29036 25844
rect 29092 25788 29102 25844
rect 29250 25788 29260 25844
rect 29316 25788 29326 25844
rect 27132 25620 27188 25788
rect 29260 25732 29316 25788
rect 27346 25676 27356 25732
rect 27412 25676 28700 25732
rect 28756 25676 28766 25732
rect 29036 25676 29316 25732
rect 29036 25620 29092 25676
rect 9202 25564 9212 25620
rect 9268 25564 10444 25620
rect 10500 25564 10510 25620
rect 12674 25564 12684 25620
rect 12740 25564 15148 25620
rect 15250 25564 15260 25620
rect 15316 25564 15708 25620
rect 15764 25564 15774 25620
rect 17714 25564 17724 25620
rect 17780 25564 18956 25620
rect 19012 25564 19022 25620
rect 19516 25564 20524 25620
rect 20580 25564 24444 25620
rect 24500 25564 27188 25620
rect 28700 25564 29092 25620
rect 29250 25564 29260 25620
rect 29316 25564 33180 25620
rect 33236 25564 33246 25620
rect 15092 25508 15148 25564
rect 19516 25508 19572 25564
rect 28700 25508 28756 25564
rect 7074 25452 7084 25508
rect 7140 25452 7150 25508
rect 10546 25452 10556 25508
rect 10612 25452 11340 25508
rect 11396 25452 11406 25508
rect 12450 25452 12460 25508
rect 12516 25452 14252 25508
rect 14308 25452 14318 25508
rect 15092 25452 16212 25508
rect 16370 25452 16380 25508
rect 16436 25452 17836 25508
rect 17892 25452 17902 25508
rect 18498 25452 18508 25508
rect 18564 25452 19572 25508
rect 19730 25452 19740 25508
rect 19796 25452 20300 25508
rect 20356 25452 20366 25508
rect 26114 25452 26124 25508
rect 26180 25452 27244 25508
rect 27300 25452 27310 25508
rect 27468 25452 28700 25508
rect 28756 25452 28766 25508
rect 29026 25452 29036 25508
rect 29092 25452 30044 25508
rect 30100 25452 30110 25508
rect 7084 25284 7140 25452
rect 16156 25396 16212 25452
rect 27468 25396 27524 25452
rect 34200 25396 35000 25424
rect 9650 25340 9660 25396
rect 9716 25340 11676 25396
rect 11732 25340 11742 25396
rect 11900 25340 12964 25396
rect 14578 25340 14588 25396
rect 14644 25340 15036 25396
rect 15092 25340 15102 25396
rect 16156 25340 16828 25396
rect 16884 25340 16894 25396
rect 18274 25340 18284 25396
rect 18340 25340 20636 25396
rect 20692 25340 23996 25396
rect 24052 25340 24062 25396
rect 24658 25340 24668 25396
rect 24724 25340 27020 25396
rect 27076 25340 27524 25396
rect 28140 25340 28588 25396
rect 28644 25340 28654 25396
rect 28914 25340 28924 25396
rect 28980 25340 35000 25396
rect 11900 25284 11956 25340
rect 2482 25228 2492 25284
rect 2548 25228 4060 25284
rect 4116 25228 4126 25284
rect 6038 25228 6076 25284
rect 6132 25228 6142 25284
rect 6290 25228 6300 25284
rect 6356 25228 6394 25284
rect 7084 25228 9548 25284
rect 9604 25228 9716 25284
rect 9986 25228 9996 25284
rect 10052 25228 11956 25284
rect 12908 25284 12964 25340
rect 28140 25284 28196 25340
rect 34200 25312 35000 25340
rect 12908 25228 18844 25284
rect 18900 25228 18910 25284
rect 19170 25228 19180 25284
rect 19236 25228 19348 25284
rect 21186 25228 21196 25284
rect 21252 25228 21980 25284
rect 22036 25228 22046 25284
rect 25218 25228 25228 25284
rect 25284 25228 27580 25284
rect 27636 25228 27646 25284
rect 28130 25228 28140 25284
rect 28196 25228 28206 25284
rect 28326 25228 28364 25284
rect 28420 25228 28430 25284
rect 28578 25228 28588 25284
rect 28644 25228 29372 25284
rect 29428 25228 29438 25284
rect 6374 25116 6412 25172
rect 6468 25116 6478 25172
rect 6636 25116 7756 25172
rect 7812 25116 8540 25172
rect 8596 25116 8606 25172
rect 6636 25060 6692 25116
rect 9266 25060 9276 25116
rect 9332 25060 9380 25116
rect 9436 25060 9484 25116
rect 9540 25060 9550 25116
rect 9660 25060 9716 25228
rect 11228 25060 11284 25228
rect 19292 25172 19348 25228
rect 11890 25116 11900 25172
rect 11956 25116 12684 25172
rect 12740 25116 12750 25172
rect 15474 25116 15484 25172
rect 15540 25116 16268 25172
rect 16324 25116 16334 25172
rect 17724 25116 19068 25172
rect 19124 25116 19134 25172
rect 19292 25116 19516 25172
rect 19572 25116 20636 25172
rect 20692 25116 20702 25172
rect 26114 25116 26124 25172
rect 26180 25116 28476 25172
rect 28532 25116 28542 25172
rect 17330 25060 17340 25116
rect 17396 25060 17444 25116
rect 17500 25060 17548 25116
rect 17604 25060 17614 25116
rect 6626 25004 6636 25060
rect 6692 25004 6702 25060
rect 9660 25004 10556 25060
rect 10612 25004 10622 25060
rect 11228 25004 11340 25060
rect 11396 25004 11406 25060
rect 13234 25004 13244 25060
rect 13300 25004 14924 25060
rect 14980 25004 14990 25060
rect 5170 24892 5180 24948
rect 5236 24892 5964 24948
rect 6020 24892 6300 24948
rect 6356 24892 6366 24948
rect 8642 24892 8652 24948
rect 8708 24892 10892 24948
rect 10948 24892 10958 24948
rect 12534 24892 12572 24948
rect 12628 24892 12638 24948
rect 13010 24892 13020 24948
rect 13076 24892 13132 24948
rect 13188 24892 13356 24948
rect 13412 24892 13422 24948
rect 14466 24892 14476 24948
rect 14532 24892 17388 24948
rect 17444 24892 17454 24948
rect 17724 24836 17780 25116
rect 25394 25060 25404 25116
rect 25460 25060 25508 25116
rect 25564 25060 25612 25116
rect 25668 25060 25678 25116
rect 33458 25060 33468 25116
rect 33524 25060 33572 25116
rect 33628 25060 33676 25116
rect 33732 25060 33742 25116
rect 18498 25004 18508 25060
rect 18564 25004 20188 25060
rect 20244 25004 20254 25060
rect 27430 25004 27468 25060
rect 27524 25004 27534 25060
rect 18386 24892 18396 24948
rect 18452 24892 19628 24948
rect 19684 24892 19694 24948
rect 19842 24892 19852 24948
rect 19908 24892 19946 24948
rect 25554 24892 25564 24948
rect 25620 24892 27244 24948
rect 27300 24892 29596 24948
rect 29652 24892 29662 24948
rect 30706 24892 30716 24948
rect 30772 24892 31276 24948
rect 31332 24892 31342 24948
rect 4498 24780 4508 24836
rect 4564 24780 5292 24836
rect 5348 24780 7308 24836
rect 7364 24780 7374 24836
rect 8754 24780 8764 24836
rect 8820 24780 9996 24836
rect 10052 24780 10062 24836
rect 10994 24780 11004 24836
rect 11060 24780 13468 24836
rect 13524 24780 13534 24836
rect 15138 24780 15148 24836
rect 15204 24780 15260 24836
rect 15316 24780 15326 24836
rect 16258 24780 16268 24836
rect 16324 24780 16716 24836
rect 16772 24780 17780 24836
rect 19506 24780 19516 24836
rect 19572 24780 20300 24836
rect 20356 24780 20366 24836
rect 5506 24668 5516 24724
rect 5572 24668 6636 24724
rect 6692 24668 6702 24724
rect 6962 24668 6972 24724
rect 7028 24668 13804 24724
rect 13860 24668 13870 24724
rect 14130 24668 14140 24724
rect 14196 24668 15932 24724
rect 15988 24668 15998 24724
rect 4610 24556 4620 24612
rect 4676 24556 6524 24612
rect 6580 24556 15260 24612
rect 15316 24556 15326 24612
rect 16268 24500 16324 24780
rect 18162 24668 18172 24724
rect 18228 24668 19292 24724
rect 19348 24668 19358 24724
rect 19730 24668 19740 24724
rect 19796 24668 20412 24724
rect 20468 24668 20478 24724
rect 27682 24668 27692 24724
rect 27748 24668 28140 24724
rect 28196 24668 28206 24724
rect 29698 24668 29708 24724
rect 29764 24668 32508 24724
rect 32564 24668 33964 24724
rect 34020 24668 34030 24724
rect 16818 24556 16828 24612
rect 16884 24556 17500 24612
rect 17556 24556 17566 24612
rect 19058 24556 19068 24612
rect 19124 24556 20300 24612
rect 20356 24556 20366 24612
rect 22642 24556 22652 24612
rect 22708 24556 31948 24612
rect 32004 24556 32014 24612
rect 6402 24444 6412 24500
rect 6468 24444 10108 24500
rect 10164 24444 10174 24500
rect 13906 24444 13916 24500
rect 13972 24444 16324 24500
rect 17602 24444 17612 24500
rect 17668 24444 19852 24500
rect 19908 24444 19918 24500
rect 20178 24444 20188 24500
rect 20244 24444 21196 24500
rect 21252 24444 21262 24500
rect 24882 24444 24892 24500
rect 24948 24444 33180 24500
rect 33236 24444 33246 24500
rect 7298 24332 7308 24388
rect 7364 24332 11900 24388
rect 11956 24332 11966 24388
rect 14354 24332 14364 24388
rect 14420 24332 18508 24388
rect 18564 24332 18574 24388
rect 5234 24276 5244 24332
rect 5300 24276 5348 24332
rect 5404 24276 5452 24332
rect 5508 24276 5518 24332
rect 13298 24276 13308 24332
rect 13364 24276 13412 24332
rect 13468 24276 13516 24332
rect 13572 24276 13582 24332
rect 19852 24276 19908 24444
rect 26198 24332 26236 24388
rect 26292 24332 26302 24388
rect 21362 24276 21372 24332
rect 21428 24276 21476 24332
rect 21532 24276 21580 24332
rect 21636 24276 21646 24332
rect 29426 24276 29436 24332
rect 29492 24276 29540 24332
rect 29596 24276 29644 24332
rect 29700 24276 29710 24332
rect 7410 24220 7420 24276
rect 7476 24220 7868 24276
rect 7924 24220 7934 24276
rect 8530 24220 8540 24276
rect 8596 24220 8876 24276
rect 8932 24220 8942 24276
rect 13794 24220 13804 24276
rect 13860 24220 15036 24276
rect 15092 24220 15102 24276
rect 15250 24220 15260 24276
rect 15316 24220 17500 24276
rect 17556 24220 17566 24276
rect 19852 24220 21196 24276
rect 21252 24220 21262 24276
rect 10434 24108 10444 24164
rect 10500 24108 12348 24164
rect 12404 24108 12414 24164
rect 14914 24108 14924 24164
rect 14980 24108 17052 24164
rect 17108 24108 17118 24164
rect 19394 24108 19404 24164
rect 19460 24108 19852 24164
rect 19908 24108 19918 24164
rect 21858 24108 21868 24164
rect 21924 24108 29428 24164
rect 29698 24108 29708 24164
rect 29764 24108 30268 24164
rect 30324 24108 30334 24164
rect 3938 23996 3948 24052
rect 4004 23996 5964 24052
rect 6020 23996 6030 24052
rect 6290 23996 6300 24052
rect 6356 23996 6636 24052
rect 6692 23996 14140 24052
rect 14196 23996 15372 24052
rect 15428 23996 16604 24052
rect 16660 23996 16670 24052
rect 16930 23996 16940 24052
rect 16996 23996 19180 24052
rect 19236 23996 19246 24052
rect 22418 23996 22428 24052
rect 22484 23996 27020 24052
rect 27076 23996 28812 24052
rect 28868 23996 28878 24052
rect 29372 23940 29428 24108
rect 4834 23884 4844 23940
rect 4900 23884 7196 23940
rect 7252 23884 7262 23940
rect 15026 23884 15036 23940
rect 15092 23884 16268 23940
rect 16324 23884 16334 23940
rect 17042 23884 17052 23940
rect 17108 23884 18732 23940
rect 18788 23884 18798 23940
rect 19282 23884 19292 23940
rect 19348 23884 20076 23940
rect 20132 23884 20142 23940
rect 21970 23884 21980 23940
rect 22036 23884 23436 23940
rect 23492 23884 23502 23940
rect 23660 23884 25900 23940
rect 25956 23884 25966 23940
rect 26898 23884 26908 23940
rect 26964 23884 29148 23940
rect 29204 23884 29214 23940
rect 29372 23884 30268 23940
rect 30324 23884 30334 23940
rect 31938 23884 31948 23940
rect 32004 23884 32732 23940
rect 32788 23884 32798 23940
rect 23660 23828 23716 23884
rect 10098 23772 10108 23828
rect 10164 23772 10668 23828
rect 10724 23772 10734 23828
rect 11218 23772 11228 23828
rect 11284 23772 11564 23828
rect 11620 23772 11630 23828
rect 16146 23772 16156 23828
rect 16212 23772 17948 23828
rect 18004 23772 18014 23828
rect 20626 23772 20636 23828
rect 20692 23772 20972 23828
rect 21028 23772 21038 23828
rect 22866 23772 22876 23828
rect 22932 23772 23716 23828
rect 24210 23772 24220 23828
rect 24276 23772 27244 23828
rect 27300 23772 27310 23828
rect 7634 23660 7644 23716
rect 7700 23660 8428 23716
rect 8484 23660 8494 23716
rect 11218 23660 11228 23716
rect 11284 23660 12236 23716
rect 12292 23660 14140 23716
rect 14196 23660 14206 23716
rect 16370 23660 16380 23716
rect 16436 23660 17164 23716
rect 17220 23660 17230 23716
rect 17602 23660 17612 23716
rect 17668 23660 18060 23716
rect 18116 23660 18126 23716
rect 20066 23660 20076 23716
rect 20132 23660 21868 23716
rect 21924 23660 21934 23716
rect 22082 23660 22092 23716
rect 22148 23660 27020 23716
rect 27076 23660 27086 23716
rect 17826 23548 17836 23604
rect 17892 23548 19964 23604
rect 20020 23548 20030 23604
rect 25890 23548 25900 23604
rect 25956 23548 26572 23604
rect 26628 23548 28476 23604
rect 28532 23548 28542 23604
rect 9266 23492 9276 23548
rect 9332 23492 9380 23548
rect 9436 23492 9484 23548
rect 9540 23492 9550 23548
rect 17330 23492 17340 23548
rect 17396 23492 17444 23548
rect 17500 23492 17548 23548
rect 17604 23492 17614 23548
rect 25394 23492 25404 23548
rect 25460 23492 25508 23548
rect 25564 23492 25612 23548
rect 25668 23492 25678 23548
rect 33458 23492 33468 23548
rect 33524 23492 33572 23548
rect 33628 23492 33676 23548
rect 33732 23492 33742 23548
rect 3332 23436 5404 23492
rect 5460 23436 5470 23492
rect 5842 23436 5852 23492
rect 5908 23436 6636 23492
rect 6692 23436 6702 23492
rect 11778 23436 11788 23492
rect 11844 23436 12236 23492
rect 12292 23436 12302 23492
rect 18610 23436 18620 23492
rect 18676 23436 19852 23492
rect 19908 23436 19918 23492
rect 20850 23436 20860 23492
rect 20916 23436 21308 23492
rect 21364 23436 21924 23492
rect 23874 23436 23884 23492
rect 23940 23436 25228 23492
rect 25284 23436 25294 23492
rect 3332 23380 3388 23436
rect 21868 23380 21924 23436
rect 2482 23324 2492 23380
rect 2548 23324 3388 23380
rect 4946 23324 4956 23380
rect 5012 23324 5740 23380
rect 5796 23324 5806 23380
rect 6962 23324 6972 23380
rect 7028 23324 14084 23380
rect 14690 23324 14700 23380
rect 14756 23324 15708 23380
rect 15764 23324 15774 23380
rect 16146 23324 16156 23380
rect 16212 23324 18508 23380
rect 18564 23324 18574 23380
rect 18946 23324 18956 23380
rect 19012 23324 20412 23380
rect 20468 23324 20478 23380
rect 20626 23324 20636 23380
rect 20692 23324 21644 23380
rect 21700 23324 21710 23380
rect 21868 23324 25844 23380
rect 27346 23324 27356 23380
rect 27412 23324 27692 23380
rect 27748 23324 27758 23380
rect 28466 23324 28476 23380
rect 28532 23324 30492 23380
rect 30548 23324 30558 23380
rect 14028 23268 14084 23324
rect 25788 23268 25844 23324
rect 5058 23212 5068 23268
rect 5124 23212 5852 23268
rect 5908 23212 5918 23268
rect 11666 23212 11676 23268
rect 11732 23212 12348 23268
rect 12404 23212 13972 23268
rect 14028 23212 16156 23268
rect 16212 23212 16222 23268
rect 16370 23212 16380 23268
rect 16436 23212 16474 23268
rect 16706 23212 16716 23268
rect 16772 23212 16782 23268
rect 18722 23212 18732 23268
rect 18788 23212 18798 23268
rect 20188 23212 21756 23268
rect 21812 23212 21822 23268
rect 25218 23212 25228 23268
rect 25284 23212 25732 23268
rect 25788 23212 29372 23268
rect 29428 23212 29438 23268
rect 29922 23212 29932 23268
rect 29988 23212 33180 23268
rect 33236 23212 33246 23268
rect 13916 23156 13972 23212
rect 16716 23156 16772 23212
rect 5282 23100 5292 23156
rect 5348 23100 7308 23156
rect 7364 23100 7374 23156
rect 10882 23100 10892 23156
rect 10948 23100 11564 23156
rect 11620 23100 12012 23156
rect 12068 23100 13692 23156
rect 13748 23100 13758 23156
rect 13916 23100 14252 23156
rect 14308 23100 14318 23156
rect 15026 23100 15036 23156
rect 15092 23100 16772 23156
rect 18732 23044 18788 23212
rect 20188 23156 20244 23212
rect 25676 23156 25732 23212
rect 19282 23100 19292 23156
rect 19348 23100 19358 23156
rect 20178 23100 20188 23156
rect 20244 23100 20254 23156
rect 21522 23100 21532 23156
rect 21588 23100 21598 23156
rect 22530 23100 22540 23156
rect 22596 23100 25452 23156
rect 25508 23100 25518 23156
rect 25676 23100 28252 23156
rect 28308 23100 28318 23156
rect 28690 23100 28700 23156
rect 28756 23100 29484 23156
rect 29540 23100 29550 23156
rect 6626 22988 6636 23044
rect 6692 22988 7196 23044
rect 7252 22988 12684 23044
rect 12740 22988 12750 23044
rect 15092 22988 18788 23044
rect 19292 23044 19348 23100
rect 21532 23044 21588 23100
rect 19292 22988 20132 23044
rect 20850 22988 20860 23044
rect 20916 22988 26796 23044
rect 26852 22988 29708 23044
rect 29764 22988 29774 23044
rect 15092 22932 15148 22988
rect 20076 22932 20132 22988
rect 11442 22876 11452 22932
rect 11508 22876 14812 22932
rect 14868 22876 15148 22932
rect 15810 22876 15820 22932
rect 15876 22876 16604 22932
rect 16660 22876 16670 22932
rect 16818 22876 16828 22932
rect 16884 22876 19852 22932
rect 19908 22876 19918 22932
rect 20076 22876 23436 22932
rect 23492 22876 23502 22932
rect 27234 22876 27244 22932
rect 27300 22876 28140 22932
rect 28196 22876 28206 22932
rect 32610 22876 32620 22932
rect 32676 22876 33068 22932
rect 33124 22876 33134 22932
rect 15698 22764 15708 22820
rect 15764 22764 17500 22820
rect 17556 22764 17566 22820
rect 18470 22764 18508 22820
rect 18564 22764 18574 22820
rect 19058 22764 19068 22820
rect 19124 22764 20188 22820
rect 20244 22764 20254 22820
rect 21858 22764 21868 22820
rect 21924 22764 22988 22820
rect 23044 22764 27132 22820
rect 27188 22764 27198 22820
rect 27906 22764 27916 22820
rect 27972 22764 28364 22820
rect 28420 22764 28430 22820
rect 5234 22708 5244 22764
rect 5300 22708 5348 22764
rect 5404 22708 5452 22764
rect 5508 22708 5518 22764
rect 13298 22708 13308 22764
rect 13364 22708 13412 22764
rect 13468 22708 13516 22764
rect 13572 22708 13582 22764
rect 21362 22708 21372 22764
rect 21428 22708 21476 22764
rect 21532 22708 21580 22764
rect 21636 22708 21646 22764
rect 29426 22708 29436 22764
rect 29492 22708 29540 22764
rect 29596 22708 29644 22764
rect 29700 22708 29710 22764
rect 34200 22708 35000 22736
rect 14802 22652 14812 22708
rect 14868 22652 16492 22708
rect 16548 22652 17836 22708
rect 17892 22652 17902 22708
rect 21746 22652 21756 22708
rect 21812 22652 25844 22708
rect 25788 22596 25844 22652
rect 30604 22652 35000 22708
rect 30604 22596 30660 22652
rect 34200 22624 35000 22652
rect 10322 22540 10332 22596
rect 10388 22540 13580 22596
rect 13636 22540 13646 22596
rect 15138 22540 15148 22596
rect 15204 22540 19180 22596
rect 19236 22540 19740 22596
rect 19796 22540 19806 22596
rect 20738 22540 20748 22596
rect 20804 22540 23884 22596
rect 23940 22540 23950 22596
rect 25228 22540 25564 22596
rect 25620 22540 25630 22596
rect 25788 22540 30660 22596
rect 25228 22484 25284 22540
rect 12898 22428 12908 22484
rect 12964 22428 13804 22484
rect 13860 22428 14588 22484
rect 14644 22428 16380 22484
rect 16436 22428 16446 22484
rect 19842 22428 19852 22484
rect 19908 22428 20636 22484
rect 20692 22428 20702 22484
rect 21644 22428 25284 22484
rect 25442 22428 25452 22484
rect 25508 22428 25788 22484
rect 25844 22428 27804 22484
rect 27860 22428 27870 22484
rect 21644 22372 21700 22428
rect 16258 22316 16268 22372
rect 16324 22316 16380 22372
rect 16436 22316 16446 22372
rect 17378 22316 17388 22372
rect 17444 22316 18844 22372
rect 18900 22316 18910 22372
rect 20412 22316 20524 22372
rect 20580 22316 21700 22372
rect 24434 22316 24444 22372
rect 24500 22316 28140 22372
rect 28196 22316 28206 22372
rect 30258 22316 30268 22372
rect 30324 22316 30940 22372
rect 30996 22316 31006 22372
rect 20412 22260 20468 22316
rect 14466 22204 14476 22260
rect 14532 22204 16772 22260
rect 17938 22204 17948 22260
rect 18004 22204 20468 22260
rect 20626 22204 20636 22260
rect 20692 22204 21420 22260
rect 21476 22204 21486 22260
rect 21634 22204 21644 22260
rect 21700 22204 23940 22260
rect 25218 22204 25228 22260
rect 25284 22204 26796 22260
rect 26852 22204 26862 22260
rect 27794 22204 27804 22260
rect 27860 22204 28476 22260
rect 28532 22204 29484 22260
rect 29540 22204 29550 22260
rect 16716 22148 16772 22204
rect 23884 22148 23940 22204
rect 1810 22092 1820 22148
rect 1876 22092 5068 22148
rect 5124 22092 5134 22148
rect 14018 22092 14028 22148
rect 14084 22092 14700 22148
rect 14756 22092 14766 22148
rect 16706 22092 16716 22148
rect 16772 22092 16782 22148
rect 21298 22092 21308 22148
rect 21364 22092 23212 22148
rect 23268 22092 23278 22148
rect 23874 22092 23884 22148
rect 23940 22092 25116 22148
rect 25172 22092 25182 22148
rect 25554 22092 25564 22148
rect 25620 22092 26124 22148
rect 26180 22092 27020 22148
rect 27076 22092 27086 22148
rect 11442 21980 11452 22036
rect 11508 21980 15036 22036
rect 15092 21980 15102 22036
rect 16006 21980 16044 22036
rect 16100 21980 16110 22036
rect 26786 21980 26796 22036
rect 26852 21980 27132 22036
rect 27188 21980 27198 22036
rect 9266 21924 9276 21980
rect 9332 21924 9380 21980
rect 9436 21924 9484 21980
rect 9540 21924 9550 21980
rect 4610 21868 4620 21924
rect 4676 21868 6244 21924
rect 6188 21812 6244 21868
rect 12908 21812 12964 21980
rect 17330 21924 17340 21980
rect 17396 21924 17444 21980
rect 17500 21924 17548 21980
rect 17604 21924 17614 21980
rect 25394 21924 25404 21980
rect 25460 21924 25508 21980
rect 25564 21924 25612 21980
rect 25668 21924 25678 21980
rect 33458 21924 33468 21980
rect 33524 21924 33572 21980
rect 33628 21924 33676 21980
rect 33732 21924 33742 21980
rect 13682 21868 13692 21924
rect 13748 21868 15820 21924
rect 15876 21868 15886 21924
rect 18274 21868 18284 21924
rect 18340 21868 19964 21924
rect 20020 21868 20030 21924
rect 26852 21868 27244 21924
rect 27300 21868 27310 21924
rect 27906 21868 27916 21924
rect 27972 21868 32620 21924
rect 32676 21868 32686 21924
rect 26852 21812 26908 21868
rect 2482 21756 2492 21812
rect 2548 21756 5292 21812
rect 5348 21756 5358 21812
rect 6178 21756 6188 21812
rect 6244 21756 6748 21812
rect 6804 21756 6814 21812
rect 12898 21756 12908 21812
rect 12964 21756 12974 21812
rect 13570 21756 13580 21812
rect 13636 21756 14364 21812
rect 14420 21756 14430 21812
rect 18386 21756 18396 21812
rect 18452 21756 19180 21812
rect 19236 21756 19246 21812
rect 22754 21756 22764 21812
rect 22820 21756 23772 21812
rect 23828 21756 23838 21812
rect 24220 21756 26348 21812
rect 26404 21756 26908 21812
rect 24220 21700 24276 21756
rect 5842 21644 5852 21700
rect 5908 21644 6076 21700
rect 6132 21644 9548 21700
rect 9604 21644 9614 21700
rect 12226 21644 12236 21700
rect 12292 21644 12572 21700
rect 12628 21644 12638 21700
rect 16482 21644 16492 21700
rect 16548 21644 19068 21700
rect 19124 21644 19134 21700
rect 19394 21644 19404 21700
rect 19460 21644 21644 21700
rect 21700 21644 21756 21700
rect 21812 21644 21822 21700
rect 22306 21644 22316 21700
rect 22372 21644 22382 21700
rect 24210 21644 24220 21700
rect 24276 21644 24286 21700
rect 24434 21644 24444 21700
rect 24500 21644 25340 21700
rect 25396 21644 28252 21700
rect 28308 21644 28318 21700
rect 5282 21532 5292 21588
rect 5348 21532 6972 21588
rect 7028 21532 7038 21588
rect 11106 21532 11116 21588
rect 11172 21532 13468 21588
rect 13524 21532 14812 21588
rect 14868 21532 14878 21588
rect 18722 21532 18732 21588
rect 18788 21532 21980 21588
rect 22036 21532 22046 21588
rect 2482 21420 2492 21476
rect 2548 21420 4172 21476
rect 4228 21420 4238 21476
rect 12450 21420 12460 21476
rect 12516 21420 18396 21476
rect 18452 21420 20524 21476
rect 20580 21420 21868 21476
rect 21924 21420 21934 21476
rect 22316 21364 22372 21644
rect 22754 21532 22764 21588
rect 22820 21532 23660 21588
rect 23716 21532 23726 21588
rect 25778 21532 25788 21588
rect 25844 21532 27468 21588
rect 27524 21532 27534 21588
rect 29810 21532 29820 21588
rect 29876 21532 30268 21588
rect 30324 21532 30334 21588
rect 22530 21420 22540 21476
rect 22596 21420 24892 21476
rect 24948 21420 24958 21476
rect 25330 21420 25340 21476
rect 25396 21420 26572 21476
rect 26628 21420 26638 21476
rect 27122 21420 27132 21476
rect 27188 21420 27244 21476
rect 27300 21420 27310 21476
rect 28130 21420 28140 21476
rect 28196 21420 32396 21476
rect 32452 21420 32462 21476
rect 15474 21308 15484 21364
rect 15540 21308 17388 21364
rect 17444 21308 22372 21364
rect 24770 21308 24780 21364
rect 24836 21308 27692 21364
rect 27748 21308 27758 21364
rect 21858 21196 21868 21252
rect 21924 21196 22316 21252
rect 22372 21196 22876 21252
rect 22932 21196 27188 21252
rect 27346 21196 27356 21252
rect 27412 21196 28924 21252
rect 28980 21196 28990 21252
rect 5234 21140 5244 21196
rect 5300 21140 5348 21196
rect 5404 21140 5452 21196
rect 5508 21140 5518 21196
rect 13298 21140 13308 21196
rect 13364 21140 13412 21196
rect 13468 21140 13516 21196
rect 13572 21140 13582 21196
rect 21362 21140 21372 21196
rect 21428 21140 21476 21196
rect 21532 21140 21580 21196
rect 21636 21140 21646 21196
rect 27132 21140 27188 21196
rect 29426 21140 29436 21196
rect 29492 21140 29540 21196
rect 29596 21140 29644 21196
rect 29700 21140 29710 21196
rect 21746 21084 21756 21140
rect 21812 21084 25788 21140
rect 25844 21084 25854 21140
rect 26870 21084 26908 21140
rect 26964 21084 26974 21140
rect 27132 21084 28588 21140
rect 28644 21084 28654 21140
rect 6626 20972 6636 21028
rect 6692 20972 7308 21028
rect 7364 20972 7374 21028
rect 13794 20972 13804 21028
rect 13860 20972 20972 21028
rect 21028 20972 21038 21028
rect 22978 20972 22988 21028
rect 23044 20972 29372 21028
rect 29428 20972 29438 21028
rect 8978 20860 8988 20916
rect 9044 20860 9660 20916
rect 9716 20860 10108 20916
rect 10164 20860 10174 20916
rect 13458 20860 13468 20916
rect 13524 20860 14252 20916
rect 14308 20860 14318 20916
rect 16930 20860 16940 20916
rect 16996 20860 22652 20916
rect 22708 20860 22718 20916
rect 26114 20860 26124 20916
rect 26180 20860 27020 20916
rect 27076 20860 27086 20916
rect 4610 20748 4620 20804
rect 4676 20748 4956 20804
rect 5012 20748 6860 20804
rect 6916 20748 7308 20804
rect 7364 20748 8428 20804
rect 8484 20748 8494 20804
rect 16594 20748 16604 20804
rect 16660 20748 17836 20804
rect 17892 20748 17902 20804
rect 27132 20748 29148 20804
rect 29204 20748 29214 20804
rect 27132 20692 27188 20748
rect 17612 20636 18844 20692
rect 18900 20636 18910 20692
rect 21746 20636 21756 20692
rect 21812 20636 27188 20692
rect 28578 20636 28588 20692
rect 28644 20636 32396 20692
rect 32452 20636 32462 20692
rect 17612 20580 17668 20636
rect 4610 20524 4620 20580
rect 4676 20524 5740 20580
rect 5796 20524 11228 20580
rect 11284 20524 11294 20580
rect 12226 20524 12236 20580
rect 12292 20524 17612 20580
rect 17668 20524 17678 20580
rect 18274 20524 18284 20580
rect 18340 20524 19628 20580
rect 19684 20524 19694 20580
rect 22642 20524 22652 20580
rect 22708 20524 24668 20580
rect 24724 20524 26796 20580
rect 26852 20524 32172 20580
rect 32228 20524 32956 20580
rect 33012 20524 33022 20580
rect 9874 20412 9884 20468
rect 9940 20412 11116 20468
rect 11172 20412 11564 20468
rect 11620 20412 11630 20468
rect 14802 20412 14812 20468
rect 14868 20412 15036 20468
rect 15092 20412 15102 20468
rect 29138 20412 29148 20468
rect 29204 20412 33180 20468
rect 33236 20412 33246 20468
rect 9266 20356 9276 20412
rect 9332 20356 9380 20412
rect 9436 20356 9484 20412
rect 9540 20356 9550 20412
rect 17330 20356 17340 20412
rect 17396 20356 17444 20412
rect 17500 20356 17548 20412
rect 17604 20356 17614 20412
rect 25394 20356 25404 20412
rect 25460 20356 25508 20412
rect 25564 20356 25612 20412
rect 25668 20356 25678 20412
rect 33458 20356 33468 20412
rect 33524 20356 33572 20412
rect 33628 20356 33676 20412
rect 33732 20356 33742 20412
rect 5058 20300 5068 20356
rect 5124 20300 5740 20356
rect 5796 20300 7196 20356
rect 7252 20300 7262 20356
rect 26534 20300 26572 20356
rect 26628 20300 26638 20356
rect 27206 20300 27244 20356
rect 27300 20300 27310 20356
rect 29250 20300 29260 20356
rect 29316 20300 31052 20356
rect 31108 20300 31118 20356
rect 7196 20244 7252 20300
rect 7196 20188 9548 20244
rect 9604 20188 10332 20244
rect 10388 20188 10398 20244
rect 15250 20188 15260 20244
rect 15316 20188 16156 20244
rect 16212 20188 16222 20244
rect 17490 20188 17500 20244
rect 17556 20188 18732 20244
rect 18788 20188 18798 20244
rect 21410 20188 21420 20244
rect 21476 20188 25228 20244
rect 25284 20188 25340 20244
rect 25396 20188 25406 20244
rect 25666 20188 25676 20244
rect 25732 20188 25788 20244
rect 25844 20188 32060 20244
rect 32116 20188 32126 20244
rect 5394 20076 5404 20132
rect 5460 20076 7980 20132
rect 8036 20076 8046 20132
rect 10882 20076 10892 20132
rect 10948 20076 11452 20132
rect 11508 20076 12572 20132
rect 12628 20076 12638 20132
rect 13682 20076 13692 20132
rect 13748 20076 14476 20132
rect 14532 20076 14542 20132
rect 15810 20076 15820 20132
rect 15876 20076 20076 20132
rect 20132 20076 20972 20132
rect 21028 20076 22204 20132
rect 22260 20076 22270 20132
rect 22866 20076 22876 20132
rect 22932 20076 23884 20132
rect 23940 20076 24892 20132
rect 24948 20076 24958 20132
rect 25452 20076 26908 20132
rect 26964 20076 26974 20132
rect 27570 20076 27580 20132
rect 27636 20076 29932 20132
rect 29988 20076 29998 20132
rect 30230 20076 30268 20132
rect 30324 20076 30334 20132
rect 31490 20076 31500 20132
rect 31556 20076 32732 20132
rect 32788 20076 32798 20132
rect 4610 19964 4620 20020
rect 4676 19964 6076 20020
rect 6132 19964 6412 20020
rect 6468 19964 6478 20020
rect 9762 19964 9772 20020
rect 9828 19964 12908 20020
rect 12964 19964 12974 20020
rect 14354 19964 14364 20020
rect 14420 19964 15036 20020
rect 15092 19964 15102 20020
rect 20514 19964 20524 20020
rect 20580 19964 21756 20020
rect 21812 19964 21822 20020
rect 21970 19964 21980 20020
rect 22036 19964 22428 20020
rect 22484 19964 24220 20020
rect 24276 19964 24286 20020
rect 25452 19908 25508 20076
rect 34200 20020 35000 20048
rect 7634 19852 7644 19908
rect 7700 19852 7980 19908
rect 8036 19852 8652 19908
rect 8708 19852 10780 19908
rect 10836 19852 10846 19908
rect 19394 19852 19404 19908
rect 19460 19852 21868 19908
rect 21924 19852 21934 19908
rect 23762 19852 23772 19908
rect 23828 19852 25508 19908
rect 25788 19964 26908 20020
rect 26964 19964 26974 20020
rect 27234 19964 27244 20020
rect 27300 19964 29148 20020
rect 29204 19964 29214 20020
rect 29362 19964 29372 20020
rect 29428 19964 31052 20020
rect 31108 19964 31118 20020
rect 31276 19964 35000 20020
rect 25788 19796 25844 19964
rect 31276 19908 31332 19964
rect 34200 19936 35000 19964
rect 26982 19852 27020 19908
rect 27076 19852 27086 19908
rect 27906 19852 27916 19908
rect 27972 19852 28364 19908
rect 28420 19852 28430 19908
rect 29026 19852 29036 19908
rect 29092 19852 31332 19908
rect 32162 19852 32172 19908
rect 32228 19852 32732 19908
rect 32788 19852 32798 19908
rect 5170 19740 5180 19796
rect 5236 19740 5852 19796
rect 5908 19740 5918 19796
rect 7522 19740 7532 19796
rect 7588 19740 21532 19796
rect 21588 19740 21980 19796
rect 22036 19740 22046 19796
rect 24770 19740 24780 19796
rect 24836 19740 25844 19796
rect 26002 19740 26012 19796
rect 26068 19740 28084 19796
rect 24098 19628 24108 19684
rect 24164 19628 27860 19684
rect 5234 19572 5244 19628
rect 5300 19572 5348 19628
rect 5404 19572 5452 19628
rect 5508 19572 5518 19628
rect 13298 19572 13308 19628
rect 13364 19572 13412 19628
rect 13468 19572 13516 19628
rect 13572 19572 13582 19628
rect 21362 19572 21372 19628
rect 21428 19572 21476 19628
rect 21532 19572 21580 19628
rect 21636 19572 21646 19628
rect 14998 19516 15036 19572
rect 15092 19516 15102 19572
rect 17042 19516 17052 19572
rect 17108 19516 17118 19572
rect 26450 19516 26460 19572
rect 26516 19516 27132 19572
rect 27188 19516 27198 19572
rect 27570 19516 27580 19572
rect 27636 19516 27646 19572
rect 17052 19460 17108 19516
rect 4050 19404 4060 19460
rect 4116 19404 5740 19460
rect 5796 19404 5806 19460
rect 17052 19404 21868 19460
rect 21924 19404 21934 19460
rect 23090 19404 23100 19460
rect 23156 19404 24332 19460
rect 24388 19404 24398 19460
rect 12898 19292 12908 19348
rect 12964 19292 14140 19348
rect 14196 19292 15148 19348
rect 19058 19292 19068 19348
rect 19124 19292 20300 19348
rect 20356 19292 20860 19348
rect 20916 19292 20926 19348
rect 22988 19292 24108 19348
rect 24164 19292 24174 19348
rect 25442 19292 25452 19348
rect 25508 19292 25788 19348
rect 25844 19292 26236 19348
rect 26292 19292 26302 19348
rect 15092 19236 15148 19292
rect 22988 19236 23044 19292
rect 27580 19236 27636 19516
rect 9650 19180 9660 19236
rect 9716 19180 13300 19236
rect 15092 19180 16828 19236
rect 16884 19180 16894 19236
rect 22978 19180 22988 19236
rect 23044 19180 23054 19236
rect 23548 19180 27636 19236
rect 13244 19124 13300 19180
rect 23548 19124 23604 19180
rect 27804 19124 27860 19628
rect 28028 19460 28084 19740
rect 29922 19628 29932 19684
rect 29988 19628 33180 19684
rect 33236 19628 33246 19684
rect 29426 19572 29436 19628
rect 29492 19572 29540 19628
rect 29596 19572 29644 19628
rect 29700 19572 29710 19628
rect 28018 19404 28028 19460
rect 28084 19404 29148 19460
rect 29204 19404 29214 19460
rect 29474 19404 29484 19460
rect 29540 19404 31612 19460
rect 31668 19404 33068 19460
rect 33124 19404 33134 19460
rect 28242 19180 28252 19236
rect 28308 19180 28476 19236
rect 28532 19180 28542 19236
rect 28690 19180 28700 19236
rect 28756 19180 30604 19236
rect 30660 19180 30670 19236
rect 33058 19180 33068 19236
rect 33124 19180 33852 19236
rect 33908 19180 33918 19236
rect 3602 19068 3612 19124
rect 3668 19068 4620 19124
rect 4676 19068 6300 19124
rect 6356 19068 6366 19124
rect 9090 19068 9100 19124
rect 9156 19068 11004 19124
rect 11060 19068 11070 19124
rect 11554 19068 11564 19124
rect 11620 19068 12348 19124
rect 12404 19068 13020 19124
rect 13076 19068 13086 19124
rect 13244 19068 15988 19124
rect 16146 19068 16156 19124
rect 16212 19068 17724 19124
rect 17780 19068 20412 19124
rect 20468 19068 20478 19124
rect 23538 19068 23548 19124
rect 23604 19068 23614 19124
rect 24994 19068 25004 19124
rect 25060 19068 26908 19124
rect 27804 19068 30268 19124
rect 30324 19068 30334 19124
rect 11004 19012 11060 19068
rect 15932 19012 15988 19068
rect 26852 19012 26908 19068
rect 4498 18956 4508 19012
rect 4564 18956 5292 19012
rect 5348 18956 5740 19012
rect 5796 18956 8876 19012
rect 8932 18956 8942 19012
rect 11004 18956 11676 19012
rect 11732 18956 11742 19012
rect 15932 18956 17500 19012
rect 17556 18956 18284 19012
rect 18340 18956 26684 19012
rect 26740 18956 26750 19012
rect 26852 18956 29148 19012
rect 29204 18956 29214 19012
rect 12086 18844 12124 18900
rect 12180 18844 12190 18900
rect 13682 18844 13692 18900
rect 13748 18844 16044 18900
rect 16100 18844 16110 18900
rect 18386 18844 18396 18900
rect 18452 18844 20748 18900
rect 20804 18844 20814 18900
rect 22306 18844 22316 18900
rect 22372 18844 23772 18900
rect 23828 18844 23838 18900
rect 25778 18844 25788 18900
rect 25844 18844 26572 18900
rect 26628 18844 27244 18900
rect 27300 18844 27310 18900
rect 27458 18844 27468 18900
rect 27524 18844 28476 18900
rect 28532 18844 28542 18900
rect 30146 18844 30156 18900
rect 30212 18844 32060 18900
rect 32116 18844 32126 18900
rect 9266 18788 9276 18844
rect 9332 18788 9380 18844
rect 9436 18788 9484 18844
rect 9540 18788 9550 18844
rect 17330 18788 17340 18844
rect 17396 18788 17444 18844
rect 17500 18788 17548 18844
rect 17604 18788 17614 18844
rect 25394 18788 25404 18844
rect 25460 18788 25508 18844
rect 25564 18788 25612 18844
rect 25668 18788 25678 18844
rect 33458 18788 33468 18844
rect 33524 18788 33572 18844
rect 33628 18788 33676 18844
rect 33732 18788 33742 18844
rect 3332 18732 3612 18788
rect 3668 18732 3678 18788
rect 8194 18732 8204 18788
rect 8260 18732 9100 18788
rect 9156 18732 9166 18788
rect 9762 18732 9772 18788
rect 9828 18732 9838 18788
rect 13906 18732 13916 18788
rect 13972 18732 15036 18788
rect 15092 18732 15102 18788
rect 21858 18732 21868 18788
rect 21924 18732 22988 18788
rect 23044 18732 23324 18788
rect 23380 18732 23390 18788
rect 27794 18732 27804 18788
rect 27860 18732 28364 18788
rect 28420 18732 30324 18788
rect 30482 18732 30492 18788
rect 30548 18732 31276 18788
rect 31332 18732 31342 18788
rect 3332 18676 3388 18732
rect 9772 18676 9828 18732
rect 30268 18676 30324 18732
rect 3042 18620 3052 18676
rect 3108 18620 3388 18676
rect 3714 18620 3724 18676
rect 3780 18620 5180 18676
rect 5236 18620 5964 18676
rect 6020 18620 6030 18676
rect 9202 18620 9212 18676
rect 9268 18620 9828 18676
rect 11778 18620 11788 18676
rect 11844 18620 12012 18676
rect 12068 18620 13132 18676
rect 13188 18620 13804 18676
rect 13860 18620 13870 18676
rect 14466 18620 14476 18676
rect 14532 18620 15484 18676
rect 15540 18620 17052 18676
rect 17108 18620 17118 18676
rect 18610 18620 18620 18676
rect 18676 18620 19404 18676
rect 19460 18620 19470 18676
rect 24098 18620 24108 18676
rect 24164 18620 26460 18676
rect 26516 18620 26526 18676
rect 26786 18620 26796 18676
rect 26852 18620 27916 18676
rect 27972 18620 27982 18676
rect 28690 18620 28700 18676
rect 28756 18620 29596 18676
rect 29652 18620 29662 18676
rect 30268 18620 32172 18676
rect 32228 18620 32238 18676
rect 5058 18508 5068 18564
rect 5124 18508 5292 18564
rect 5348 18508 5358 18564
rect 8530 18508 8540 18564
rect 8596 18508 8988 18564
rect 9044 18508 9660 18564
rect 9716 18508 9726 18564
rect 15586 18508 15596 18564
rect 15652 18508 16156 18564
rect 16212 18508 16222 18564
rect 19058 18508 19068 18564
rect 19124 18508 19964 18564
rect 20020 18508 20030 18564
rect 20178 18508 20188 18564
rect 20244 18508 20860 18564
rect 20916 18508 22316 18564
rect 22372 18508 22382 18564
rect 22754 18508 22764 18564
rect 22820 18508 23436 18564
rect 23492 18508 23502 18564
rect 23762 18508 23772 18564
rect 23828 18508 26124 18564
rect 26180 18508 26190 18564
rect 26898 18508 26908 18564
rect 26964 18508 27692 18564
rect 27748 18508 28364 18564
rect 28420 18508 28430 18564
rect 29484 18508 29932 18564
rect 29988 18508 29998 18564
rect 8540 18452 8596 18508
rect 29484 18452 29540 18508
rect 3266 18396 3276 18452
rect 3332 18396 3948 18452
rect 4004 18396 4014 18452
rect 4386 18396 4396 18452
rect 4452 18396 4844 18452
rect 4900 18396 4910 18452
rect 6290 18396 6300 18452
rect 6356 18396 6748 18452
rect 6804 18396 8596 18452
rect 11106 18396 11116 18452
rect 11172 18396 12012 18452
rect 12068 18396 12078 18452
rect 13906 18396 13916 18452
rect 13972 18396 13982 18452
rect 14802 18396 14812 18452
rect 14868 18396 15260 18452
rect 15316 18396 15326 18452
rect 15810 18396 15820 18452
rect 15876 18396 15886 18452
rect 16034 18396 16044 18452
rect 16100 18396 16138 18452
rect 19842 18396 19852 18452
rect 19908 18396 20188 18452
rect 20244 18396 21644 18452
rect 21700 18396 21710 18452
rect 22082 18396 22092 18452
rect 22148 18396 25004 18452
rect 25060 18396 25070 18452
rect 25890 18396 25900 18452
rect 25956 18396 27804 18452
rect 27860 18396 27870 18452
rect 28028 18396 28588 18452
rect 28644 18396 29148 18452
rect 29204 18396 29214 18452
rect 29474 18396 29484 18452
rect 29540 18396 29550 18452
rect 30902 18396 30940 18452
rect 30996 18396 31006 18452
rect 32498 18396 32508 18452
rect 32564 18396 33292 18452
rect 33348 18396 33358 18452
rect 13916 18340 13972 18396
rect 15820 18340 15876 18396
rect 28028 18340 28084 18396
rect 2482 18284 2492 18340
rect 2548 18284 4172 18340
rect 4228 18284 4238 18340
rect 9874 18284 9884 18340
rect 9940 18284 11228 18340
rect 11284 18284 11294 18340
rect 13916 18284 15876 18340
rect 20738 18284 20748 18340
rect 20804 18284 25452 18340
rect 25508 18284 25518 18340
rect 27244 18284 28084 18340
rect 28242 18284 28252 18340
rect 28308 18284 29260 18340
rect 29316 18284 29326 18340
rect 29698 18284 29708 18340
rect 29764 18284 31052 18340
rect 31108 18284 31118 18340
rect 27244 18228 27300 18284
rect 3490 18172 3500 18228
rect 3556 18172 5628 18228
rect 5684 18172 5694 18228
rect 10882 18172 10892 18228
rect 10948 18172 14028 18228
rect 14084 18172 14476 18228
rect 14532 18172 14542 18228
rect 21858 18172 21868 18228
rect 21924 18172 27300 18228
rect 27458 18172 27468 18228
rect 27524 18172 28812 18228
rect 28868 18172 29820 18228
rect 29876 18172 29886 18228
rect 28690 18060 28700 18116
rect 28756 18060 28868 18116
rect 30258 18060 30268 18116
rect 30324 18060 31724 18116
rect 31780 18060 31790 18116
rect 5234 18004 5244 18060
rect 5300 18004 5348 18060
rect 5404 18004 5452 18060
rect 5508 18004 5518 18060
rect 13298 18004 13308 18060
rect 13364 18004 13412 18060
rect 13468 18004 13516 18060
rect 13572 18004 13582 18060
rect 21362 18004 21372 18060
rect 21428 18004 21476 18060
rect 21532 18004 21580 18060
rect 21636 18004 21646 18060
rect 19954 17948 19964 18004
rect 20020 17948 20524 18004
rect 20580 17948 20590 18004
rect 21970 17948 21980 18004
rect 22036 17948 28588 18004
rect 28644 17948 28654 18004
rect 28812 17892 28868 18060
rect 29426 18004 29436 18060
rect 29492 18004 29540 18060
rect 29596 18004 29644 18060
rect 29700 18004 29710 18060
rect 7158 17836 7196 17892
rect 7252 17836 7262 17892
rect 17602 17836 17612 17892
rect 17668 17836 18620 17892
rect 18676 17836 29372 17892
rect 29428 17836 29438 17892
rect 31490 17836 31500 17892
rect 31556 17836 31566 17892
rect 31500 17780 31556 17836
rect 3938 17724 3948 17780
rect 4004 17724 4508 17780
rect 4564 17724 6748 17780
rect 6804 17724 6814 17780
rect 11732 17724 15932 17780
rect 15988 17724 15998 17780
rect 20626 17724 20636 17780
rect 20692 17724 21980 17780
rect 22036 17724 22046 17780
rect 22194 17724 22204 17780
rect 22260 17724 23212 17780
rect 23268 17724 23278 17780
rect 24770 17724 24780 17780
rect 24836 17724 26348 17780
rect 26404 17724 26414 17780
rect 28476 17724 31556 17780
rect 11732 17668 11788 17724
rect 28476 17668 28532 17724
rect 5814 17612 5852 17668
rect 5908 17612 11340 17668
rect 11396 17612 11788 17668
rect 12450 17612 12460 17668
rect 12516 17612 12908 17668
rect 12964 17612 13580 17668
rect 13636 17612 13646 17668
rect 18722 17612 18732 17668
rect 18788 17612 20300 17668
rect 20356 17612 21308 17668
rect 21364 17612 21374 17668
rect 24658 17612 24668 17668
rect 24724 17612 25900 17668
rect 25956 17612 26236 17668
rect 26292 17612 26302 17668
rect 26758 17612 26796 17668
rect 26852 17612 26862 17668
rect 27234 17612 27244 17668
rect 27300 17612 27916 17668
rect 27972 17612 27982 17668
rect 28130 17612 28140 17668
rect 28196 17612 28476 17668
rect 28532 17612 28542 17668
rect 29250 17612 29260 17668
rect 29316 17612 30044 17668
rect 30100 17612 30110 17668
rect 2482 17500 2492 17556
rect 2548 17500 4508 17556
rect 4564 17500 4574 17556
rect 8530 17500 8540 17556
rect 8596 17500 12236 17556
rect 12292 17500 12302 17556
rect 16706 17500 16716 17556
rect 16772 17500 22540 17556
rect 22596 17500 23884 17556
rect 23940 17500 23950 17556
rect 25330 17500 25340 17556
rect 25396 17500 26124 17556
rect 26180 17500 26190 17556
rect 32050 17500 32060 17556
rect 32116 17500 32956 17556
rect 33012 17500 33022 17556
rect 7074 17388 7084 17444
rect 7140 17388 7756 17444
rect 7812 17388 8204 17444
rect 8260 17388 10668 17444
rect 10724 17388 10734 17444
rect 18610 17388 18620 17444
rect 18676 17388 19404 17444
rect 19460 17388 19470 17444
rect 19842 17388 19852 17444
rect 19908 17388 20524 17444
rect 20580 17388 22204 17444
rect 22260 17388 22270 17444
rect 24546 17388 24556 17444
rect 24612 17388 27356 17444
rect 27412 17388 27692 17444
rect 27748 17388 27758 17444
rect 28438 17388 28476 17444
rect 28532 17388 28542 17444
rect 34200 17332 35000 17360
rect 21970 17276 21980 17332
rect 22036 17276 22988 17332
rect 23044 17276 23054 17332
rect 26982 17276 27020 17332
rect 27076 17276 27086 17332
rect 27234 17276 27244 17332
rect 27300 17276 28140 17332
rect 28196 17276 28206 17332
rect 33852 17276 35000 17332
rect 9266 17220 9276 17276
rect 9332 17220 9380 17276
rect 9436 17220 9484 17276
rect 9540 17220 9550 17276
rect 17330 17220 17340 17276
rect 17396 17220 17444 17276
rect 17500 17220 17548 17276
rect 17604 17220 17614 17276
rect 25394 17220 25404 17276
rect 25460 17220 25508 17276
rect 25564 17220 25612 17276
rect 25668 17220 25678 17276
rect 33458 17220 33468 17276
rect 33524 17220 33572 17276
rect 33628 17220 33676 17276
rect 33732 17220 33742 17276
rect 5170 17164 5180 17220
rect 5236 17164 5404 17220
rect 5460 17164 7532 17220
rect 7588 17164 7598 17220
rect 11778 17164 11788 17220
rect 11844 17164 12684 17220
rect 12740 17164 15148 17220
rect 17938 17164 17948 17220
rect 18004 17164 19628 17220
rect 19684 17164 21084 17220
rect 21140 17164 21150 17220
rect 26114 17164 26124 17220
rect 26180 17164 28252 17220
rect 28308 17164 28318 17220
rect 30482 17164 30492 17220
rect 30548 17164 31164 17220
rect 31220 17164 31230 17220
rect 15092 17108 15148 17164
rect 33852 17108 33908 17276
rect 34200 17248 35000 17276
rect 4722 17052 4732 17108
rect 4788 17052 6636 17108
rect 6692 17052 6702 17108
rect 15092 17052 26572 17108
rect 26628 17052 26638 17108
rect 26786 17052 26796 17108
rect 26852 17052 27132 17108
rect 27188 17052 28364 17108
rect 28420 17052 28430 17108
rect 29810 17052 29820 17108
rect 29876 17052 33908 17108
rect 6290 16940 6300 16996
rect 6356 16940 7644 16996
rect 7700 16940 7868 16996
rect 7924 16940 8428 16996
rect 8484 16940 8494 16996
rect 12562 16940 12572 16996
rect 12628 16940 20636 16996
rect 20692 16940 20702 16996
rect 21634 16940 21644 16996
rect 21700 16940 23548 16996
rect 23604 16940 23614 16996
rect 26002 16940 26012 16996
rect 26068 16940 26684 16996
rect 26740 16940 28700 16996
rect 28756 16940 28766 16996
rect 29362 16940 29372 16996
rect 29428 16940 31948 16996
rect 32004 16940 33180 16996
rect 33236 16940 33246 16996
rect 7074 16828 7084 16884
rect 7140 16828 7532 16884
rect 7588 16828 7598 16884
rect 11554 16828 11564 16884
rect 11620 16828 12460 16884
rect 12516 16828 13132 16884
rect 13188 16828 13916 16884
rect 13972 16828 13982 16884
rect 16818 16828 16828 16884
rect 16884 16828 17948 16884
rect 18004 16828 18014 16884
rect 23202 16828 23212 16884
rect 23268 16828 23436 16884
rect 23492 16828 27020 16884
rect 27076 16828 27356 16884
rect 27412 16828 27422 16884
rect 27804 16828 31500 16884
rect 31556 16828 31566 16884
rect 27804 16772 27860 16828
rect 30268 16772 30324 16828
rect 18834 16716 18844 16772
rect 18900 16716 20412 16772
rect 20468 16716 20478 16772
rect 23538 16716 23548 16772
rect 23604 16716 24444 16772
rect 24500 16716 25116 16772
rect 25172 16716 25182 16772
rect 27794 16716 27804 16772
rect 27860 16716 27870 16772
rect 30258 16716 30268 16772
rect 30324 16716 30334 16772
rect 4162 16604 4172 16660
rect 4228 16604 4844 16660
rect 4900 16604 4910 16660
rect 18162 16604 18172 16660
rect 18228 16604 18732 16660
rect 18788 16604 18798 16660
rect 25554 16604 25564 16660
rect 25620 16604 26124 16660
rect 26180 16604 26190 16660
rect 19394 16492 19404 16548
rect 19460 16492 20188 16548
rect 20244 16492 20254 16548
rect 5234 16436 5244 16492
rect 5300 16436 5348 16492
rect 5404 16436 5452 16492
rect 5508 16436 5518 16492
rect 13298 16436 13308 16492
rect 13364 16436 13412 16492
rect 13468 16436 13516 16492
rect 13572 16436 13582 16492
rect 21362 16436 21372 16492
rect 21428 16436 21476 16492
rect 21532 16436 21580 16492
rect 21636 16436 21646 16492
rect 29426 16436 29436 16492
rect 29492 16436 29540 16492
rect 29596 16436 29644 16492
rect 29700 16436 29710 16492
rect 15026 16268 15036 16324
rect 15092 16268 23548 16324
rect 23604 16268 23614 16324
rect 25106 16156 25116 16212
rect 25172 16156 28308 16212
rect 28690 16156 28700 16212
rect 28756 16156 28766 16212
rect 28252 16100 28308 16156
rect 28700 16100 28756 16156
rect 4946 16044 4956 16100
rect 5012 16044 5628 16100
rect 5684 16044 5694 16100
rect 10882 16044 10892 16100
rect 10948 16044 11676 16100
rect 11732 16044 11742 16100
rect 17826 16044 17836 16100
rect 17892 16044 19068 16100
rect 19124 16044 19292 16100
rect 19348 16044 19358 16100
rect 22642 16044 22652 16100
rect 22708 16044 27020 16100
rect 27076 16044 27086 16100
rect 28242 16044 28252 16100
rect 28308 16044 28318 16100
rect 28700 16044 28924 16100
rect 28980 16044 28990 16100
rect 29138 16044 29148 16100
rect 29204 16044 29372 16100
rect 29428 16044 32956 16100
rect 33012 16044 33022 16100
rect 17602 15932 17612 15988
rect 17668 15932 21532 15988
rect 21588 15932 21598 15988
rect 22530 15932 22540 15988
rect 22596 15932 24556 15988
rect 24612 15932 24622 15988
rect 24994 15932 25004 15988
rect 25060 15932 25844 15988
rect 26002 15932 26012 15988
rect 26068 15932 28308 15988
rect 25788 15876 25844 15932
rect 2482 15820 2492 15876
rect 2548 15820 4508 15876
rect 4564 15820 4574 15876
rect 6626 15820 6636 15876
rect 6692 15820 6702 15876
rect 18162 15820 18172 15876
rect 18228 15820 18620 15876
rect 18676 15820 18686 15876
rect 19282 15820 19292 15876
rect 19348 15820 19740 15876
rect 19796 15820 19806 15876
rect 20076 15820 21644 15876
rect 21700 15820 23212 15876
rect 23268 15820 23278 15876
rect 24658 15820 24668 15876
rect 24724 15820 25564 15876
rect 25620 15820 25630 15876
rect 25788 15820 26068 15876
rect 6636 15764 6692 15820
rect 20076 15764 20132 15820
rect 3938 15708 3948 15764
rect 4004 15708 5852 15764
rect 5908 15708 6692 15764
rect 18834 15708 18844 15764
rect 18900 15708 20076 15764
rect 20132 15708 20142 15764
rect 24098 15708 24108 15764
rect 24164 15708 25116 15764
rect 25172 15708 25182 15764
rect 9266 15652 9276 15708
rect 9332 15652 9380 15708
rect 9436 15652 9484 15708
rect 9540 15652 9550 15708
rect 17330 15652 17340 15708
rect 17396 15652 17444 15708
rect 17500 15652 17548 15708
rect 17604 15652 17614 15708
rect 25394 15652 25404 15708
rect 25460 15652 25508 15708
rect 25564 15652 25612 15708
rect 25668 15652 25678 15708
rect 26012 15652 26068 15820
rect 28252 15764 28308 15932
rect 27010 15708 27020 15764
rect 27076 15708 27468 15764
rect 27524 15708 27534 15764
rect 28242 15708 28252 15764
rect 28308 15708 29260 15764
rect 29316 15708 30156 15764
rect 30212 15708 30222 15764
rect 33458 15652 33468 15708
rect 33524 15652 33572 15708
rect 33628 15652 33676 15708
rect 33732 15652 33742 15708
rect 17836 15596 20188 15652
rect 20244 15596 20254 15652
rect 26002 15596 26012 15652
rect 26068 15596 28476 15652
rect 28532 15596 28542 15652
rect 30258 15596 30268 15652
rect 30324 15596 32508 15652
rect 32564 15596 32574 15652
rect 17836 15540 17892 15596
rect 4610 15484 4620 15540
rect 4676 15484 5292 15540
rect 5348 15484 5740 15540
rect 5796 15484 5806 15540
rect 6178 15484 6188 15540
rect 6244 15484 6748 15540
rect 6804 15484 6814 15540
rect 12562 15484 12572 15540
rect 12628 15484 17836 15540
rect 17892 15484 17902 15540
rect 18050 15484 18060 15540
rect 18116 15484 18508 15540
rect 18564 15484 18574 15540
rect 18834 15484 18844 15540
rect 18900 15484 19292 15540
rect 19348 15484 21196 15540
rect 21252 15484 21262 15540
rect 22866 15484 22876 15540
rect 22932 15484 23884 15540
rect 23940 15484 25116 15540
rect 25172 15484 25182 15540
rect 25554 15484 25564 15540
rect 25620 15484 29932 15540
rect 29988 15484 29998 15540
rect 6402 15372 6412 15428
rect 6468 15372 6972 15428
rect 7028 15372 7038 15428
rect 7186 15372 7196 15428
rect 7252 15372 8316 15428
rect 8372 15372 8652 15428
rect 8708 15372 10220 15428
rect 10276 15372 10286 15428
rect 13346 15372 13356 15428
rect 13412 15372 14028 15428
rect 14084 15372 14700 15428
rect 14756 15372 14766 15428
rect 16594 15372 16604 15428
rect 16660 15372 17948 15428
rect 18004 15372 18014 15428
rect 18722 15372 18732 15428
rect 18788 15372 19964 15428
rect 20020 15372 20524 15428
rect 20580 15372 20590 15428
rect 21634 15372 21644 15428
rect 21700 15372 21710 15428
rect 23538 15372 23548 15428
rect 23604 15372 24444 15428
rect 24500 15372 24510 15428
rect 25778 15372 25788 15428
rect 25844 15372 25900 15428
rect 25956 15372 25966 15428
rect 26114 15372 26124 15428
rect 26180 15372 26796 15428
rect 26852 15372 26862 15428
rect 28662 15372 28700 15428
rect 28756 15372 33180 15428
rect 33236 15372 33246 15428
rect 21644 15316 21700 15372
rect 5394 15260 5404 15316
rect 5460 15260 6300 15316
rect 6356 15260 6366 15316
rect 6514 15260 6524 15316
rect 6580 15260 7980 15316
rect 8036 15260 8046 15316
rect 10546 15260 10556 15316
rect 10612 15260 11228 15316
rect 11284 15260 11452 15316
rect 11508 15260 11518 15316
rect 17154 15260 17164 15316
rect 17220 15260 18284 15316
rect 18340 15260 18350 15316
rect 18498 15260 18508 15316
rect 18564 15260 19628 15316
rect 19684 15260 20412 15316
rect 20468 15260 21700 15316
rect 21970 15260 21980 15316
rect 22036 15260 23884 15316
rect 23940 15260 23950 15316
rect 24770 15260 24780 15316
rect 24836 15260 25564 15316
rect 25620 15260 25630 15316
rect 26450 15260 26460 15316
rect 26516 15260 28476 15316
rect 28532 15260 28542 15316
rect 6300 15204 6356 15260
rect 2482 15148 2492 15204
rect 2548 15148 5964 15204
rect 6020 15148 6030 15204
rect 6300 15148 6748 15204
rect 6804 15148 7532 15204
rect 7588 15148 7598 15204
rect 19394 15148 19404 15204
rect 19460 15148 22428 15204
rect 22484 15148 22494 15204
rect 27906 15148 27916 15204
rect 27972 15148 30380 15204
rect 30436 15148 30828 15204
rect 30884 15148 30894 15204
rect 21298 15036 21308 15092
rect 21364 15036 21980 15092
rect 22036 15036 22046 15092
rect 22194 15036 22204 15092
rect 22260 15036 30940 15092
rect 30996 15036 31006 15092
rect 10546 14924 10556 14980
rect 10612 14924 11340 14980
rect 11396 14924 11406 14980
rect 16818 14924 16828 14980
rect 16884 14924 17836 14980
rect 17892 14924 18172 14980
rect 18228 14924 18238 14980
rect 22978 14924 22988 14980
rect 23044 14924 28364 14980
rect 28420 14924 28430 14980
rect 28578 14924 28588 14980
rect 28644 14924 28682 14980
rect 5234 14868 5244 14924
rect 5300 14868 5348 14924
rect 5404 14868 5452 14924
rect 5508 14868 5518 14924
rect 13298 14868 13308 14924
rect 13364 14868 13412 14924
rect 13468 14868 13516 14924
rect 13572 14868 13582 14924
rect 21362 14868 21372 14924
rect 21428 14868 21476 14924
rect 21532 14868 21580 14924
rect 21636 14868 21646 14924
rect 29426 14868 29436 14924
rect 29492 14868 29540 14924
rect 29596 14868 29644 14924
rect 29700 14868 29710 14924
rect 19618 14812 19628 14868
rect 19684 14812 19694 14868
rect 27570 14812 27580 14868
rect 27636 14812 28476 14868
rect 28532 14812 28868 14868
rect 19628 14756 19684 14812
rect 16370 14700 16380 14756
rect 16436 14700 17164 14756
rect 17220 14700 17230 14756
rect 19628 14700 19740 14756
rect 19796 14700 19806 14756
rect 21980 14700 26572 14756
rect 26628 14700 26638 14756
rect 26898 14700 26908 14756
rect 26964 14700 28588 14756
rect 28644 14700 28654 14756
rect 21980 14644 22036 14700
rect 28812 14644 28868 14812
rect 34200 14644 35000 14672
rect 14466 14588 14476 14644
rect 14532 14588 18508 14644
rect 18564 14588 18574 14644
rect 18844 14588 19628 14644
rect 19684 14588 22036 14644
rect 25666 14588 25676 14644
rect 25732 14588 28252 14644
rect 28308 14588 28318 14644
rect 28812 14588 35000 14644
rect 7186 14476 7196 14532
rect 7252 14476 7644 14532
rect 7700 14476 8540 14532
rect 8596 14476 8606 14532
rect 16930 14476 16940 14532
rect 16996 14476 18620 14532
rect 18676 14476 18686 14532
rect 18844 14420 18900 14588
rect 34200 14560 35000 14588
rect 19058 14476 19068 14532
rect 19124 14476 20076 14532
rect 20132 14476 20142 14532
rect 20514 14476 20524 14532
rect 20580 14476 21196 14532
rect 21252 14476 22876 14532
rect 22932 14476 23772 14532
rect 23828 14476 23838 14532
rect 26852 14476 31724 14532
rect 31780 14476 31790 14532
rect 20076 14420 20132 14476
rect 14018 14364 14028 14420
rect 14084 14364 15148 14420
rect 15204 14364 18900 14420
rect 19254 14364 19292 14420
rect 19348 14364 19358 14420
rect 19506 14364 19516 14420
rect 19572 14364 19852 14420
rect 19908 14364 19918 14420
rect 20076 14364 21084 14420
rect 21140 14364 21150 14420
rect 21298 14364 21308 14420
rect 21364 14364 25900 14420
rect 25956 14364 25966 14420
rect 26852 14308 26908 14476
rect 7298 14252 7308 14308
rect 7364 14252 8540 14308
rect 8596 14252 8606 14308
rect 11554 14252 11564 14308
rect 11620 14252 12236 14308
rect 12292 14252 12572 14308
rect 12628 14252 12638 14308
rect 14466 14252 14476 14308
rect 14532 14252 16828 14308
rect 16884 14252 16894 14308
rect 18722 14252 18732 14308
rect 18788 14252 19404 14308
rect 19460 14252 20636 14308
rect 20692 14252 20702 14308
rect 21410 14252 21420 14308
rect 21476 14252 26908 14308
rect 29026 14252 29036 14308
rect 29092 14252 29708 14308
rect 29764 14252 30604 14308
rect 30660 14252 30670 14308
rect 21420 14196 21476 14252
rect 7186 14140 7196 14196
rect 7252 14140 7868 14196
rect 7924 14140 7934 14196
rect 17826 14140 17836 14196
rect 17892 14140 19068 14196
rect 19124 14140 21476 14196
rect 25890 14140 25900 14196
rect 25956 14140 28588 14196
rect 28644 14140 29820 14196
rect 29876 14140 29886 14196
rect 30034 14140 30044 14196
rect 30100 14140 33068 14196
rect 33124 14140 33134 14196
rect 9266 14084 9276 14140
rect 9332 14084 9380 14140
rect 9436 14084 9484 14140
rect 9540 14084 9550 14140
rect 17330 14084 17340 14140
rect 17396 14084 17444 14140
rect 17500 14084 17548 14140
rect 17604 14084 17614 14140
rect 25394 14084 25404 14140
rect 25460 14084 25508 14140
rect 25564 14084 25612 14140
rect 25668 14084 25678 14140
rect 33458 14084 33468 14140
rect 33524 14084 33572 14140
rect 33628 14084 33676 14140
rect 33732 14084 33742 14140
rect 21858 14028 21868 14084
rect 21924 14028 22204 14084
rect 22260 14028 22270 14084
rect 26870 14028 26908 14084
rect 26964 14028 26974 14084
rect 31154 14028 31164 14084
rect 31220 14028 32396 14084
rect 32452 14028 32462 14084
rect 8978 13916 8988 13972
rect 9044 13916 10780 13972
rect 10836 13916 10846 13972
rect 12002 13916 12012 13972
rect 12068 13916 12460 13972
rect 12516 13916 12526 13972
rect 17042 13916 17052 13972
rect 17108 13916 18508 13972
rect 18564 13916 18574 13972
rect 19282 13916 19292 13972
rect 19348 13916 20188 13972
rect 20244 13916 20254 13972
rect 20402 13916 20412 13972
rect 20468 13916 22092 13972
rect 22148 13916 22158 13972
rect 23314 13916 23324 13972
rect 23380 13916 23996 13972
rect 24052 13916 24062 13972
rect 24210 13916 24220 13972
rect 24276 13916 25452 13972
rect 25508 13916 25518 13972
rect 28242 13916 28252 13972
rect 28308 13916 31724 13972
rect 31780 13916 31790 13972
rect 16706 13804 16716 13860
rect 16772 13804 19180 13860
rect 19236 13804 19246 13860
rect 21746 13804 21756 13860
rect 21812 13804 23436 13860
rect 23492 13804 23772 13860
rect 23828 13804 27916 13860
rect 27972 13804 27982 13860
rect 12898 13692 12908 13748
rect 12964 13692 14812 13748
rect 14868 13692 14878 13748
rect 17602 13692 17612 13748
rect 17668 13692 20524 13748
rect 20580 13692 20590 13748
rect 21634 13692 21644 13748
rect 21700 13692 23100 13748
rect 23156 13692 23660 13748
rect 23716 13692 23726 13748
rect 26562 13692 26572 13748
rect 26628 13692 27468 13748
rect 27524 13692 27534 13748
rect 28578 13692 28588 13748
rect 28644 13692 30828 13748
rect 30884 13692 30894 13748
rect 15922 13580 15932 13636
rect 15988 13580 16380 13636
rect 16436 13580 20300 13636
rect 20356 13580 20366 13636
rect 20626 13580 20636 13636
rect 20692 13580 21308 13636
rect 21364 13580 21374 13636
rect 22082 13580 22092 13636
rect 22148 13580 25228 13636
rect 25284 13580 25294 13636
rect 28354 13580 28364 13636
rect 28420 13580 29596 13636
rect 29652 13580 30604 13636
rect 30660 13580 30670 13636
rect 10770 13468 10780 13524
rect 10836 13468 11676 13524
rect 11732 13468 11742 13524
rect 14914 13468 14924 13524
rect 14980 13468 15596 13524
rect 15652 13468 15662 13524
rect 17714 13468 17724 13524
rect 17780 13468 18732 13524
rect 18788 13468 19852 13524
rect 19908 13468 19918 13524
rect 27794 13468 27804 13524
rect 27860 13468 28924 13524
rect 28980 13468 29820 13524
rect 29876 13468 29886 13524
rect 31724 13412 31780 13916
rect 20822 13356 20860 13412
rect 20916 13356 20926 13412
rect 31724 13356 32396 13412
rect 32452 13356 32462 13412
rect 5234 13300 5244 13356
rect 5300 13300 5348 13356
rect 5404 13300 5452 13356
rect 5508 13300 5518 13356
rect 13298 13300 13308 13356
rect 13364 13300 13412 13356
rect 13468 13300 13516 13356
rect 13572 13300 13582 13356
rect 21362 13300 21372 13356
rect 21428 13300 21476 13356
rect 21532 13300 21580 13356
rect 21636 13300 21646 13356
rect 29426 13300 29436 13356
rect 29492 13300 29540 13356
rect 29596 13300 29644 13356
rect 29700 13300 29710 13356
rect 18386 13244 18396 13300
rect 18452 13244 21084 13300
rect 21140 13244 21150 13300
rect 23762 13244 23772 13300
rect 23828 13244 26684 13300
rect 26740 13244 26750 13300
rect 19590 13132 19628 13188
rect 19684 13132 19694 13188
rect 20038 13132 20076 13188
rect 20132 13132 20142 13188
rect 22418 13132 22428 13188
rect 22484 13132 24220 13188
rect 24276 13132 24892 13188
rect 24948 13132 24958 13188
rect 26460 13132 28476 13188
rect 28532 13132 30156 13188
rect 30212 13132 30222 13188
rect 26460 13076 26516 13132
rect 13346 13020 13356 13076
rect 13412 13020 26124 13076
rect 26180 13020 26190 13076
rect 26450 13020 26460 13076
rect 26516 13020 26526 13076
rect 26674 13020 26684 13076
rect 26740 13020 30716 13076
rect 30772 13020 30782 13076
rect 6178 12908 6188 12964
rect 6244 12908 8540 12964
rect 8596 12908 9212 12964
rect 9268 12908 9996 12964
rect 10052 12908 10062 12964
rect 16594 12908 16604 12964
rect 16660 12908 17164 12964
rect 17220 12908 19068 12964
rect 19124 12908 19134 12964
rect 23314 12908 23324 12964
rect 23380 12908 23996 12964
rect 24052 12908 24062 12964
rect 24546 12908 24556 12964
rect 24612 12908 25228 12964
rect 25284 12908 25294 12964
rect 29586 12908 29596 12964
rect 29652 12908 31052 12964
rect 31108 12908 31118 12964
rect 6738 12796 6748 12852
rect 6804 12796 7756 12852
rect 7812 12796 7822 12852
rect 26562 12796 26572 12852
rect 26628 12796 29988 12852
rect 30146 12796 30156 12852
rect 30212 12796 31276 12852
rect 31332 12796 32396 12852
rect 32452 12796 32956 12852
rect 33012 12796 33022 12852
rect 29932 12740 29988 12796
rect 25890 12684 25900 12740
rect 25956 12684 26348 12740
rect 26404 12684 26908 12740
rect 27682 12684 27692 12740
rect 27748 12684 28700 12740
rect 28756 12684 28766 12740
rect 29110 12684 29148 12740
rect 29204 12684 29214 12740
rect 29932 12684 32508 12740
rect 32564 12684 32732 12740
rect 32788 12684 32798 12740
rect 26852 12628 26908 12684
rect 26852 12572 27244 12628
rect 27300 12572 30716 12628
rect 30772 12572 32284 12628
rect 32340 12572 32350 12628
rect 9266 12516 9276 12572
rect 9332 12516 9380 12572
rect 9436 12516 9484 12572
rect 9540 12516 9550 12572
rect 17330 12516 17340 12572
rect 17396 12516 17444 12572
rect 17500 12516 17548 12572
rect 17604 12516 17614 12572
rect 25394 12516 25404 12572
rect 25460 12516 25508 12572
rect 25564 12516 25612 12572
rect 25668 12516 25678 12572
rect 33458 12516 33468 12572
rect 33524 12516 33572 12572
rect 33628 12516 33676 12572
rect 33732 12516 33742 12572
rect 12086 12460 12124 12516
rect 12180 12460 12190 12516
rect 19964 12460 24780 12516
rect 24836 12460 24846 12516
rect 28690 12460 28700 12516
rect 28756 12460 30044 12516
rect 30100 12460 30110 12516
rect 11442 12348 11452 12404
rect 11508 12348 15148 12404
rect 15092 12292 15148 12348
rect 19964 12292 20020 12460
rect 23202 12348 23212 12404
rect 23268 12348 23884 12404
rect 23940 12348 23950 12404
rect 12002 12236 12012 12292
rect 12068 12236 12348 12292
rect 12404 12236 12796 12292
rect 12852 12236 13356 12292
rect 13412 12236 13422 12292
rect 15092 12236 20020 12292
rect 24210 12236 24220 12292
rect 24276 12236 25228 12292
rect 25284 12236 25294 12292
rect 25218 12124 25228 12180
rect 25284 12124 25340 12180
rect 25396 12124 25406 12180
rect 28914 12124 28924 12180
rect 28980 12124 32060 12180
rect 32116 12124 33180 12180
rect 33236 12124 33246 12180
rect 7522 12012 7532 12068
rect 7588 12012 8092 12068
rect 8148 12012 19964 12068
rect 20020 12012 20030 12068
rect 28018 12012 28028 12068
rect 28084 12012 29036 12068
rect 29092 12012 29102 12068
rect 34200 11956 35000 11984
rect 16706 11900 16716 11956
rect 16772 11900 21868 11956
rect 21924 11900 21934 11956
rect 28578 11900 28588 11956
rect 28644 11900 30156 11956
rect 30212 11900 30222 11956
rect 33842 11900 33852 11956
rect 33908 11900 35000 11956
rect 34200 11872 35000 11900
rect 25890 11788 25900 11844
rect 25956 11788 27356 11844
rect 27412 11788 29036 11844
rect 29092 11788 29102 11844
rect 5234 11732 5244 11788
rect 5300 11732 5348 11788
rect 5404 11732 5452 11788
rect 5508 11732 5518 11788
rect 13298 11732 13308 11788
rect 13364 11732 13412 11788
rect 13468 11732 13516 11788
rect 13572 11732 13582 11788
rect 21362 11732 21372 11788
rect 21428 11732 21476 11788
rect 21532 11732 21580 11788
rect 21636 11732 21646 11788
rect 29426 11732 29436 11788
rect 29492 11732 29540 11788
rect 29596 11732 29644 11788
rect 29700 11732 29710 11788
rect 10882 11676 10892 11732
rect 10948 11676 12572 11732
rect 12628 11676 13132 11732
rect 13188 11676 13198 11732
rect 11554 11564 11564 11620
rect 11620 11564 12236 11620
rect 12292 11564 12302 11620
rect 12786 11564 12796 11620
rect 12852 11564 26012 11620
rect 26068 11564 26078 11620
rect 7858 11452 7868 11508
rect 7924 11452 8652 11508
rect 8708 11452 8988 11508
rect 9044 11452 9054 11508
rect 9426 11452 9436 11508
rect 9492 11452 16716 11508
rect 16772 11452 16782 11508
rect 27234 11452 27244 11508
rect 27300 11452 28252 11508
rect 28308 11452 28318 11508
rect 29922 11452 29932 11508
rect 29988 11452 29998 11508
rect 30146 11452 30156 11508
rect 30212 11452 33180 11508
rect 33236 11452 33246 11508
rect 9436 11396 9492 11452
rect 29932 11396 29988 11452
rect 6402 11340 6412 11396
rect 6468 11340 8428 11396
rect 8484 11340 9492 11396
rect 12226 11340 12236 11396
rect 12292 11340 13468 11396
rect 13524 11340 13534 11396
rect 13682 11340 13692 11396
rect 13748 11340 17052 11396
rect 17108 11340 17118 11396
rect 21522 11340 21532 11396
rect 21588 11340 32620 11396
rect 32676 11340 32686 11396
rect 24994 11228 25004 11284
rect 25060 11228 25452 11284
rect 25508 11228 25518 11284
rect 28354 11228 28364 11284
rect 28420 11228 29932 11284
rect 29988 11228 29998 11284
rect 9874 11116 9884 11172
rect 9940 11116 10892 11172
rect 10948 11116 10958 11172
rect 28242 11116 28252 11172
rect 28308 11116 29372 11172
rect 29428 11116 30156 11172
rect 30212 11116 30222 11172
rect 3714 11004 3724 11060
rect 3780 11004 7644 11060
rect 7700 11004 8316 11060
rect 8372 11004 8382 11060
rect 9266 10948 9276 11004
rect 9332 10948 9380 11004
rect 9436 10948 9484 11004
rect 9540 10948 9550 11004
rect 17330 10948 17340 11004
rect 17396 10948 17444 11004
rect 17500 10948 17548 11004
rect 17604 10948 17614 11004
rect 25394 10948 25404 11004
rect 25460 10948 25508 11004
rect 25564 10948 25612 11004
rect 25668 10948 25678 11004
rect 33458 10948 33468 11004
rect 33524 10948 33572 11004
rect 33628 10948 33676 11004
rect 33732 10948 33742 11004
rect 4498 10780 4508 10836
rect 4564 10780 5964 10836
rect 6020 10780 6412 10836
rect 6468 10780 6478 10836
rect 8194 10780 8204 10836
rect 8260 10780 8652 10836
rect 8708 10780 10668 10836
rect 10724 10780 10734 10836
rect 19730 10780 19740 10836
rect 19796 10780 21308 10836
rect 21364 10780 22876 10836
rect 22932 10780 22942 10836
rect 28802 10780 28812 10836
rect 28868 10780 32956 10836
rect 33012 10780 33022 10836
rect 9650 10668 9660 10724
rect 9716 10668 24556 10724
rect 24612 10668 24622 10724
rect 25554 10668 25564 10724
rect 25620 10668 26460 10724
rect 26516 10668 26526 10724
rect 2818 10556 2828 10612
rect 2884 10556 3724 10612
rect 3780 10556 3790 10612
rect 14130 10556 14140 10612
rect 14196 10556 15708 10612
rect 15764 10556 17612 10612
rect 17668 10556 20300 10612
rect 20356 10556 20972 10612
rect 21028 10556 21038 10612
rect 24658 10556 24668 10612
rect 24724 10556 25452 10612
rect 25508 10556 26348 10612
rect 26404 10556 26414 10612
rect 26562 10556 26572 10612
rect 26628 10556 27132 10612
rect 27188 10556 27198 10612
rect 27458 10556 27468 10612
rect 27524 10556 31836 10612
rect 31892 10556 31902 10612
rect 9986 10444 9996 10500
rect 10052 10444 10780 10500
rect 10836 10444 10846 10500
rect 14242 10444 14252 10500
rect 14308 10444 15932 10500
rect 15988 10444 15998 10500
rect 22530 10444 22540 10500
rect 22596 10444 23324 10500
rect 23380 10444 23390 10500
rect 23874 10444 23884 10500
rect 23940 10444 25340 10500
rect 25396 10444 25406 10500
rect 26002 10444 26012 10500
rect 26068 10444 29260 10500
rect 29316 10444 31724 10500
rect 31780 10444 33068 10500
rect 33124 10444 33134 10500
rect 5058 10332 5068 10388
rect 5124 10332 5404 10388
rect 5460 10332 5470 10388
rect 22978 10332 22988 10388
rect 23044 10332 28700 10388
rect 28756 10332 28766 10388
rect 21858 10220 21868 10276
rect 21924 10220 22316 10276
rect 22372 10220 25004 10276
rect 25060 10220 25070 10276
rect 5234 10164 5244 10220
rect 5300 10164 5348 10220
rect 5404 10164 5452 10220
rect 5508 10164 5518 10220
rect 13298 10164 13308 10220
rect 13364 10164 13412 10220
rect 13468 10164 13516 10220
rect 13572 10164 13582 10220
rect 21362 10164 21372 10220
rect 21428 10164 21476 10220
rect 21532 10164 21580 10220
rect 21636 10164 21646 10220
rect 29426 10164 29436 10220
rect 29492 10164 29540 10220
rect 29596 10164 29644 10220
rect 29700 10164 29710 10220
rect 14354 10108 14364 10164
rect 14420 10108 15148 10164
rect 15204 10108 15214 10164
rect 22754 10108 22764 10164
rect 22820 10108 24892 10164
rect 24948 10108 24958 10164
rect 30482 10108 30492 10164
rect 30548 10108 31052 10164
rect 31108 10108 31118 10164
rect 4834 9996 4844 10052
rect 4900 9996 5516 10052
rect 5572 9996 7196 10052
rect 7252 9996 7262 10052
rect 13794 9996 13804 10052
rect 13860 9996 20636 10052
rect 20692 9996 20702 10052
rect 25218 9996 25228 10052
rect 25284 9996 27020 10052
rect 27076 9996 29148 10052
rect 29204 9996 29214 10052
rect 13010 9884 13020 9940
rect 13076 9884 13916 9940
rect 13972 9884 13982 9940
rect 15092 9884 22204 9940
rect 22260 9884 22540 9940
rect 22596 9884 22606 9940
rect 23538 9884 23548 9940
rect 23604 9884 25452 9940
rect 25508 9884 25518 9940
rect 26674 9884 26684 9940
rect 26740 9884 27132 9940
rect 27188 9884 27198 9940
rect 15092 9828 15148 9884
rect 25452 9828 25508 9884
rect 5702 9772 5740 9828
rect 5796 9772 6412 9828
rect 6468 9772 6478 9828
rect 7074 9772 7084 9828
rect 7140 9772 8764 9828
rect 8820 9772 8830 9828
rect 13122 9772 13132 9828
rect 13188 9772 15148 9828
rect 17938 9772 17948 9828
rect 18004 9772 19292 9828
rect 19348 9772 19964 9828
rect 20020 9772 20030 9828
rect 20290 9772 20300 9828
rect 20356 9772 21868 9828
rect 21924 9772 24444 9828
rect 24500 9772 24510 9828
rect 25452 9772 28140 9828
rect 28196 9772 28206 9828
rect 3266 9660 3276 9716
rect 3332 9660 6748 9716
rect 6804 9660 7420 9716
rect 7476 9660 7486 9716
rect 8306 9660 8316 9716
rect 8372 9660 8652 9716
rect 8708 9660 8718 9716
rect 13794 9660 13804 9716
rect 13860 9660 18172 9716
rect 18228 9660 18238 9716
rect 23314 9660 23324 9716
rect 23380 9660 24332 9716
rect 24388 9660 24398 9716
rect 25218 9660 25228 9716
rect 25284 9660 29260 9716
rect 29316 9660 29326 9716
rect 4050 9548 4060 9604
rect 4116 9548 4956 9604
rect 5012 9548 6076 9604
rect 6132 9548 7532 9604
rect 7588 9548 7598 9604
rect 7970 9548 7980 9604
rect 8036 9548 9100 9604
rect 9156 9548 9660 9604
rect 9716 9548 9726 9604
rect 11890 9548 11900 9604
rect 11956 9548 14812 9604
rect 14868 9548 14878 9604
rect 15586 9548 15596 9604
rect 15652 9548 17948 9604
rect 18004 9548 18014 9604
rect 20626 9548 20636 9604
rect 20692 9548 25340 9604
rect 25396 9548 25406 9604
rect 25666 9548 25676 9604
rect 25732 9548 26572 9604
rect 26628 9548 26638 9604
rect 26852 9548 27468 9604
rect 27524 9548 29596 9604
rect 29652 9548 29662 9604
rect 10434 9436 10444 9492
rect 10500 9436 10892 9492
rect 10948 9436 10958 9492
rect 9266 9380 9276 9436
rect 9332 9380 9380 9436
rect 9436 9380 9484 9436
rect 9540 9380 9550 9436
rect 7298 9324 7308 9380
rect 7364 9324 7756 9380
rect 7812 9324 7822 9380
rect 14812 9268 14868 9548
rect 26852 9492 26908 9548
rect 25890 9436 25900 9492
rect 25956 9436 26908 9492
rect 31826 9436 31836 9492
rect 31892 9436 32732 9492
rect 32788 9436 32798 9492
rect 17330 9380 17340 9436
rect 17396 9380 17444 9436
rect 17500 9380 17548 9436
rect 17604 9380 17614 9436
rect 25394 9380 25404 9436
rect 25460 9380 25508 9436
rect 25564 9380 25612 9436
rect 25668 9380 25678 9436
rect 33458 9380 33468 9436
rect 33524 9380 33572 9436
rect 33628 9380 33676 9436
rect 33732 9380 33742 9436
rect 34200 9268 35000 9296
rect 14812 9212 16268 9268
rect 16324 9212 17500 9268
rect 17556 9212 17566 9268
rect 19058 9212 19068 9268
rect 19124 9212 22316 9268
rect 22372 9212 22382 9268
rect 23762 9212 23772 9268
rect 23828 9212 24332 9268
rect 24388 9212 25564 9268
rect 25620 9212 26908 9268
rect 26964 9212 26974 9268
rect 28578 9212 28588 9268
rect 28644 9212 29260 9268
rect 29316 9212 29326 9268
rect 30258 9212 30268 9268
rect 30324 9212 33292 9268
rect 33348 9212 33358 9268
rect 33516 9212 35000 9268
rect 33516 9156 33572 9212
rect 34200 9184 35000 9212
rect 4610 9100 4620 9156
rect 4676 9100 6188 9156
rect 6244 9100 6254 9156
rect 10210 9100 10220 9156
rect 10276 9100 11564 9156
rect 11620 9100 11630 9156
rect 12226 9100 12236 9156
rect 12292 9100 13692 9156
rect 13748 9100 15148 9156
rect 16146 9100 16156 9156
rect 16212 9100 16828 9156
rect 16884 9100 16894 9156
rect 24546 9100 24556 9156
rect 24612 9100 26124 9156
rect 26180 9100 28028 9156
rect 28084 9100 29148 9156
rect 29204 9100 29214 9156
rect 32498 9100 32508 9156
rect 32564 9100 33572 9156
rect 15092 9044 15148 9100
rect 10882 8988 10892 9044
rect 10948 8988 11340 9044
rect 11396 8988 12572 9044
rect 12628 8988 12908 9044
rect 12964 8988 12974 9044
rect 15092 8988 16716 9044
rect 16772 8988 16782 9044
rect 17714 8988 17724 9044
rect 17780 8988 19628 9044
rect 19684 8988 19694 9044
rect 26852 8988 30940 9044
rect 30996 8988 31006 9044
rect 3490 8876 3500 8932
rect 3556 8876 5068 8932
rect 5124 8876 5134 8932
rect 9762 8876 9772 8932
rect 9828 8876 11788 8932
rect 11844 8876 12460 8932
rect 12516 8876 12526 8932
rect 15810 8876 15820 8932
rect 15876 8876 16604 8932
rect 16660 8876 16670 8932
rect 22530 8876 22540 8932
rect 22596 8876 24444 8932
rect 24500 8876 24510 8932
rect 26852 8820 26908 8988
rect 1698 8764 1708 8820
rect 1764 8764 4284 8820
rect 4340 8764 4350 8820
rect 4610 8764 4620 8820
rect 4676 8764 5180 8820
rect 5236 8764 5246 8820
rect 10770 8764 10780 8820
rect 10836 8764 23212 8820
rect 23268 8764 26908 8820
rect 4620 8708 4676 8764
rect 3938 8652 3948 8708
rect 4004 8652 4676 8708
rect 25106 8652 25116 8708
rect 25172 8652 25340 8708
rect 25396 8652 25406 8708
rect 5234 8596 5244 8652
rect 5300 8596 5348 8652
rect 5404 8596 5452 8652
rect 5508 8596 5518 8652
rect 13298 8596 13308 8652
rect 13364 8596 13412 8652
rect 13468 8596 13516 8652
rect 13572 8596 13582 8652
rect 21362 8596 21372 8652
rect 21428 8596 21476 8652
rect 21532 8596 21580 8652
rect 21636 8596 21646 8652
rect 29426 8596 29436 8652
rect 29492 8596 29540 8652
rect 29596 8596 29644 8652
rect 29700 8596 29710 8652
rect 31602 8540 31612 8596
rect 31668 8540 32396 8596
rect 32452 8540 32462 8596
rect 11554 8428 11564 8484
rect 11620 8428 12012 8484
rect 12068 8428 12078 8484
rect 16706 8428 16716 8484
rect 16772 8428 17836 8484
rect 17892 8428 17902 8484
rect 18050 8428 18060 8484
rect 18116 8428 23436 8484
rect 23492 8428 23502 8484
rect 25564 8428 28420 8484
rect 29474 8428 29484 8484
rect 29540 8428 31724 8484
rect 31780 8428 31790 8484
rect 25564 8372 25620 8428
rect 28364 8372 28420 8428
rect 2146 8316 2156 8372
rect 2212 8316 2716 8372
rect 2772 8316 2782 8372
rect 6178 8316 6188 8372
rect 6244 8316 7868 8372
rect 7924 8316 7934 8372
rect 22306 8316 22316 8372
rect 22372 8316 25620 8372
rect 25778 8316 25788 8372
rect 25844 8316 26908 8372
rect 28364 8316 33852 8372
rect 33908 8316 33918 8372
rect 26852 8260 26908 8316
rect 1810 8204 1820 8260
rect 1876 8204 4508 8260
rect 4564 8204 4574 8260
rect 11666 8204 11676 8260
rect 11732 8204 12460 8260
rect 12516 8204 14924 8260
rect 14980 8204 19180 8260
rect 19236 8204 19740 8260
rect 19796 8204 22092 8260
rect 22148 8204 26236 8260
rect 26292 8204 26302 8260
rect 26852 8204 28140 8260
rect 28196 8204 28206 8260
rect 3154 8092 3164 8148
rect 3220 8092 5740 8148
rect 5796 8092 5806 8148
rect 19282 8092 19292 8148
rect 19348 8092 20300 8148
rect 20356 8092 20366 8148
rect 21858 8092 21868 8148
rect 21924 8092 32508 8148
rect 32564 8092 32574 8148
rect 4386 7980 4396 8036
rect 4452 7980 6748 8036
rect 6804 7980 6814 8036
rect 19842 7980 19852 8036
rect 19908 7980 23996 8036
rect 24052 7980 24062 8036
rect 24322 7980 24332 8036
rect 24388 7980 24668 8036
rect 24724 7980 24734 8036
rect 26786 7980 26796 8036
rect 26852 7980 28588 8036
rect 28644 7980 28654 8036
rect 2034 7868 2044 7924
rect 2100 7868 3836 7924
rect 3892 7868 3902 7924
rect 5170 7868 5180 7924
rect 5236 7868 9156 7924
rect 19506 7868 19516 7924
rect 19572 7868 19964 7924
rect 20020 7868 20030 7924
rect 32050 7868 32060 7924
rect 32116 7868 32396 7924
rect 32452 7868 32462 7924
rect 5506 7756 5516 7812
rect 5572 7756 5852 7812
rect 5908 7756 5918 7812
rect 9100 7700 9156 7868
rect 9266 7812 9276 7868
rect 9332 7812 9380 7868
rect 9436 7812 9484 7868
rect 9540 7812 9550 7868
rect 17330 7812 17340 7868
rect 17396 7812 17444 7868
rect 17500 7812 17548 7868
rect 17604 7812 17614 7868
rect 25394 7812 25404 7868
rect 25460 7812 25508 7868
rect 25564 7812 25612 7868
rect 25668 7812 25678 7868
rect 33458 7812 33468 7868
rect 33524 7812 33572 7868
rect 33628 7812 33676 7868
rect 33732 7812 33742 7868
rect 18386 7756 18396 7812
rect 18452 7756 21644 7812
rect 21700 7756 21756 7812
rect 21812 7756 21822 7812
rect 23286 7756 23324 7812
rect 23380 7756 23390 7812
rect 2146 7644 2156 7700
rect 2212 7644 4172 7700
rect 4228 7644 4238 7700
rect 4946 7644 4956 7700
rect 5012 7644 5964 7700
rect 6020 7644 6030 7700
rect 9100 7644 9212 7700
rect 9268 7644 9996 7700
rect 10052 7644 10062 7700
rect 12338 7644 12348 7700
rect 12404 7644 13692 7700
rect 13748 7644 13758 7700
rect 16594 7644 16604 7700
rect 16660 7644 17612 7700
rect 17668 7644 17678 7700
rect 20626 7644 20636 7700
rect 20692 7644 25116 7700
rect 25172 7644 26796 7700
rect 26852 7644 26862 7700
rect 28588 7644 29148 7700
rect 29204 7644 29214 7700
rect 30258 7644 30268 7700
rect 30324 7644 31052 7700
rect 31108 7644 31118 7700
rect 28588 7588 28644 7644
rect 2482 7532 2492 7588
rect 2548 7532 6300 7588
rect 6356 7532 6366 7588
rect 16482 7532 16492 7588
rect 16548 7532 16716 7588
rect 16772 7532 19292 7588
rect 19348 7532 20076 7588
rect 20132 7532 20142 7588
rect 21746 7532 21756 7588
rect 21812 7532 22092 7588
rect 22148 7532 23548 7588
rect 23604 7532 23614 7588
rect 26646 7532 26684 7588
rect 26740 7532 26750 7588
rect 27010 7532 27020 7588
rect 27076 7532 28588 7588
rect 28644 7532 28654 7588
rect 28914 7532 28924 7588
rect 28980 7532 31948 7588
rect 32004 7532 32014 7588
rect 4274 7420 4284 7476
rect 4340 7420 6076 7476
rect 6132 7420 6142 7476
rect 6738 7420 6748 7476
rect 6804 7420 8316 7476
rect 8372 7420 8382 7476
rect 17378 7420 17388 7476
rect 17444 7420 18508 7476
rect 18564 7420 19180 7476
rect 19236 7420 19246 7476
rect 22754 7420 22764 7476
rect 22820 7420 23100 7476
rect 23156 7420 23166 7476
rect 23426 7420 23436 7476
rect 23492 7420 24556 7476
rect 24612 7420 24622 7476
rect 24770 7420 24780 7476
rect 24836 7420 26908 7476
rect 26964 7420 26974 7476
rect 27122 7420 27132 7476
rect 27188 7420 27692 7476
rect 27748 7420 29148 7476
rect 29204 7420 29214 7476
rect 30482 7420 30492 7476
rect 30548 7420 32172 7476
rect 32228 7420 32238 7476
rect 33170 7420 33180 7476
rect 33236 7420 33852 7476
rect 33908 7420 33918 7476
rect 5954 7308 5964 7364
rect 6020 7308 6972 7364
rect 7028 7308 7038 7364
rect 10770 7308 10780 7364
rect 10836 7308 12124 7364
rect 12180 7308 12190 7364
rect 13346 7308 13356 7364
rect 13412 7308 19404 7364
rect 19460 7308 19470 7364
rect 23650 7308 23660 7364
rect 23716 7308 24444 7364
rect 24500 7308 24510 7364
rect 24658 7308 24668 7364
rect 24724 7308 25228 7364
rect 25284 7308 25294 7364
rect 31154 7308 31164 7364
rect 31220 7308 31500 7364
rect 31556 7308 31566 7364
rect 2594 7196 2604 7252
rect 2660 7196 4396 7252
rect 4452 7196 4462 7252
rect 4834 7196 4844 7252
rect 4900 7196 8428 7252
rect 8484 7196 8494 7252
rect 16930 7196 16940 7252
rect 16996 7196 17612 7252
rect 17668 7196 17678 7252
rect 24322 7084 24332 7140
rect 24388 7084 27692 7140
rect 27748 7084 27758 7140
rect 5234 7028 5244 7084
rect 5300 7028 5348 7084
rect 5404 7028 5452 7084
rect 5508 7028 5518 7084
rect 13298 7028 13308 7084
rect 13364 7028 13412 7084
rect 13468 7028 13516 7084
rect 13572 7028 13582 7084
rect 21362 7028 21372 7084
rect 21428 7028 21476 7084
rect 21532 7028 21580 7084
rect 21636 7028 21646 7084
rect 29426 7028 29436 7084
rect 29492 7028 29540 7084
rect 29596 7028 29644 7084
rect 29700 7028 29710 7084
rect 5852 6972 7420 7028
rect 7476 6972 7486 7028
rect 27010 6972 27020 7028
rect 27076 6972 27692 7028
rect 27748 6972 28252 7028
rect 28308 6972 28318 7028
rect 5852 6916 5908 6972
rect 3826 6860 3836 6916
rect 3892 6860 5908 6916
rect 6514 6860 6524 6916
rect 6580 6860 9436 6916
rect 9492 6860 9502 6916
rect 9650 6860 9660 6916
rect 9716 6860 12124 6916
rect 12180 6860 12190 6916
rect 24182 6860 24220 6916
rect 24276 6860 24286 6916
rect 25890 6860 25900 6916
rect 25956 6860 26460 6916
rect 26516 6860 26526 6916
rect 27010 6860 27020 6916
rect 27076 6860 27086 6916
rect 28690 6860 28700 6916
rect 28756 6860 30604 6916
rect 30660 6860 30670 6916
rect 5506 6748 5516 6804
rect 5572 6748 6860 6804
rect 6916 6748 6926 6804
rect 7410 6748 7420 6804
rect 7476 6748 8764 6804
rect 8820 6748 8830 6804
rect 12124 6748 12572 6804
rect 12628 6748 13020 6804
rect 13076 6748 13086 6804
rect 20738 6748 20748 6804
rect 20804 6748 22540 6804
rect 22596 6748 22606 6804
rect 24546 6748 24556 6804
rect 24612 6748 26796 6804
rect 26852 6748 26862 6804
rect 12124 6692 12180 6748
rect 27020 6692 27076 6860
rect 28130 6748 28140 6804
rect 28196 6748 30716 6804
rect 30772 6748 30782 6804
rect 3332 6636 5852 6692
rect 5908 6636 5918 6692
rect 6402 6636 6412 6692
rect 6468 6636 9100 6692
rect 9156 6636 9660 6692
rect 9716 6636 9726 6692
rect 10994 6636 11004 6692
rect 11060 6636 11340 6692
rect 11396 6636 12180 6692
rect 12338 6636 12348 6692
rect 12404 6636 13580 6692
rect 13636 6636 13646 6692
rect 15026 6636 15036 6692
rect 15092 6636 17052 6692
rect 17108 6636 17118 6692
rect 22642 6636 22652 6692
rect 22708 6636 22718 6692
rect 25666 6636 25676 6692
rect 25732 6636 26348 6692
rect 26404 6636 27076 6692
rect 3332 6580 3388 6636
rect 22652 6580 22708 6636
rect 34200 6580 35000 6608
rect 2370 6524 2380 6580
rect 2436 6524 3388 6580
rect 4834 6524 4844 6580
rect 4900 6524 5740 6580
rect 5796 6524 5806 6580
rect 9538 6524 9548 6580
rect 9604 6524 10332 6580
rect 10388 6524 11788 6580
rect 11844 6524 11854 6580
rect 12012 6524 12796 6580
rect 12852 6524 12862 6580
rect 14018 6524 14028 6580
rect 14084 6524 16604 6580
rect 16660 6524 16670 6580
rect 22652 6524 29820 6580
rect 29876 6524 35000 6580
rect 12012 6468 12068 6524
rect 34200 6496 35000 6524
rect 3826 6412 3836 6468
rect 3892 6412 5740 6468
rect 5796 6412 5806 6468
rect 9874 6412 9884 6468
rect 9940 6412 12068 6468
rect 12562 6412 12572 6468
rect 12628 6412 14140 6468
rect 14196 6412 14206 6468
rect 17266 6412 17276 6468
rect 17332 6412 18452 6468
rect 18610 6412 18620 6468
rect 18676 6412 21756 6468
rect 21812 6412 21822 6468
rect 21970 6412 21980 6468
rect 22036 6412 22764 6468
rect 22820 6412 24780 6468
rect 24836 6412 25340 6468
rect 25396 6412 25406 6468
rect 25554 6412 25564 6468
rect 25620 6412 26684 6468
rect 26740 6412 30156 6468
rect 30212 6412 31164 6468
rect 31220 6412 31230 6468
rect 18396 6356 18452 6412
rect 9650 6300 9660 6356
rect 9716 6300 10220 6356
rect 10276 6300 10286 6356
rect 11890 6300 11900 6356
rect 11956 6300 13692 6356
rect 13748 6300 13758 6356
rect 18396 6300 22876 6356
rect 22932 6300 22942 6356
rect 23538 6300 23548 6356
rect 23604 6300 24220 6356
rect 24276 6300 24286 6356
rect 24406 6300 24444 6356
rect 24500 6300 24510 6356
rect 27570 6300 27580 6356
rect 27636 6300 28588 6356
rect 28644 6300 28654 6356
rect 29586 6300 29596 6356
rect 29652 6300 31948 6356
rect 32004 6300 32014 6356
rect 9266 6244 9276 6300
rect 9332 6244 9380 6300
rect 9436 6244 9484 6300
rect 9540 6244 9550 6300
rect 17330 6244 17340 6300
rect 17396 6244 17444 6300
rect 17500 6244 17548 6300
rect 17604 6244 17614 6300
rect 25394 6244 25404 6300
rect 25460 6244 25508 6300
rect 25564 6244 25612 6300
rect 25668 6244 25678 6300
rect 33458 6244 33468 6300
rect 33524 6244 33572 6300
rect 33628 6244 33676 6300
rect 33732 6244 33742 6300
rect 5282 6188 5292 6244
rect 5348 6188 8092 6244
rect 8148 6188 8158 6244
rect 12786 6188 12796 6244
rect 12852 6188 14252 6244
rect 14308 6188 14318 6244
rect 22754 6188 22764 6244
rect 22820 6188 24108 6244
rect 24164 6188 24174 6244
rect 24882 6188 24892 6244
rect 24948 6188 25116 6244
rect 25172 6188 25182 6244
rect 28466 6188 28476 6244
rect 28532 6188 29148 6244
rect 29204 6188 33068 6244
rect 33124 6188 33134 6244
rect 5170 6076 5180 6132
rect 5236 6076 5740 6132
rect 5796 6076 5806 6132
rect 11900 6076 13244 6132
rect 13300 6076 13310 6132
rect 22194 6076 22204 6132
rect 22260 6076 23436 6132
rect 23492 6076 24332 6132
rect 24388 6076 26012 6132
rect 26068 6076 26078 6132
rect 26338 6076 26348 6132
rect 26404 6076 26796 6132
rect 26852 6076 26862 6132
rect 28242 6076 28252 6132
rect 28308 6076 30044 6132
rect 30100 6076 30110 6132
rect 30482 6076 30492 6132
rect 30548 6076 31724 6132
rect 31780 6076 31790 6132
rect 11900 6020 11956 6076
rect 5030 5964 5068 6020
rect 5124 5964 5134 6020
rect 9762 5964 9772 6020
rect 9828 5964 11900 6020
rect 11956 5964 11966 6020
rect 13122 5964 13132 6020
rect 13188 5964 17276 6020
rect 17332 5964 17342 6020
rect 19730 5964 19740 6020
rect 19796 5964 22652 6020
rect 22708 5964 22718 6020
rect 29810 5964 29820 6020
rect 29876 5964 30828 6020
rect 30884 5964 30894 6020
rect 14354 5852 14364 5908
rect 14420 5852 17500 5908
rect 17556 5852 17566 5908
rect 19058 5852 19068 5908
rect 19124 5852 20748 5908
rect 20804 5852 20814 5908
rect 23090 5852 23100 5908
rect 23156 5852 23548 5908
rect 23604 5852 24780 5908
rect 24836 5852 24846 5908
rect 25330 5852 25340 5908
rect 25396 5852 25676 5908
rect 25732 5852 25742 5908
rect 26338 5852 26348 5908
rect 26404 5852 27692 5908
rect 27748 5852 27758 5908
rect 28802 5852 28812 5908
rect 28868 5852 30380 5908
rect 30436 5852 30446 5908
rect 16930 5740 16940 5796
rect 16996 5740 19292 5796
rect 19348 5740 19358 5796
rect 21858 5740 21868 5796
rect 21924 5740 23324 5796
rect 23380 5740 23390 5796
rect 30594 5740 30604 5796
rect 30660 5740 33180 5796
rect 33236 5740 33246 5796
rect 3826 5628 3836 5684
rect 3892 5628 6300 5684
rect 6356 5628 6366 5684
rect 9762 5628 9772 5684
rect 9828 5628 12124 5684
rect 12180 5628 12190 5684
rect 12450 5628 12460 5684
rect 12516 5628 13580 5684
rect 13636 5628 15820 5684
rect 15876 5628 15886 5684
rect 16594 5628 16604 5684
rect 16660 5628 17724 5684
rect 17780 5628 18396 5684
rect 18452 5628 18462 5684
rect 21746 5628 21756 5684
rect 21812 5628 23660 5684
rect 23716 5628 23726 5684
rect 28018 5628 28028 5684
rect 28084 5628 29372 5684
rect 29428 5628 32284 5684
rect 32340 5628 32350 5684
rect 16370 5516 16380 5572
rect 16436 5516 17948 5572
rect 18004 5516 18014 5572
rect 23314 5516 23324 5572
rect 23380 5516 24108 5572
rect 24164 5516 24174 5572
rect 5234 5460 5244 5516
rect 5300 5460 5348 5516
rect 5404 5460 5452 5516
rect 5508 5460 5518 5516
rect 13298 5460 13308 5516
rect 13364 5460 13412 5516
rect 13468 5460 13516 5516
rect 13572 5460 13582 5516
rect 21362 5460 21372 5516
rect 21428 5460 21476 5516
rect 21532 5460 21580 5516
rect 21636 5460 21646 5516
rect 29426 5460 29436 5516
rect 29492 5460 29540 5516
rect 29596 5460 29644 5516
rect 29700 5460 29710 5516
rect 1698 5404 1708 5460
rect 1764 5404 2044 5460
rect 2100 5404 2380 5460
rect 2436 5404 2446 5460
rect 18834 5404 18844 5460
rect 18900 5404 19740 5460
rect 19796 5404 19806 5460
rect 24210 5404 24220 5460
rect 24276 5404 24286 5460
rect 26450 5404 26460 5460
rect 26516 5404 26908 5460
rect 26964 5404 26974 5460
rect 24220 5348 24276 5404
rect 2258 5292 2268 5348
rect 2324 5292 5628 5348
rect 5684 5292 5694 5348
rect 24220 5292 26348 5348
rect 26404 5292 26796 5348
rect 26852 5292 26862 5348
rect 27346 5292 27356 5348
rect 27412 5292 28364 5348
rect 28420 5292 28430 5348
rect 28578 5292 28588 5348
rect 28644 5292 32844 5348
rect 32900 5292 32910 5348
rect 5954 5180 5964 5236
rect 6020 5180 6412 5236
rect 6468 5180 6478 5236
rect 9762 5180 9772 5236
rect 9828 5180 10556 5236
rect 10612 5180 10622 5236
rect 14802 5180 14812 5236
rect 14868 5180 15148 5236
rect 15204 5180 16380 5236
rect 16436 5180 16446 5236
rect 21298 5180 21308 5236
rect 21364 5180 22540 5236
rect 22596 5180 22606 5236
rect 22764 5180 24556 5236
rect 24612 5180 24622 5236
rect 22764 5124 22820 5180
rect 6066 5068 6076 5124
rect 6132 5068 6860 5124
rect 6916 5068 6926 5124
rect 11666 5068 11676 5124
rect 11732 5068 12348 5124
rect 12404 5068 12414 5124
rect 14578 5068 14588 5124
rect 14644 5068 15372 5124
rect 15428 5068 15438 5124
rect 18386 5068 18396 5124
rect 18452 5068 20300 5124
rect 20356 5068 20366 5124
rect 21634 5068 21644 5124
rect 21700 5068 22820 5124
rect 23202 5068 23212 5124
rect 23268 5068 24332 5124
rect 24388 5068 24398 5124
rect 24770 5068 24780 5124
rect 24836 5068 25340 5124
rect 25396 5068 26684 5124
rect 26740 5068 26750 5124
rect 28018 5068 28028 5124
rect 28084 5068 29036 5124
rect 29092 5068 29102 5124
rect 31938 5068 31948 5124
rect 32004 5068 32396 5124
rect 32452 5068 32462 5124
rect 19404 5012 19460 5068
rect 1922 4956 1932 5012
rect 1988 4956 6524 5012
rect 6580 4956 6590 5012
rect 19282 4956 19292 5012
rect 19348 4956 19460 5012
rect 23986 4956 23996 5012
rect 24052 4956 25620 5012
rect 25564 4900 25620 4956
rect 17154 4844 17164 4900
rect 17220 4844 18732 4900
rect 18788 4844 19740 4900
rect 19796 4844 19806 4900
rect 25554 4844 25564 4900
rect 25620 4844 25630 4900
rect 9266 4676 9276 4732
rect 9332 4676 9380 4732
rect 9436 4676 9484 4732
rect 9540 4676 9550 4732
rect 17330 4676 17340 4732
rect 17396 4676 17444 4732
rect 17500 4676 17548 4732
rect 17604 4676 17614 4732
rect 25394 4676 25404 4732
rect 25460 4676 25508 4732
rect 25564 4676 25612 4732
rect 25668 4676 25678 4732
rect 33458 4676 33468 4732
rect 33524 4676 33572 4732
rect 33628 4676 33676 4732
rect 33732 4676 33742 4732
rect 24406 4508 24444 4564
rect 24500 4508 24510 4564
rect 25330 4508 25340 4564
rect 25396 4508 26684 4564
rect 26740 4508 28644 4564
rect 24994 4396 25004 4452
rect 25060 4396 28420 4452
rect 7858 4284 7868 4340
rect 7924 4284 8428 4340
rect 8484 4284 8494 4340
rect 15586 4284 15596 4340
rect 15652 4284 17388 4340
rect 17444 4284 17454 4340
rect 20850 4284 20860 4340
rect 20916 4284 25564 4340
rect 25620 4284 25630 4340
rect 26338 4284 26348 4340
rect 26404 4284 26908 4340
rect 19170 4172 19180 4228
rect 19236 4172 20300 4228
rect 20356 4172 21532 4228
rect 21588 4172 21598 4228
rect 24658 4172 24668 4228
rect 24724 4172 26236 4228
rect 26292 4172 26302 4228
rect 26852 4116 26908 4284
rect 28364 4228 28420 4396
rect 28588 4340 28644 4508
rect 31714 4396 31724 4452
rect 31780 4396 32172 4452
rect 32228 4396 32238 4452
rect 28578 4284 28588 4340
rect 28644 4284 28654 4340
rect 28364 4172 30268 4228
rect 30324 4172 30334 4228
rect 31266 4172 31276 4228
rect 31332 4172 33180 4228
rect 33236 4172 33246 4228
rect 19730 4060 19740 4116
rect 19796 4060 20748 4116
rect 20804 4060 20814 4116
rect 26852 4060 33236 4116
rect 33180 4004 33236 4060
rect 33170 3948 33180 4004
rect 33236 3948 33246 4004
rect 5234 3892 5244 3948
rect 5300 3892 5348 3948
rect 5404 3892 5452 3948
rect 5508 3892 5518 3948
rect 13298 3892 13308 3948
rect 13364 3892 13412 3948
rect 13468 3892 13516 3948
rect 13572 3892 13582 3948
rect 21362 3892 21372 3948
rect 21428 3892 21476 3948
rect 21532 3892 21580 3948
rect 21636 3892 21646 3948
rect 29426 3892 29436 3948
rect 29492 3892 29540 3948
rect 29596 3892 29644 3948
rect 29700 3892 29710 3948
rect 33180 3892 33236 3948
rect 34200 3892 35000 3920
rect 22082 3836 22092 3892
rect 22148 3836 29316 3892
rect 33180 3836 35000 3892
rect 29260 3780 29316 3836
rect 34200 3808 35000 3836
rect 21074 3724 21084 3780
rect 21140 3724 27580 3780
rect 27636 3724 28588 3780
rect 28644 3724 28654 3780
rect 29260 3724 32284 3780
rect 32340 3724 32350 3780
rect 19842 3612 19852 3668
rect 19908 3612 21868 3668
rect 21924 3612 21934 3668
rect 26562 3612 26572 3668
rect 26628 3612 30716 3668
rect 30772 3612 30782 3668
rect 914 3500 924 3556
rect 980 3500 3276 3556
rect 3332 3500 3342 3556
rect 24770 3500 24780 3556
rect 24836 3500 27020 3556
rect 27076 3500 27086 3556
rect 27682 3500 27692 3556
rect 27748 3500 29148 3556
rect 29204 3500 29596 3556
rect 29652 3500 29662 3556
rect 30258 3500 30268 3556
rect 30324 3500 33852 3556
rect 33908 3500 33918 3556
rect 2034 3388 2044 3444
rect 2100 3388 7868 3444
rect 7924 3388 7934 3444
rect 12674 3388 12684 3444
rect 12740 3388 13356 3444
rect 13412 3388 13804 3444
rect 13860 3388 13870 3444
rect 22866 3388 22876 3444
rect 22932 3388 23996 3444
rect 24052 3388 25900 3444
rect 25956 3388 25966 3444
rect 26338 3388 26348 3444
rect 26404 3388 27468 3444
rect 27524 3388 27534 3444
rect 28690 3388 28700 3444
rect 28756 3388 29372 3444
rect 29428 3388 29438 3444
rect 2146 3276 2156 3332
rect 2212 3276 3164 3332
rect 3220 3276 3230 3332
rect 5506 3276 5516 3332
rect 5572 3276 5852 3332
rect 5908 3276 5918 3332
rect 9266 3108 9276 3164
rect 9332 3108 9380 3164
rect 9436 3108 9484 3164
rect 9540 3108 9550 3164
rect 17330 3108 17340 3164
rect 17396 3108 17444 3164
rect 17500 3108 17548 3164
rect 17604 3108 17614 3164
rect 25394 3108 25404 3164
rect 25460 3108 25508 3164
rect 25564 3108 25612 3164
rect 25668 3108 25678 3164
rect 33458 3108 33468 3164
rect 33524 3108 33572 3164
rect 33628 3108 33676 3164
rect 33732 3108 33742 3164
rect 34200 1204 35000 1232
rect 25106 1148 25116 1204
rect 25172 1148 35000 1204
rect 34200 1120 35000 1148
<< via3 >>
rect 27468 33068 27524 33124
rect 28924 31948 28980 32004
rect 26236 31724 26292 31780
rect 10444 31612 10500 31668
rect 9276 31332 9332 31388
rect 9380 31332 9436 31388
rect 9484 31332 9540 31388
rect 17340 31332 17396 31388
rect 17444 31332 17500 31388
rect 17548 31332 17604 31388
rect 25404 31332 25460 31388
rect 25508 31332 25564 31388
rect 25612 31332 25668 31388
rect 33468 31332 33524 31388
rect 33572 31332 33628 31388
rect 33676 31332 33732 31388
rect 5244 30548 5300 30604
rect 5348 30548 5404 30604
rect 5452 30548 5508 30604
rect 13308 30548 13364 30604
rect 13412 30548 13468 30604
rect 13516 30548 13572 30604
rect 21372 30548 21428 30604
rect 21476 30548 21532 30604
rect 21580 30548 21636 30604
rect 29436 30548 29492 30604
rect 29540 30548 29596 30604
rect 29644 30548 29700 30604
rect 28700 30492 28756 30548
rect 14924 30156 14980 30212
rect 9276 29764 9332 29820
rect 9380 29764 9436 29820
rect 9484 29764 9540 29820
rect 17340 29764 17396 29820
rect 17444 29764 17500 29820
rect 17548 29764 17604 29820
rect 25404 29764 25460 29820
rect 25508 29764 25564 29820
rect 25612 29764 25668 29820
rect 33468 29764 33524 29820
rect 33572 29764 33628 29820
rect 33676 29764 33732 29820
rect 15036 29484 15092 29540
rect 26236 29372 26292 29428
rect 29820 29036 29876 29092
rect 5244 28980 5300 29036
rect 5348 28980 5404 29036
rect 5452 28980 5508 29036
rect 13308 28980 13364 29036
rect 13412 28980 13468 29036
rect 13516 28980 13572 29036
rect 21372 28980 21428 29036
rect 21476 28980 21532 29036
rect 21580 28980 21636 29036
rect 29436 28980 29492 29036
rect 29540 28980 29596 29036
rect 29644 28980 29700 29036
rect 20972 28812 21028 28868
rect 15036 28476 15092 28532
rect 29036 28476 29092 28532
rect 10332 28364 10388 28420
rect 9276 28196 9332 28252
rect 9380 28196 9436 28252
rect 9484 28196 9540 28252
rect 17340 28196 17396 28252
rect 17444 28196 17500 28252
rect 17548 28196 17604 28252
rect 25404 28196 25460 28252
rect 25508 28196 25564 28252
rect 25612 28196 25668 28252
rect 33468 28196 33524 28252
rect 33572 28196 33628 28252
rect 33676 28196 33732 28252
rect 22540 28140 22596 28196
rect 30268 28028 30324 28084
rect 13132 27804 13188 27860
rect 8988 27692 9044 27748
rect 22540 27692 22596 27748
rect 5244 27412 5300 27468
rect 5348 27412 5404 27468
rect 5452 27412 5508 27468
rect 13308 27412 13364 27468
rect 13412 27412 13468 27468
rect 13516 27412 13572 27468
rect 21372 27412 21428 27468
rect 21476 27412 21532 27468
rect 21580 27412 21636 27468
rect 29436 27412 29492 27468
rect 29540 27412 29596 27468
rect 29644 27412 29700 27468
rect 14140 27356 14196 27412
rect 14812 27356 14868 27412
rect 7196 26908 7252 26964
rect 11228 26908 11284 26964
rect 12572 26908 12628 26964
rect 10332 26684 10388 26740
rect 9276 26628 9332 26684
rect 9380 26628 9436 26684
rect 9484 26628 9540 26684
rect 17340 26628 17396 26684
rect 17444 26628 17500 26684
rect 17548 26628 17604 26684
rect 25404 26628 25460 26684
rect 25508 26628 25564 26684
rect 25612 26628 25668 26684
rect 33468 26628 33524 26684
rect 33572 26628 33628 26684
rect 33676 26628 33732 26684
rect 14812 26572 14868 26628
rect 18508 26572 18564 26628
rect 20972 26572 21028 26628
rect 29820 26572 29876 26628
rect 6412 26460 6468 26516
rect 15260 26460 15316 26516
rect 8988 26236 9044 26292
rect 29036 26236 29092 26292
rect 16156 26124 16212 26180
rect 6300 25900 6356 25956
rect 5244 25844 5300 25900
rect 5348 25844 5404 25900
rect 5452 25844 5508 25900
rect 13308 25844 13364 25900
rect 13412 25844 13468 25900
rect 13516 25844 13572 25900
rect 21372 25844 21428 25900
rect 21476 25844 21532 25900
rect 21580 25844 21636 25900
rect 6076 25788 6132 25844
rect 12684 25788 12740 25844
rect 29436 25844 29492 25900
rect 29540 25844 29596 25900
rect 29644 25844 29700 25900
rect 10444 25564 10500 25620
rect 28924 25340 28980 25396
rect 6076 25228 6132 25284
rect 6300 25228 6356 25284
rect 28140 25228 28196 25284
rect 28364 25228 28420 25284
rect 28588 25228 28644 25284
rect 6412 25116 6468 25172
rect 9276 25060 9332 25116
rect 9380 25060 9436 25116
rect 9484 25060 9540 25116
rect 12684 25116 12740 25172
rect 17340 25060 17396 25116
rect 17444 25060 17500 25116
rect 17548 25060 17604 25116
rect 14924 25004 14980 25060
rect 12572 24892 12628 24948
rect 13132 24892 13188 24948
rect 25404 25060 25460 25116
rect 25508 25060 25564 25116
rect 25612 25060 25668 25116
rect 33468 25060 33524 25116
rect 33572 25060 33628 25116
rect 33676 25060 33732 25116
rect 27468 25004 27524 25060
rect 19852 24892 19908 24948
rect 15260 24780 15316 24836
rect 28140 24668 28196 24724
rect 19852 24444 19908 24500
rect 5244 24276 5300 24332
rect 5348 24276 5404 24332
rect 5452 24276 5508 24332
rect 13308 24276 13364 24332
rect 13412 24276 13468 24332
rect 13516 24276 13572 24332
rect 26236 24332 26292 24388
rect 21372 24276 21428 24332
rect 21476 24276 21532 24332
rect 21580 24276 21636 24332
rect 29436 24276 29492 24332
rect 29540 24276 29596 24332
rect 29644 24276 29700 24332
rect 21868 24108 21924 24164
rect 14140 23996 14196 24052
rect 11228 23772 11284 23828
rect 9276 23492 9332 23548
rect 9380 23492 9436 23548
rect 9484 23492 9540 23548
rect 17340 23492 17396 23548
rect 17444 23492 17500 23548
rect 17548 23492 17604 23548
rect 25404 23492 25460 23548
rect 25508 23492 25564 23548
rect 25612 23492 25668 23548
rect 33468 23492 33524 23548
rect 33572 23492 33628 23548
rect 33676 23492 33732 23548
rect 16156 23212 16212 23268
rect 16380 23212 16436 23268
rect 21756 23212 21812 23268
rect 28700 23100 28756 23156
rect 26796 22988 26852 23044
rect 18508 22764 18564 22820
rect 5244 22708 5300 22764
rect 5348 22708 5404 22764
rect 5452 22708 5508 22764
rect 13308 22708 13364 22764
rect 13412 22708 13468 22764
rect 13516 22708 13572 22764
rect 21372 22708 21428 22764
rect 21476 22708 21532 22764
rect 21580 22708 21636 22764
rect 29436 22708 29492 22764
rect 29540 22708 29596 22764
rect 29644 22708 29700 22764
rect 21756 22652 21812 22708
rect 16380 22316 16436 22372
rect 27020 22092 27076 22148
rect 16044 21980 16100 22036
rect 9276 21924 9332 21980
rect 9380 21924 9436 21980
rect 9484 21924 9540 21980
rect 17340 21924 17396 21980
rect 17444 21924 17500 21980
rect 17548 21924 17604 21980
rect 25404 21924 25460 21980
rect 25508 21924 25564 21980
rect 25612 21924 25668 21980
rect 33468 21924 33524 21980
rect 33572 21924 33628 21980
rect 33676 21924 33732 21980
rect 12572 21644 12628 21700
rect 21756 21644 21812 21700
rect 27244 21420 27300 21476
rect 5244 21140 5300 21196
rect 5348 21140 5404 21196
rect 5452 21140 5508 21196
rect 13308 21140 13364 21196
rect 13412 21140 13468 21196
rect 13516 21140 13572 21196
rect 21372 21140 21428 21196
rect 21476 21140 21532 21196
rect 21580 21140 21636 21196
rect 29436 21140 29492 21196
rect 29540 21140 29596 21196
rect 29644 21140 29700 21196
rect 25788 21084 25844 21140
rect 26908 21084 26964 21140
rect 28588 21084 28644 21140
rect 21756 20636 21812 20692
rect 15036 20412 15092 20468
rect 29148 20412 29204 20468
rect 9276 20356 9332 20412
rect 9380 20356 9436 20412
rect 9484 20356 9540 20412
rect 17340 20356 17396 20412
rect 17444 20356 17500 20412
rect 17548 20356 17604 20412
rect 25404 20356 25460 20412
rect 25508 20356 25564 20412
rect 25612 20356 25668 20412
rect 33468 20356 33524 20412
rect 33572 20356 33628 20412
rect 33676 20356 33732 20412
rect 26572 20300 26628 20356
rect 27244 20300 27300 20356
rect 25228 20188 25284 20244
rect 25788 20188 25844 20244
rect 26908 20076 26964 20132
rect 30268 20076 30324 20132
rect 21868 19852 21924 19908
rect 27244 19964 27300 20020
rect 29148 19964 29204 20020
rect 27020 19852 27076 19908
rect 29036 19852 29092 19908
rect 5852 19740 5908 19796
rect 5244 19572 5300 19628
rect 5348 19572 5404 19628
rect 5452 19572 5508 19628
rect 13308 19572 13364 19628
rect 13412 19572 13468 19628
rect 13516 19572 13572 19628
rect 21372 19572 21428 19628
rect 21476 19572 21532 19628
rect 21580 19572 21636 19628
rect 15036 19516 15092 19572
rect 20860 19292 20916 19348
rect 29436 19572 29492 19628
rect 29540 19572 29596 19628
rect 29644 19572 29700 19628
rect 28252 19180 28308 19236
rect 28476 19180 28532 19236
rect 12124 18844 12180 18900
rect 16044 18844 16100 18900
rect 26572 18844 26628 18900
rect 27244 18844 27300 18900
rect 28476 18844 28532 18900
rect 9276 18788 9332 18844
rect 9380 18788 9436 18844
rect 9484 18788 9540 18844
rect 17340 18788 17396 18844
rect 17444 18788 17500 18844
rect 17548 18788 17604 18844
rect 25404 18788 25460 18844
rect 25508 18788 25564 18844
rect 25612 18788 25668 18844
rect 33468 18788 33524 18844
rect 33572 18788 33628 18844
rect 33676 18788 33732 18844
rect 27804 18732 27860 18788
rect 28364 18732 28420 18788
rect 20188 18508 20244 18564
rect 16044 18396 16100 18452
rect 27804 18396 27860 18452
rect 29148 18396 29204 18452
rect 30940 18396 30996 18452
rect 5244 18004 5300 18060
rect 5348 18004 5404 18060
rect 5452 18004 5508 18060
rect 13308 18004 13364 18060
rect 13412 18004 13468 18060
rect 13516 18004 13572 18060
rect 21372 18004 21428 18060
rect 21476 18004 21532 18060
rect 21580 18004 21636 18060
rect 29436 18004 29492 18060
rect 29540 18004 29596 18060
rect 29644 18004 29700 18060
rect 7196 17836 7252 17892
rect 5852 17612 5908 17668
rect 26796 17612 26852 17668
rect 28476 17388 28532 17444
rect 27020 17276 27076 17332
rect 9276 17220 9332 17276
rect 9380 17220 9436 17276
rect 9484 17220 9540 17276
rect 17340 17220 17396 17276
rect 17444 17220 17500 17276
rect 17548 17220 17604 17276
rect 25404 17220 25460 17276
rect 25508 17220 25564 17276
rect 25612 17220 25668 17276
rect 33468 17220 33524 17276
rect 33572 17220 33628 17276
rect 33676 17220 33732 17276
rect 28700 16940 28756 16996
rect 5244 16436 5300 16492
rect 5348 16436 5404 16492
rect 5452 16436 5508 16492
rect 13308 16436 13364 16492
rect 13412 16436 13468 16492
rect 13516 16436 13572 16492
rect 21372 16436 21428 16492
rect 21476 16436 21532 16492
rect 21580 16436 21636 16492
rect 29436 16436 29492 16492
rect 29540 16436 29596 16492
rect 29644 16436 29700 16492
rect 19292 16044 19348 16100
rect 27020 16044 27076 16100
rect 29148 16044 29204 16100
rect 9276 15652 9332 15708
rect 9380 15652 9436 15708
rect 9484 15652 9540 15708
rect 17340 15652 17396 15708
rect 17444 15652 17500 15708
rect 17548 15652 17604 15708
rect 25404 15652 25460 15708
rect 25508 15652 25564 15708
rect 25612 15652 25668 15708
rect 27020 15708 27076 15764
rect 30156 15708 30212 15764
rect 33468 15652 33524 15708
rect 33572 15652 33628 15708
rect 33676 15652 33732 15708
rect 12572 15484 12628 15540
rect 25900 15372 25956 15428
rect 28700 15372 28756 15428
rect 19628 15260 19684 15316
rect 30940 15036 30996 15092
rect 28588 14924 28644 14980
rect 5244 14868 5300 14924
rect 5348 14868 5404 14924
rect 5452 14868 5508 14924
rect 13308 14868 13364 14924
rect 13412 14868 13468 14924
rect 13516 14868 13572 14924
rect 21372 14868 21428 14924
rect 21476 14868 21532 14924
rect 21580 14868 21636 14924
rect 29436 14868 29492 14924
rect 29540 14868 29596 14924
rect 29644 14868 29700 14924
rect 19628 14812 19684 14868
rect 19628 14588 19684 14644
rect 19292 14364 19348 14420
rect 19068 14140 19124 14196
rect 25900 14140 25956 14196
rect 28588 14140 28644 14196
rect 9276 14084 9332 14140
rect 9380 14084 9436 14140
rect 9484 14084 9540 14140
rect 17340 14084 17396 14140
rect 17444 14084 17500 14140
rect 17548 14084 17604 14140
rect 25404 14084 25460 14140
rect 25508 14084 25564 14140
rect 25612 14084 25668 14140
rect 33468 14084 33524 14140
rect 33572 14084 33628 14140
rect 33676 14084 33732 14140
rect 26908 14028 26964 14084
rect 28252 13916 28308 13972
rect 20860 13356 20916 13412
rect 5244 13300 5300 13356
rect 5348 13300 5404 13356
rect 5452 13300 5508 13356
rect 13308 13300 13364 13356
rect 13412 13300 13468 13356
rect 13516 13300 13572 13356
rect 21372 13300 21428 13356
rect 21476 13300 21532 13356
rect 21580 13300 21636 13356
rect 29436 13300 29492 13356
rect 29540 13300 29596 13356
rect 29644 13300 29700 13356
rect 19628 13132 19684 13188
rect 20076 13132 20132 13188
rect 19068 12908 19124 12964
rect 29148 12684 29204 12740
rect 9276 12516 9332 12572
rect 9380 12516 9436 12572
rect 9484 12516 9540 12572
rect 17340 12516 17396 12572
rect 17444 12516 17500 12572
rect 17548 12516 17604 12572
rect 25404 12516 25460 12572
rect 25508 12516 25564 12572
rect 25612 12516 25668 12572
rect 33468 12516 33524 12572
rect 33572 12516 33628 12572
rect 33676 12516 33732 12572
rect 12124 12460 12180 12516
rect 25228 12124 25284 12180
rect 29036 11788 29092 11844
rect 5244 11732 5300 11788
rect 5348 11732 5404 11788
rect 5452 11732 5508 11788
rect 13308 11732 13364 11788
rect 13412 11732 13468 11788
rect 13516 11732 13572 11788
rect 21372 11732 21428 11788
rect 21476 11732 21532 11788
rect 21580 11732 21636 11788
rect 29436 11732 29492 11788
rect 29540 11732 29596 11788
rect 29644 11732 29700 11788
rect 30156 11452 30212 11508
rect 9276 10948 9332 11004
rect 9380 10948 9436 11004
rect 9484 10948 9540 11004
rect 17340 10948 17396 11004
rect 17444 10948 17500 11004
rect 17548 10948 17604 11004
rect 25404 10948 25460 11004
rect 25508 10948 25564 11004
rect 25612 10948 25668 11004
rect 33468 10948 33524 11004
rect 33572 10948 33628 11004
rect 33676 10948 33732 11004
rect 5068 10332 5124 10388
rect 5244 10164 5300 10220
rect 5348 10164 5404 10220
rect 5452 10164 5508 10220
rect 13308 10164 13364 10220
rect 13412 10164 13468 10220
rect 13516 10164 13572 10220
rect 21372 10164 21428 10220
rect 21476 10164 21532 10220
rect 21580 10164 21636 10220
rect 29436 10164 29492 10220
rect 29540 10164 29596 10220
rect 29644 10164 29700 10220
rect 5740 9772 5796 9828
rect 9276 9380 9332 9436
rect 9380 9380 9436 9436
rect 9484 9380 9540 9436
rect 17340 9380 17396 9436
rect 17444 9380 17500 9436
rect 17548 9380 17604 9436
rect 25404 9380 25460 9436
rect 25508 9380 25564 9436
rect 25612 9380 25668 9436
rect 33468 9380 33524 9436
rect 33572 9380 33628 9436
rect 33676 9380 33732 9436
rect 30268 9212 30324 9268
rect 5244 8596 5300 8652
rect 5348 8596 5404 8652
rect 5452 8596 5508 8652
rect 13308 8596 13364 8652
rect 13412 8596 13468 8652
rect 13516 8596 13572 8652
rect 21372 8596 21428 8652
rect 21476 8596 21532 8652
rect 21580 8596 21636 8652
rect 29436 8596 29492 8652
rect 29540 8596 29596 8652
rect 29644 8596 29700 8652
rect 5852 7756 5908 7812
rect 9276 7812 9332 7868
rect 9380 7812 9436 7868
rect 9484 7812 9540 7868
rect 17340 7812 17396 7868
rect 17444 7812 17500 7868
rect 17548 7812 17604 7868
rect 25404 7812 25460 7868
rect 25508 7812 25564 7868
rect 25612 7812 25668 7868
rect 33468 7812 33524 7868
rect 33572 7812 33628 7868
rect 33676 7812 33732 7868
rect 21756 7756 21812 7812
rect 23324 7756 23380 7812
rect 23548 7532 23604 7588
rect 26684 7532 26740 7588
rect 27020 7532 27076 7588
rect 27692 7084 27748 7140
rect 5244 7028 5300 7084
rect 5348 7028 5404 7084
rect 5452 7028 5508 7084
rect 13308 7028 13364 7084
rect 13412 7028 13468 7084
rect 13516 7028 13572 7084
rect 21372 7028 21428 7084
rect 21476 7028 21532 7084
rect 21580 7028 21636 7084
rect 29436 7028 29492 7084
rect 29540 7028 29596 7084
rect 29644 7028 29700 7084
rect 24220 6860 24276 6916
rect 27020 6860 27076 6916
rect 5740 6524 5796 6580
rect 24444 6300 24500 6356
rect 9276 6244 9332 6300
rect 9380 6244 9436 6300
rect 9484 6244 9540 6300
rect 17340 6244 17396 6300
rect 17444 6244 17500 6300
rect 17548 6244 17604 6300
rect 25404 6244 25460 6300
rect 25508 6244 25564 6300
rect 25612 6244 25668 6300
rect 33468 6244 33524 6300
rect 33572 6244 33628 6300
rect 33676 6244 33732 6300
rect 5068 5964 5124 6020
rect 23548 5852 23604 5908
rect 24780 5852 24836 5908
rect 21756 5628 21812 5684
rect 23324 5516 23380 5572
rect 5244 5460 5300 5516
rect 5348 5460 5404 5516
rect 5452 5460 5508 5516
rect 13308 5460 13364 5516
rect 13412 5460 13468 5516
rect 13516 5460 13572 5516
rect 21372 5460 21428 5516
rect 21476 5460 21532 5516
rect 21580 5460 21636 5516
rect 29436 5460 29492 5516
rect 29540 5460 29596 5516
rect 29644 5460 29700 5516
rect 24220 5404 24276 5460
rect 24780 5068 24836 5124
rect 26684 5068 26740 5124
rect 9276 4676 9332 4732
rect 9380 4676 9436 4732
rect 9484 4676 9540 4732
rect 17340 4676 17396 4732
rect 17444 4676 17500 4732
rect 17548 4676 17604 4732
rect 25404 4676 25460 4732
rect 25508 4676 25564 4732
rect 25612 4676 25668 4732
rect 33468 4676 33524 4732
rect 33572 4676 33628 4732
rect 33676 4676 33732 4732
rect 24444 4508 24500 4564
rect 5244 3892 5300 3948
rect 5348 3892 5404 3948
rect 5452 3892 5508 3948
rect 13308 3892 13364 3948
rect 13412 3892 13468 3948
rect 13516 3892 13572 3948
rect 21372 3892 21428 3948
rect 21476 3892 21532 3948
rect 21580 3892 21636 3948
rect 29436 3892 29492 3948
rect 29540 3892 29596 3948
rect 29644 3892 29700 3948
rect 27692 3500 27748 3556
rect 5852 3276 5908 3332
rect 9276 3108 9332 3164
rect 9380 3108 9436 3164
rect 9484 3108 9540 3164
rect 17340 3108 17396 3164
rect 17444 3108 17500 3164
rect 17548 3108 17604 3164
rect 25404 3108 25460 3164
rect 25508 3108 25564 3164
rect 25612 3108 25668 3164
rect 33468 3108 33524 3164
rect 33572 3108 33628 3164
rect 33676 3108 33732 3164
<< metal4 >>
rect 27468 33124 27524 33134
rect 26236 31780 26292 31790
rect 10444 31668 10500 31678
rect 5216 30604 5536 31420
rect 5216 30548 5244 30604
rect 5300 30548 5348 30604
rect 5404 30548 5452 30604
rect 5508 30548 5536 30604
rect 5216 29036 5536 30548
rect 5216 28980 5244 29036
rect 5300 28980 5348 29036
rect 5404 28980 5452 29036
rect 5508 28980 5536 29036
rect 5216 27468 5536 28980
rect 9248 31388 9568 31420
rect 9248 31332 9276 31388
rect 9332 31332 9380 31388
rect 9436 31332 9484 31388
rect 9540 31332 9568 31388
rect 9248 29820 9568 31332
rect 9248 29764 9276 29820
rect 9332 29764 9380 29820
rect 9436 29764 9484 29820
rect 9540 29764 9568 29820
rect 9248 28252 9568 29764
rect 9248 28196 9276 28252
rect 9332 28196 9380 28252
rect 9436 28196 9484 28252
rect 9540 28196 9568 28252
rect 5216 27412 5244 27468
rect 5300 27412 5348 27468
rect 5404 27412 5452 27468
rect 5508 27412 5536 27468
rect 5216 25900 5536 27412
rect 8988 27748 9044 27758
rect 7196 26964 7252 26974
rect 6412 26516 6468 26526
rect 5216 25844 5244 25900
rect 5300 25844 5348 25900
rect 5404 25844 5452 25900
rect 5508 25844 5536 25900
rect 6300 25956 6356 25966
rect 5216 24332 5536 25844
rect 6076 25844 6132 25854
rect 6076 25284 6132 25788
rect 6076 25218 6132 25228
rect 6300 25284 6356 25900
rect 6300 25218 6356 25228
rect 6412 25172 6468 26460
rect 6412 25106 6468 25116
rect 5216 24276 5244 24332
rect 5300 24276 5348 24332
rect 5404 24276 5452 24332
rect 5508 24276 5536 24332
rect 5216 22764 5536 24276
rect 5216 22708 5244 22764
rect 5300 22708 5348 22764
rect 5404 22708 5452 22764
rect 5508 22708 5536 22764
rect 5216 21196 5536 22708
rect 5216 21140 5244 21196
rect 5300 21140 5348 21196
rect 5404 21140 5452 21196
rect 5508 21140 5536 21196
rect 5216 19628 5536 21140
rect 5216 19572 5244 19628
rect 5300 19572 5348 19628
rect 5404 19572 5452 19628
rect 5508 19572 5536 19628
rect 5216 18060 5536 19572
rect 5216 18004 5244 18060
rect 5300 18004 5348 18060
rect 5404 18004 5452 18060
rect 5508 18004 5536 18060
rect 5216 16492 5536 18004
rect 5852 19796 5908 19806
rect 5852 17668 5908 19740
rect 7196 17892 7252 26908
rect 8988 26292 9044 27692
rect 8988 26226 9044 26236
rect 9248 26684 9568 28196
rect 9248 26628 9276 26684
rect 9332 26628 9380 26684
rect 9436 26628 9484 26684
rect 9540 26628 9568 26684
rect 10332 28420 10388 28430
rect 10332 26740 10388 28364
rect 10332 26674 10388 26684
rect 7196 17826 7252 17836
rect 9248 25116 9568 26628
rect 10444 25620 10500 31612
rect 13280 30604 13600 31420
rect 13280 30548 13308 30604
rect 13364 30548 13412 30604
rect 13468 30548 13516 30604
rect 13572 30548 13600 30604
rect 13280 29036 13600 30548
rect 17312 31388 17632 31420
rect 17312 31332 17340 31388
rect 17396 31332 17444 31388
rect 17500 31332 17548 31388
rect 17604 31332 17632 31388
rect 13280 28980 13308 29036
rect 13364 28980 13412 29036
rect 13468 28980 13516 29036
rect 13572 28980 13600 29036
rect 13132 27860 13188 27870
rect 10444 25554 10500 25564
rect 11228 26964 11284 26974
rect 9248 25060 9276 25116
rect 9332 25060 9380 25116
rect 9436 25060 9484 25116
rect 9540 25060 9568 25116
rect 9248 23548 9568 25060
rect 11228 23828 11284 26908
rect 12572 26964 12628 26974
rect 12572 24948 12628 26908
rect 12684 25844 12740 25854
rect 12684 25172 12740 25788
rect 12684 25106 12740 25116
rect 12572 24882 12628 24892
rect 13132 24948 13188 27804
rect 13132 24882 13188 24892
rect 13280 27468 13600 28980
rect 13280 27412 13308 27468
rect 13364 27412 13412 27468
rect 13468 27412 13516 27468
rect 13572 27412 13600 27468
rect 14924 30212 14980 30222
rect 13280 25900 13600 27412
rect 13280 25844 13308 25900
rect 13364 25844 13412 25900
rect 13468 25844 13516 25900
rect 13572 25844 13600 25900
rect 11228 23762 11284 23772
rect 13280 24332 13600 25844
rect 13280 24276 13308 24332
rect 13364 24276 13412 24332
rect 13468 24276 13516 24332
rect 13572 24276 13600 24332
rect 9248 23492 9276 23548
rect 9332 23492 9380 23548
rect 9436 23492 9484 23548
rect 9540 23492 9568 23548
rect 9248 21980 9568 23492
rect 9248 21924 9276 21980
rect 9332 21924 9380 21980
rect 9436 21924 9484 21980
rect 9540 21924 9568 21980
rect 9248 20412 9568 21924
rect 13280 22764 13600 24276
rect 14140 27412 14196 27422
rect 14140 24052 14196 27356
rect 14812 27412 14868 27422
rect 14812 26628 14868 27356
rect 14812 26562 14868 26572
rect 14924 25060 14980 30156
rect 17312 29820 17632 31332
rect 17312 29764 17340 29820
rect 17396 29764 17444 29820
rect 17500 29764 17548 29820
rect 17604 29764 17632 29820
rect 15036 29540 15092 29550
rect 15036 28532 15092 29484
rect 15036 28466 15092 28476
rect 17312 28252 17632 29764
rect 21344 30604 21664 31420
rect 21344 30548 21372 30604
rect 21428 30548 21476 30604
rect 21532 30548 21580 30604
rect 21636 30548 21664 30604
rect 21344 29036 21664 30548
rect 21344 28980 21372 29036
rect 21428 28980 21476 29036
rect 21532 28980 21580 29036
rect 21636 28980 21664 29036
rect 17312 28196 17340 28252
rect 17396 28196 17444 28252
rect 17500 28196 17548 28252
rect 17604 28196 17632 28252
rect 17312 26684 17632 28196
rect 17312 26628 17340 26684
rect 17396 26628 17444 26684
rect 17500 26628 17548 26684
rect 17604 26628 17632 26684
rect 20972 28868 21028 28878
rect 14924 24994 14980 25004
rect 15260 26516 15316 26526
rect 15260 24836 15316 26460
rect 15260 24770 15316 24780
rect 16156 26180 16212 26190
rect 14140 23986 14196 23996
rect 16156 23268 16212 26124
rect 17312 25116 17632 26628
rect 17312 25060 17340 25116
rect 17396 25060 17444 25116
rect 17500 25060 17548 25116
rect 17604 25060 17632 25116
rect 17312 23548 17632 25060
rect 17312 23492 17340 23548
rect 17396 23492 17444 23548
rect 17500 23492 17548 23548
rect 17604 23492 17632 23548
rect 16156 23202 16212 23212
rect 16380 23268 16436 23278
rect 13280 22708 13308 22764
rect 13364 22708 13412 22764
rect 13468 22708 13516 22764
rect 13572 22708 13600 22764
rect 9248 20356 9276 20412
rect 9332 20356 9380 20412
rect 9436 20356 9484 20412
rect 9540 20356 9568 20412
rect 9248 18844 9568 20356
rect 12572 21700 12628 21710
rect 9248 18788 9276 18844
rect 9332 18788 9380 18844
rect 9436 18788 9484 18844
rect 9540 18788 9568 18844
rect 5852 17602 5908 17612
rect 5216 16436 5244 16492
rect 5300 16436 5348 16492
rect 5404 16436 5452 16492
rect 5508 16436 5536 16492
rect 5216 14924 5536 16436
rect 5216 14868 5244 14924
rect 5300 14868 5348 14924
rect 5404 14868 5452 14924
rect 5508 14868 5536 14924
rect 5216 13356 5536 14868
rect 5216 13300 5244 13356
rect 5300 13300 5348 13356
rect 5404 13300 5452 13356
rect 5508 13300 5536 13356
rect 5216 11788 5536 13300
rect 5216 11732 5244 11788
rect 5300 11732 5348 11788
rect 5404 11732 5452 11788
rect 5508 11732 5536 11788
rect 5068 10388 5124 10398
rect 5068 6020 5124 10332
rect 5068 5954 5124 5964
rect 5216 10220 5536 11732
rect 5216 10164 5244 10220
rect 5300 10164 5348 10220
rect 5404 10164 5452 10220
rect 5508 10164 5536 10220
rect 5216 8652 5536 10164
rect 9248 17276 9568 18788
rect 9248 17220 9276 17276
rect 9332 17220 9380 17276
rect 9436 17220 9484 17276
rect 9540 17220 9568 17276
rect 9248 15708 9568 17220
rect 9248 15652 9276 15708
rect 9332 15652 9380 15708
rect 9436 15652 9484 15708
rect 9540 15652 9568 15708
rect 9248 14140 9568 15652
rect 9248 14084 9276 14140
rect 9332 14084 9380 14140
rect 9436 14084 9484 14140
rect 9540 14084 9568 14140
rect 9248 12572 9568 14084
rect 9248 12516 9276 12572
rect 9332 12516 9380 12572
rect 9436 12516 9484 12572
rect 9540 12516 9568 12572
rect 9248 11004 9568 12516
rect 12124 18900 12180 18910
rect 12124 12516 12180 18844
rect 12572 15540 12628 21644
rect 12572 15474 12628 15484
rect 13280 21196 13600 22708
rect 16380 22372 16436 23212
rect 16380 22306 16436 22316
rect 13280 21140 13308 21196
rect 13364 21140 13412 21196
rect 13468 21140 13516 21196
rect 13572 21140 13600 21196
rect 13280 19628 13600 21140
rect 16044 22036 16100 22046
rect 13280 19572 13308 19628
rect 13364 19572 13412 19628
rect 13468 19572 13516 19628
rect 13572 19572 13600 19628
rect 13280 18060 13600 19572
rect 15036 20468 15092 20478
rect 15036 19572 15092 20412
rect 15036 19506 15092 19516
rect 16044 18900 16100 21980
rect 16044 18452 16100 18844
rect 16044 18386 16100 18396
rect 17312 21980 17632 23492
rect 18508 26628 18564 26638
rect 18508 22820 18564 26572
rect 20972 26628 21028 28812
rect 20972 26562 21028 26572
rect 21344 27468 21664 28980
rect 25376 31388 25696 31420
rect 25376 31332 25404 31388
rect 25460 31332 25508 31388
rect 25564 31332 25612 31388
rect 25668 31332 25696 31388
rect 25376 29820 25696 31332
rect 25376 29764 25404 29820
rect 25460 29764 25508 29820
rect 25564 29764 25612 29820
rect 25668 29764 25696 29820
rect 25376 28252 25696 29764
rect 22540 28196 22596 28206
rect 22540 27748 22596 28140
rect 22540 27682 22596 27692
rect 25376 28196 25404 28252
rect 25460 28196 25508 28252
rect 25564 28196 25612 28252
rect 25668 28196 25696 28252
rect 21344 27412 21372 27468
rect 21428 27412 21476 27468
rect 21532 27412 21580 27468
rect 21636 27412 21664 27468
rect 21344 25900 21664 27412
rect 21344 25844 21372 25900
rect 21428 25844 21476 25900
rect 21532 25844 21580 25900
rect 21636 25844 21664 25900
rect 19852 24948 19908 24958
rect 19852 24500 19908 24892
rect 19852 24434 19908 24444
rect 18508 22754 18564 22764
rect 21344 24332 21664 25844
rect 21344 24276 21372 24332
rect 21428 24276 21476 24332
rect 21532 24276 21580 24332
rect 21636 24276 21664 24332
rect 21344 22764 21664 24276
rect 25376 26684 25696 28196
rect 25376 26628 25404 26684
rect 25460 26628 25508 26684
rect 25564 26628 25612 26684
rect 25668 26628 25696 26684
rect 25376 25116 25696 26628
rect 25376 25060 25404 25116
rect 25460 25060 25508 25116
rect 25564 25060 25612 25116
rect 25668 25060 25696 25116
rect 21868 24164 21924 24174
rect 17312 21924 17340 21980
rect 17396 21924 17444 21980
rect 17500 21924 17548 21980
rect 17604 21924 17632 21980
rect 17312 20412 17632 21924
rect 17312 20356 17340 20412
rect 17396 20356 17444 20412
rect 17500 20356 17548 20412
rect 17604 20356 17632 20412
rect 17312 18844 17632 20356
rect 21344 22708 21372 22764
rect 21428 22708 21476 22764
rect 21532 22708 21580 22764
rect 21636 22708 21664 22764
rect 21344 21196 21664 22708
rect 21756 23268 21812 23278
rect 21756 22708 21812 23212
rect 21756 22642 21812 22652
rect 21344 21140 21372 21196
rect 21428 21140 21476 21196
rect 21532 21140 21580 21196
rect 21636 21140 21664 21196
rect 21344 19628 21664 21140
rect 21756 21700 21812 21710
rect 21756 20692 21812 21644
rect 21756 20626 21812 20636
rect 21868 19908 21924 24108
rect 25376 23548 25696 25060
rect 26236 29428 26292 31724
rect 26236 24388 26292 29372
rect 27468 25060 27524 33068
rect 28924 32004 28980 32014
rect 28700 30548 28756 30558
rect 27468 24994 27524 25004
rect 28140 25284 28196 25294
rect 28140 24724 28196 25228
rect 28140 24658 28196 24668
rect 28364 25284 28420 25294
rect 26236 24322 26292 24332
rect 25376 23492 25404 23548
rect 25460 23492 25508 23548
rect 25564 23492 25612 23548
rect 25668 23492 25696 23548
rect 25376 21980 25696 23492
rect 25376 21924 25404 21980
rect 25460 21924 25508 21980
rect 25564 21924 25612 21980
rect 25668 21924 25696 21980
rect 25376 20412 25696 21924
rect 26796 23044 26852 23054
rect 25376 20356 25404 20412
rect 25460 20356 25508 20412
rect 25564 20356 25612 20412
rect 25668 20356 25696 20412
rect 21868 19842 21924 19852
rect 25228 20244 25284 20254
rect 21344 19572 21372 19628
rect 21428 19572 21476 19628
rect 21532 19572 21580 19628
rect 21636 19572 21664 19628
rect 17312 18788 17340 18844
rect 17396 18788 17444 18844
rect 17500 18788 17548 18844
rect 17604 18788 17632 18844
rect 13280 18004 13308 18060
rect 13364 18004 13412 18060
rect 13468 18004 13516 18060
rect 13572 18004 13600 18060
rect 13280 16492 13600 18004
rect 13280 16436 13308 16492
rect 13364 16436 13412 16492
rect 13468 16436 13516 16492
rect 13572 16436 13600 16492
rect 12124 12450 12180 12460
rect 13280 14924 13600 16436
rect 13280 14868 13308 14924
rect 13364 14868 13412 14924
rect 13468 14868 13516 14924
rect 13572 14868 13600 14924
rect 13280 13356 13600 14868
rect 13280 13300 13308 13356
rect 13364 13300 13412 13356
rect 13468 13300 13516 13356
rect 13572 13300 13600 13356
rect 9248 10948 9276 11004
rect 9332 10948 9380 11004
rect 9436 10948 9484 11004
rect 9540 10948 9568 11004
rect 5216 8596 5244 8652
rect 5300 8596 5348 8652
rect 5404 8596 5452 8652
rect 5508 8596 5536 8652
rect 5216 7084 5536 8596
rect 5216 7028 5244 7084
rect 5300 7028 5348 7084
rect 5404 7028 5452 7084
rect 5508 7028 5536 7084
rect 5216 5516 5536 7028
rect 5740 9828 5796 9838
rect 5740 6580 5796 9772
rect 9248 9436 9568 10948
rect 9248 9380 9276 9436
rect 9332 9380 9380 9436
rect 9436 9380 9484 9436
rect 9540 9380 9568 9436
rect 9248 7868 9568 9380
rect 5740 6514 5796 6524
rect 5852 7812 5908 7822
rect 5216 5460 5244 5516
rect 5300 5460 5348 5516
rect 5404 5460 5452 5516
rect 5508 5460 5536 5516
rect 5216 3948 5536 5460
rect 5216 3892 5244 3948
rect 5300 3892 5348 3948
rect 5404 3892 5452 3948
rect 5508 3892 5536 3948
rect 5216 3076 5536 3892
rect 5852 3332 5908 7756
rect 5852 3266 5908 3276
rect 9248 7812 9276 7868
rect 9332 7812 9380 7868
rect 9436 7812 9484 7868
rect 9540 7812 9568 7868
rect 9248 6300 9568 7812
rect 9248 6244 9276 6300
rect 9332 6244 9380 6300
rect 9436 6244 9484 6300
rect 9540 6244 9568 6300
rect 9248 4732 9568 6244
rect 9248 4676 9276 4732
rect 9332 4676 9380 4732
rect 9436 4676 9484 4732
rect 9540 4676 9568 4732
rect 9248 3164 9568 4676
rect 9248 3108 9276 3164
rect 9332 3108 9380 3164
rect 9436 3108 9484 3164
rect 9540 3108 9568 3164
rect 9248 3076 9568 3108
rect 13280 11788 13600 13300
rect 13280 11732 13308 11788
rect 13364 11732 13412 11788
rect 13468 11732 13516 11788
rect 13572 11732 13600 11788
rect 13280 10220 13600 11732
rect 13280 10164 13308 10220
rect 13364 10164 13412 10220
rect 13468 10164 13516 10220
rect 13572 10164 13600 10220
rect 13280 8652 13600 10164
rect 13280 8596 13308 8652
rect 13364 8596 13412 8652
rect 13468 8596 13516 8652
rect 13572 8596 13600 8652
rect 13280 7084 13600 8596
rect 13280 7028 13308 7084
rect 13364 7028 13412 7084
rect 13468 7028 13516 7084
rect 13572 7028 13600 7084
rect 13280 5516 13600 7028
rect 13280 5460 13308 5516
rect 13364 5460 13412 5516
rect 13468 5460 13516 5516
rect 13572 5460 13600 5516
rect 13280 3948 13600 5460
rect 13280 3892 13308 3948
rect 13364 3892 13412 3948
rect 13468 3892 13516 3948
rect 13572 3892 13600 3948
rect 13280 3076 13600 3892
rect 17312 17276 17632 18788
rect 20860 19348 20916 19358
rect 17312 17220 17340 17276
rect 17396 17220 17444 17276
rect 17500 17220 17548 17276
rect 17604 17220 17632 17276
rect 17312 15708 17632 17220
rect 20188 18564 20244 18574
rect 17312 15652 17340 15708
rect 17396 15652 17444 15708
rect 17500 15652 17548 15708
rect 17604 15652 17632 15708
rect 17312 14140 17632 15652
rect 19292 16100 19348 16110
rect 19292 14420 19348 16044
rect 19628 15316 19684 15326
rect 19628 14868 19684 15260
rect 20188 15148 20244 18508
rect 19628 14802 19684 14812
rect 20076 15092 20244 15148
rect 19292 14354 19348 14364
rect 19628 14644 19684 14654
rect 17312 14084 17340 14140
rect 17396 14084 17444 14140
rect 17500 14084 17548 14140
rect 17604 14084 17632 14140
rect 17312 12572 17632 14084
rect 19068 14196 19124 14206
rect 19068 12964 19124 14140
rect 19628 13188 19684 14588
rect 19628 13122 19684 13132
rect 20076 13188 20132 15092
rect 20860 13412 20916 19292
rect 20860 13346 20916 13356
rect 21344 18060 21664 19572
rect 21344 18004 21372 18060
rect 21428 18004 21476 18060
rect 21532 18004 21580 18060
rect 21636 18004 21664 18060
rect 21344 16492 21664 18004
rect 21344 16436 21372 16492
rect 21428 16436 21476 16492
rect 21532 16436 21580 16492
rect 21636 16436 21664 16492
rect 21344 14924 21664 16436
rect 21344 14868 21372 14924
rect 21428 14868 21476 14924
rect 21532 14868 21580 14924
rect 21636 14868 21664 14924
rect 21344 13356 21664 14868
rect 20076 13122 20132 13132
rect 21344 13300 21372 13356
rect 21428 13300 21476 13356
rect 21532 13300 21580 13356
rect 21636 13300 21664 13356
rect 19068 12898 19124 12908
rect 17312 12516 17340 12572
rect 17396 12516 17444 12572
rect 17500 12516 17548 12572
rect 17604 12516 17632 12572
rect 17312 11004 17632 12516
rect 17312 10948 17340 11004
rect 17396 10948 17444 11004
rect 17500 10948 17548 11004
rect 17604 10948 17632 11004
rect 17312 9436 17632 10948
rect 17312 9380 17340 9436
rect 17396 9380 17444 9436
rect 17500 9380 17548 9436
rect 17604 9380 17632 9436
rect 17312 7868 17632 9380
rect 17312 7812 17340 7868
rect 17396 7812 17444 7868
rect 17500 7812 17548 7868
rect 17604 7812 17632 7868
rect 17312 6300 17632 7812
rect 17312 6244 17340 6300
rect 17396 6244 17444 6300
rect 17500 6244 17548 6300
rect 17604 6244 17632 6300
rect 17312 4732 17632 6244
rect 17312 4676 17340 4732
rect 17396 4676 17444 4732
rect 17500 4676 17548 4732
rect 17604 4676 17632 4732
rect 17312 3164 17632 4676
rect 17312 3108 17340 3164
rect 17396 3108 17444 3164
rect 17500 3108 17548 3164
rect 17604 3108 17632 3164
rect 17312 3076 17632 3108
rect 21344 11788 21664 13300
rect 25228 12180 25284 20188
rect 25228 12114 25284 12124
rect 25376 18844 25696 20356
rect 25788 21140 25844 21150
rect 25788 20244 25844 21084
rect 25788 20178 25844 20188
rect 26572 20356 26628 20366
rect 25376 18788 25404 18844
rect 25460 18788 25508 18844
rect 25564 18788 25612 18844
rect 25668 18788 25696 18844
rect 26572 18900 26628 20300
rect 26572 18834 26628 18844
rect 25376 17276 25696 18788
rect 26796 17668 26852 22988
rect 27020 22148 27076 22158
rect 26796 17602 26852 17612
rect 26908 21140 26964 21150
rect 26908 20132 26964 21084
rect 25376 17220 25404 17276
rect 25460 17220 25508 17276
rect 25564 17220 25612 17276
rect 25668 17220 25696 17276
rect 25376 15708 25696 17220
rect 25376 15652 25404 15708
rect 25460 15652 25508 15708
rect 25564 15652 25612 15708
rect 25668 15652 25696 15708
rect 25376 14140 25696 15652
rect 25376 14084 25404 14140
rect 25460 14084 25508 14140
rect 25564 14084 25612 14140
rect 25668 14084 25696 14140
rect 25900 15428 25956 15438
rect 25900 14196 25956 15372
rect 25900 14130 25956 14140
rect 25376 12572 25696 14084
rect 26908 14084 26964 20076
rect 27020 19908 27076 22092
rect 27244 21476 27300 21486
rect 27244 20356 27300 21420
rect 27244 20290 27300 20300
rect 27020 19842 27076 19852
rect 27244 20020 27300 20030
rect 27244 18900 27300 19964
rect 27244 18834 27300 18844
rect 28252 19236 28308 19246
rect 27804 18788 27860 18798
rect 27804 18452 27860 18732
rect 27804 18386 27860 18396
rect 27020 17332 27076 17342
rect 27020 16100 27076 17276
rect 27020 16034 27076 16044
rect 26908 14018 26964 14028
rect 27020 15764 27076 15774
rect 25376 12516 25404 12572
rect 25460 12516 25508 12572
rect 25564 12516 25612 12572
rect 25668 12516 25696 12572
rect 21344 11732 21372 11788
rect 21428 11732 21476 11788
rect 21532 11732 21580 11788
rect 21636 11732 21664 11788
rect 21344 10220 21664 11732
rect 21344 10164 21372 10220
rect 21428 10164 21476 10220
rect 21532 10164 21580 10220
rect 21636 10164 21664 10220
rect 21344 8652 21664 10164
rect 21344 8596 21372 8652
rect 21428 8596 21476 8652
rect 21532 8596 21580 8652
rect 21636 8596 21664 8652
rect 21344 7084 21664 8596
rect 25376 11004 25696 12516
rect 25376 10948 25404 11004
rect 25460 10948 25508 11004
rect 25564 10948 25612 11004
rect 25668 10948 25696 11004
rect 25376 9436 25696 10948
rect 25376 9380 25404 9436
rect 25460 9380 25508 9436
rect 25564 9380 25612 9436
rect 25668 9380 25696 9436
rect 25376 7868 25696 9380
rect 21344 7028 21372 7084
rect 21428 7028 21476 7084
rect 21532 7028 21580 7084
rect 21636 7028 21664 7084
rect 21344 5516 21664 7028
rect 21756 7812 21812 7822
rect 21756 5684 21812 7756
rect 21756 5618 21812 5628
rect 23324 7812 23380 7822
rect 21344 5460 21372 5516
rect 21428 5460 21476 5516
rect 21532 5460 21580 5516
rect 21636 5460 21664 5516
rect 23324 5572 23380 7756
rect 25376 7812 25404 7868
rect 25460 7812 25508 7868
rect 25564 7812 25612 7868
rect 25668 7812 25696 7868
rect 23548 7588 23604 7598
rect 23548 5908 23604 7532
rect 23548 5842 23604 5852
rect 24220 6916 24276 6926
rect 23324 5506 23380 5516
rect 21344 3948 21664 5460
rect 24220 5460 24276 6860
rect 24220 5394 24276 5404
rect 24444 6356 24500 6366
rect 24444 4564 24500 6300
rect 25376 6300 25696 7812
rect 25376 6244 25404 6300
rect 25460 6244 25508 6300
rect 25564 6244 25612 6300
rect 25668 6244 25696 6300
rect 24780 5908 24836 5918
rect 24780 5124 24836 5852
rect 24780 5058 24836 5068
rect 24444 4498 24500 4508
rect 25376 4732 25696 6244
rect 26684 7588 26740 7598
rect 26684 5124 26740 7532
rect 27020 7588 27076 15708
rect 28252 13972 28308 19180
rect 28364 18788 28420 25228
rect 28588 25284 28644 25294
rect 28588 21140 28644 25228
rect 28700 23156 28756 30492
rect 28924 25396 28980 31948
rect 29408 30604 29728 31420
rect 29408 30548 29436 30604
rect 29492 30548 29540 30604
rect 29596 30548 29644 30604
rect 29700 30548 29728 30604
rect 29408 29036 29728 30548
rect 33440 31388 33760 31420
rect 33440 31332 33468 31388
rect 33524 31332 33572 31388
rect 33628 31332 33676 31388
rect 33732 31332 33760 31388
rect 33440 29820 33760 31332
rect 33440 29764 33468 29820
rect 33524 29764 33572 29820
rect 33628 29764 33676 29820
rect 33732 29764 33760 29820
rect 29408 28980 29436 29036
rect 29492 28980 29540 29036
rect 29596 28980 29644 29036
rect 29700 28980 29728 29036
rect 29036 28532 29092 28542
rect 29036 26292 29092 28476
rect 29036 26226 29092 26236
rect 29408 27468 29728 28980
rect 29408 27412 29436 27468
rect 29492 27412 29540 27468
rect 29596 27412 29644 27468
rect 29700 27412 29728 27468
rect 28924 25330 28980 25340
rect 29408 25900 29728 27412
rect 29820 29092 29876 29102
rect 29820 26628 29876 29036
rect 33440 28252 33760 29764
rect 33440 28196 33468 28252
rect 33524 28196 33572 28252
rect 33628 28196 33676 28252
rect 33732 28196 33760 28252
rect 29820 26562 29876 26572
rect 30268 28084 30324 28094
rect 29408 25844 29436 25900
rect 29492 25844 29540 25900
rect 29596 25844 29644 25900
rect 29700 25844 29728 25900
rect 28700 23090 28756 23100
rect 29408 24332 29728 25844
rect 29408 24276 29436 24332
rect 29492 24276 29540 24332
rect 29596 24276 29644 24332
rect 29700 24276 29728 24332
rect 28588 20098 28644 21084
rect 29408 22764 29728 24276
rect 29408 22708 29436 22764
rect 29492 22708 29540 22764
rect 29596 22708 29644 22764
rect 29700 22708 29728 22764
rect 29408 21196 29728 22708
rect 29408 21140 29436 21196
rect 29492 21140 29540 21196
rect 29596 21140 29644 21196
rect 29700 21140 29728 21196
rect 28476 20042 28644 20098
rect 29148 20468 29204 20478
rect 28476 19236 28532 20042
rect 29148 20020 29204 20412
rect 29148 19954 29204 19964
rect 28476 19170 28532 19180
rect 29036 19908 29092 19918
rect 28364 18722 28420 18732
rect 28476 18900 28532 18910
rect 28476 17444 28532 18844
rect 28476 17378 28532 17388
rect 28700 16996 28756 17006
rect 28700 15428 28756 16940
rect 28700 15362 28756 15372
rect 28588 14980 28644 14990
rect 28588 14196 28644 14924
rect 28588 14130 28644 14140
rect 28252 13906 28308 13916
rect 29036 11844 29092 19852
rect 29408 19628 29728 21140
rect 29408 19572 29436 19628
rect 29492 19572 29540 19628
rect 29596 19572 29644 19628
rect 29700 19572 29728 19628
rect 29148 18452 29204 18462
rect 29148 16100 29204 18396
rect 29148 12740 29204 16044
rect 29148 12674 29204 12684
rect 29408 18060 29728 19572
rect 29408 18004 29436 18060
rect 29492 18004 29540 18060
rect 29596 18004 29644 18060
rect 29700 18004 29728 18060
rect 29408 16492 29728 18004
rect 29408 16436 29436 16492
rect 29492 16436 29540 16492
rect 29596 16436 29644 16492
rect 29700 16436 29728 16492
rect 29408 14924 29728 16436
rect 30268 20132 30324 28028
rect 29408 14868 29436 14924
rect 29492 14868 29540 14924
rect 29596 14868 29644 14924
rect 29700 14868 29728 14924
rect 29408 13356 29728 14868
rect 29408 13300 29436 13356
rect 29492 13300 29540 13356
rect 29596 13300 29644 13356
rect 29700 13300 29728 13356
rect 29036 11778 29092 11788
rect 29408 11788 29728 13300
rect 27020 6916 27076 7532
rect 29408 11732 29436 11788
rect 29492 11732 29540 11788
rect 29596 11732 29644 11788
rect 29700 11732 29728 11788
rect 29408 10220 29728 11732
rect 30156 15764 30212 15774
rect 30156 11508 30212 15708
rect 30156 11442 30212 11452
rect 29408 10164 29436 10220
rect 29492 10164 29540 10220
rect 29596 10164 29644 10220
rect 29700 10164 29728 10220
rect 29408 8652 29728 10164
rect 30268 9268 30324 20076
rect 33440 26684 33760 28196
rect 33440 26628 33468 26684
rect 33524 26628 33572 26684
rect 33628 26628 33676 26684
rect 33732 26628 33760 26684
rect 33440 25116 33760 26628
rect 33440 25060 33468 25116
rect 33524 25060 33572 25116
rect 33628 25060 33676 25116
rect 33732 25060 33760 25116
rect 33440 23548 33760 25060
rect 33440 23492 33468 23548
rect 33524 23492 33572 23548
rect 33628 23492 33676 23548
rect 33732 23492 33760 23548
rect 33440 21980 33760 23492
rect 33440 21924 33468 21980
rect 33524 21924 33572 21980
rect 33628 21924 33676 21980
rect 33732 21924 33760 21980
rect 33440 20412 33760 21924
rect 33440 20356 33468 20412
rect 33524 20356 33572 20412
rect 33628 20356 33676 20412
rect 33732 20356 33760 20412
rect 33440 18844 33760 20356
rect 33440 18788 33468 18844
rect 33524 18788 33572 18844
rect 33628 18788 33676 18844
rect 33732 18788 33760 18844
rect 30940 18452 30996 18462
rect 30940 15092 30996 18396
rect 30940 15026 30996 15036
rect 33440 17276 33760 18788
rect 33440 17220 33468 17276
rect 33524 17220 33572 17276
rect 33628 17220 33676 17276
rect 33732 17220 33760 17276
rect 33440 15708 33760 17220
rect 33440 15652 33468 15708
rect 33524 15652 33572 15708
rect 33628 15652 33676 15708
rect 33732 15652 33760 15708
rect 30268 9202 30324 9212
rect 33440 14140 33760 15652
rect 33440 14084 33468 14140
rect 33524 14084 33572 14140
rect 33628 14084 33676 14140
rect 33732 14084 33760 14140
rect 33440 12572 33760 14084
rect 33440 12516 33468 12572
rect 33524 12516 33572 12572
rect 33628 12516 33676 12572
rect 33732 12516 33760 12572
rect 33440 11004 33760 12516
rect 33440 10948 33468 11004
rect 33524 10948 33572 11004
rect 33628 10948 33676 11004
rect 33732 10948 33760 11004
rect 33440 9436 33760 10948
rect 33440 9380 33468 9436
rect 33524 9380 33572 9436
rect 33628 9380 33676 9436
rect 33732 9380 33760 9436
rect 29408 8596 29436 8652
rect 29492 8596 29540 8652
rect 29596 8596 29644 8652
rect 29700 8596 29728 8652
rect 27020 6850 27076 6860
rect 27692 7140 27748 7150
rect 26684 5058 26740 5068
rect 25376 4676 25404 4732
rect 25460 4676 25508 4732
rect 25564 4676 25612 4732
rect 25668 4676 25696 4732
rect 21344 3892 21372 3948
rect 21428 3892 21476 3948
rect 21532 3892 21580 3948
rect 21636 3892 21664 3948
rect 21344 3076 21664 3892
rect 25376 3164 25696 4676
rect 27692 3556 27748 7084
rect 27692 3490 27748 3500
rect 29408 7084 29728 8596
rect 29408 7028 29436 7084
rect 29492 7028 29540 7084
rect 29596 7028 29644 7084
rect 29700 7028 29728 7084
rect 29408 5516 29728 7028
rect 29408 5460 29436 5516
rect 29492 5460 29540 5516
rect 29596 5460 29644 5516
rect 29700 5460 29728 5516
rect 29408 3948 29728 5460
rect 29408 3892 29436 3948
rect 29492 3892 29540 3948
rect 29596 3892 29644 3948
rect 29700 3892 29728 3948
rect 25376 3108 25404 3164
rect 25460 3108 25508 3164
rect 25564 3108 25612 3164
rect 25668 3108 25696 3164
rect 25376 3076 25696 3108
rect 29408 3076 29728 3892
rect 33440 7868 33760 9380
rect 33440 7812 33468 7868
rect 33524 7812 33572 7868
rect 33628 7812 33676 7868
rect 33732 7812 33760 7868
rect 33440 6300 33760 7812
rect 33440 6244 33468 6300
rect 33524 6244 33572 6300
rect 33628 6244 33676 6300
rect 33732 6244 33760 6300
rect 33440 4732 33760 6244
rect 33440 4676 33468 4732
rect 33524 4676 33572 4732
rect 33628 4676 33676 4732
rect 33732 4676 33760 4732
rect 33440 3164 33760 4676
rect 33440 3108 33468 3164
rect 33524 3108 33572 3164
rect 33628 3108 33676 3164
rect 33732 3108 33760 3164
rect 33440 3076 33760 3108
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0511_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 30464 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0512_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 30464 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0513_
timestamp 1698175906
transform 1 0 27664 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0514_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0515_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23632 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0516_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24752 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0517_
timestamp 1698175906
transform 1 0 29792 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0518_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28784 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0519_
timestamp 1698175906
transform 1 0 29680 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0520_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 25760 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0521_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23744 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0522_
timestamp 1698175906
transform 1 0 25424 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0523_
timestamp 1698175906
transform -1 0 29904 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0524_
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0525_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24752 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0526_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23632 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0527_
timestamp 1698175906
transform -1 0 21952 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0528_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0529_
timestamp 1698175906
transform -1 0 26208 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0530_
timestamp 1698175906
transform -1 0 23072 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0531_
timestamp 1698175906
transform 1 0 21168 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0532_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28560 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0533_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0534_
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0535_
timestamp 1698175906
transform -1 0 33376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0536_
timestamp 1698175906
transform -1 0 32704 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0537_
timestamp 1698175906
transform -1 0 33264 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0538_
timestamp 1698175906
transform -1 0 22848 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0539_
timestamp 1698175906
transform -1 0 32704 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0540_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0541_
timestamp 1698175906
transform -1 0 32256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0542_
timestamp 1698175906
transform -1 0 27664 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0543_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 25200 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0544_
timestamp 1698175906
transform -1 0 24864 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0545_
timestamp 1698175906
transform 1 0 21840 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0546_
timestamp 1698175906
transform 1 0 21952 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0547_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23856 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0548_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23408 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0549_
timestamp 1698175906
transform -1 0 24864 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0550_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26432 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0551_
timestamp 1698175906
transform 1 0 21952 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0552_
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0553_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0554_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 29792 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0555_
timestamp 1698175906
transform -1 0 30800 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0556_
timestamp 1698175906
transform 1 0 25536 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0557_
timestamp 1698175906
transform -1 0 29680 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0558_
timestamp 1698175906
transform -1 0 33376 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0559_
timestamp 1698175906
transform -1 0 25648 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0560_
timestamp 1698175906
transform -1 0 28784 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0561_
timestamp 1698175906
transform -1 0 26768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0562_
timestamp 1698175906
transform 1 0 26432 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0563_
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0564_
timestamp 1698175906
transform 1 0 25984 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0565_
timestamp 1698175906
transform -1 0 26432 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0566_
timestamp 1698175906
transform 1 0 21392 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0567_
timestamp 1698175906
transform 1 0 32032 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0568_
timestamp 1698175906
transform -1 0 23520 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0569_
timestamp 1698175906
transform 1 0 26656 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0570_
timestamp 1698175906
transform -1 0 27776 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0571_
timestamp 1698175906
transform 1 0 23632 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0572_
timestamp 1698175906
transform -1 0 22736 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0573_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0574_
timestamp 1698175906
transform -1 0 21840 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0575_
timestamp 1698175906
transform -1 0 24080 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0576_
timestamp 1698175906
transform -1 0 24640 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0577_
timestamp 1698175906
transform 1 0 24864 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0578_
timestamp 1698175906
transform -1 0 24080 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0579_
timestamp 1698175906
transform 1 0 22736 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0580_
timestamp 1698175906
transform -1 0 23520 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0581_
timestamp 1698175906
transform 1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0582_
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0583_
timestamp 1698175906
transform -1 0 28000 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0584_
timestamp 1698175906
transform -1 0 27552 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0585_
timestamp 1698175906
transform 1 0 28000 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0586_
timestamp 1698175906
transform -1 0 21616 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0587_
timestamp 1698175906
transform -1 0 21056 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0588_
timestamp 1698175906
transform -1 0 21504 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0589_
timestamp 1698175906
transform -1 0 19600 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0590_
timestamp 1698175906
transform 1 0 11760 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0591_
timestamp 1698175906
transform 1 0 11872 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0592_
timestamp 1698175906
transform 1 0 19600 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0593_
timestamp 1698175906
transform -1 0 22176 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0594_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0595_
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0596_
timestamp 1698175906
transform -1 0 18256 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0597_
timestamp 1698175906
transform -1 0 27440 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0598_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24080 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0599_
timestamp 1698175906
transform 1 0 25200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0600_
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0601_
timestamp 1698175906
transform -1 0 33376 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0602_
timestamp 1698175906
transform -1 0 26768 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0603_
timestamp 1698175906
transform -1 0 28784 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0604_
timestamp 1698175906
transform -1 0 28672 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0605_
timestamp 1698175906
transform 1 0 27552 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0606_
timestamp 1698175906
transform -1 0 33376 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0607_
timestamp 1698175906
transform -1 0 23296 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _0608_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32704 0 -1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0609_
timestamp 1698175906
transform -1 0 33376 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0610_
timestamp 1698175906
transform -1 0 33040 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0611_
timestamp 1698175906
transform 1 0 22512 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _0612_
timestamp 1698175906
transform -1 0 32704 0 -1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0613_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 30240 0 -1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0614_
timestamp 1698175906
transform -1 0 33376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0615_
timestamp 1698175906
transform -1 0 30464 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0616_
timestamp 1698175906
transform -1 0 33376 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0617_
timestamp 1698175906
transform -1 0 29568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0618_
timestamp 1698175906
transform 1 0 28224 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0619_
timestamp 1698175906
transform 1 0 31472 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _0620_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 29456 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0621_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32592 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0622_
timestamp 1698175906
transform 1 0 28336 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0623_
timestamp 1698175906
transform 1 0 29904 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _0624_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 29232 0 1 17248
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0625_
timestamp 1698175906
transform 1 0 18256 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0626_
timestamp 1698175906
transform -1 0 17248 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0627_
timestamp 1698175906
transform -1 0 21840 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0628_
timestamp 1698175906
transform -1 0 23744 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0629_
timestamp 1698175906
transform -1 0 21840 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0630_
timestamp 1698175906
transform -1 0 18368 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0631_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0632_
timestamp 1698175906
transform 1 0 18816 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0633_
timestamp 1698175906
transform 1 0 18368 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0634_
timestamp 1698175906
transform 1 0 18368 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0635_
timestamp 1698175906
transform -1 0 18368 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0636_
timestamp 1698175906
transform 1 0 19264 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0637_
timestamp 1698175906
transform 1 0 18256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0638_
timestamp 1698175906
transform 1 0 21952 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0639_
timestamp 1698175906
transform 1 0 23856 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0640_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28336 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0641_
timestamp 1698175906
transform 1 0 22736 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0642_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23408 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0643_
timestamp 1698175906
transform 1 0 6272 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0644_
timestamp 1698175906
transform 1 0 7840 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0645_
timestamp 1698175906
transform -1 0 3024 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0646_
timestamp 1698175906
transform 1 0 5600 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0647_
timestamp 1698175906
transform 1 0 4816 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0648_
timestamp 1698175906
transform 1 0 2800 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0649_
timestamp 1698175906
transform -1 0 3920 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0650_
timestamp 1698175906
transform 1 0 3920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0651_
timestamp 1698175906
transform 1 0 3024 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0652_
timestamp 1698175906
transform 1 0 23744 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0653_
timestamp 1698175906
transform -1 0 30128 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0654_
timestamp 1698175906
transform -1 0 26544 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0655_
timestamp 1698175906
transform -1 0 11200 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0656_
timestamp 1698175906
transform 1 0 11424 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0657_
timestamp 1698175906
transform 1 0 11200 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0658_
timestamp 1698175906
transform 1 0 10528 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0659_
timestamp 1698175906
transform -1 0 25536 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0660_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25536 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0661_
timestamp 1698175906
transform -1 0 14112 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0662_
timestamp 1698175906
transform -1 0 12096 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0663_
timestamp 1698175906
transform 1 0 9968 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0664_
timestamp 1698175906
transform 1 0 12096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0665_
timestamp 1698175906
transform -1 0 12768 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0666_
timestamp 1698175906
transform 1 0 10640 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0667_
timestamp 1698175906
transform -1 0 12656 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0668_
timestamp 1698175906
transform 1 0 10080 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0669_
timestamp 1698175906
transform 1 0 10304 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0670_
timestamp 1698175906
transform -1 0 9968 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0671_
timestamp 1698175906
transform 1 0 9520 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0672_
timestamp 1698175906
transform 1 0 12096 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0673_
timestamp 1698175906
transform 1 0 13104 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0674_
timestamp 1698175906
transform 1 0 12432 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0675_
timestamp 1698175906
transform -1 0 13104 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0676_
timestamp 1698175906
transform 1 0 12880 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0677_
timestamp 1698175906
transform -1 0 15680 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0678_
timestamp 1698175906
transform 1 0 14112 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0679_
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0680_
timestamp 1698175906
transform 1 0 12992 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0681_
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0682_
timestamp 1698175906
transform -1 0 17472 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0683_
timestamp 1698175906
transform -1 0 19600 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0684_
timestamp 1698175906
transform -1 0 17024 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0685_
timestamp 1698175906
transform -1 0 19488 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0686_
timestamp 1698175906
transform 1 0 19488 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0687_
timestamp 1698175906
transform -1 0 19040 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0688_
timestamp 1698175906
transform -1 0 23296 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0689_
timestamp 1698175906
transform 1 0 25872 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0690_
timestamp 1698175906
transform -1 0 23968 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0691_
timestamp 1698175906
transform -1 0 21504 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0692_
timestamp 1698175906
transform -1 0 28336 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0693_
timestamp 1698175906
transform -1 0 25760 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0694_
timestamp 1698175906
transform -1 0 20832 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0695_
timestamp 1698175906
transform -1 0 18704 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0696_
timestamp 1698175906
transform -1 0 19936 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0697_
timestamp 1698175906
transform -1 0 15456 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0698_
timestamp 1698175906
transform 1 0 13664 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0699_
timestamp 1698175906
transform -1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0700_
timestamp 1698175906
transform -1 0 24080 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0701_
timestamp 1698175906
transform -1 0 23408 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0702_
timestamp 1698175906
transform 1 0 16688 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0703_
timestamp 1698175906
transform 1 0 15456 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0704_
timestamp 1698175906
transform -1 0 16240 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0705_
timestamp 1698175906
transform -1 0 24864 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0706_
timestamp 1698175906
transform -1 0 23968 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0707_
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0708_
timestamp 1698175906
transform -1 0 18144 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0709_
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0710_
timestamp 1698175906
transform -1 0 27104 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0711_
timestamp 1698175906
transform -1 0 24528 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0712_
timestamp 1698175906
transform 1 0 19264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0713_
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0714_
timestamp 1698175906
transform 1 0 19824 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0715_
timestamp 1698175906
transform 1 0 19936 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0716_
timestamp 1698175906
transform 1 0 23072 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0717_
timestamp 1698175906
transform 1 0 24080 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0718_
timestamp 1698175906
transform -1 0 28784 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0719_
timestamp 1698175906
transform 1 0 24528 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0720_
timestamp 1698175906
transform 1 0 24080 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0721_
timestamp 1698175906
transform 1 0 23744 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0722_
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0723_
timestamp 1698175906
transform 1 0 23184 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0724_
timestamp 1698175906
transform -1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0725_
timestamp 1698175906
transform -1 0 27888 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0726_
timestamp 1698175906
transform 1 0 25984 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0727_
timestamp 1698175906
transform 1 0 26880 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0728_
timestamp 1698175906
transform 1 0 25984 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0729_
timestamp 1698175906
transform -1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0730_
timestamp 1698175906
transform 1 0 29120 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0731_
timestamp 1698175906
transform 1 0 27888 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0732_
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0733_
timestamp 1698175906
transform -1 0 25984 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0734_
timestamp 1698175906
transform -1 0 33376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0735_
timestamp 1698175906
transform 1 0 28896 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0736_
timestamp 1698175906
transform 1 0 29008 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0737_
timestamp 1698175906
transform -1 0 13104 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0738_
timestamp 1698175906
transform 1 0 22400 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0739_
timestamp 1698175906
transform -1 0 29344 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0740_
timestamp 1698175906
transform -1 0 28672 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0741_
timestamp 1698175906
transform -1 0 29680 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0742_
timestamp 1698175906
transform -1 0 28224 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0743_
timestamp 1698175906
transform -1 0 28896 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0744_
timestamp 1698175906
transform 1 0 26768 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0745_
timestamp 1698175906
transform -1 0 25872 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0746_
timestamp 1698175906
transform 1 0 27328 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0747_
timestamp 1698175906
transform -1 0 27216 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0748_
timestamp 1698175906
transform -1 0 21952 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0749_
timestamp 1698175906
transform -1 0 26544 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0750_
timestamp 1698175906
transform 1 0 22064 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0751_
timestamp 1698175906
transform 1 0 21504 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0752_
timestamp 1698175906
transform -1 0 27328 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0753_
timestamp 1698175906
transform -1 0 23632 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0754_
timestamp 1698175906
transform 1 0 21952 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0755_
timestamp 1698175906
transform 1 0 23296 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0756_
timestamp 1698175906
transform 1 0 22400 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0757_
timestamp 1698175906
transform -1 0 24752 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0758_
timestamp 1698175906
transform 1 0 22960 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0759_
timestamp 1698175906
transform -1 0 24752 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0760_
timestamp 1698175906
transform 1 0 24304 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0761_
timestamp 1698175906
transform -1 0 26656 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0762_
timestamp 1698175906
transform 1 0 25200 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0763_
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0764_
timestamp 1698175906
transform 1 0 25984 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0765_
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0766_
timestamp 1698175906
transform 1 0 28448 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0767_
timestamp 1698175906
transform 1 0 27328 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0768_
timestamp 1698175906
transform 1 0 27104 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0769_
timestamp 1698175906
transform -1 0 28336 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0770_
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0771_
timestamp 1698175906
transform 1 0 29456 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0772_
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0773_
timestamp 1698175906
transform 1 0 28336 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0774_
timestamp 1698175906
transform -1 0 31248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0775_
timestamp 1698175906
transform -1 0 32144 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0776_
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0777_
timestamp 1698175906
transform 1 0 27776 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0778_
timestamp 1698175906
transform -1 0 30912 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0779_
timestamp 1698175906
transform -1 0 31808 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0780_
timestamp 1698175906
transform -1 0 32368 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0781_
timestamp 1698175906
transform 1 0 28224 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0782_
timestamp 1698175906
transform -1 0 31472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0783_
timestamp 1698175906
transform 1 0 9744 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0784_
timestamp 1698175906
transform -1 0 31696 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0785_
timestamp 1698175906
transform -1 0 32592 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0786_
timestamp 1698175906
transform -1 0 28784 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0787_
timestamp 1698175906
transform -1 0 33376 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0788_
timestamp 1698175906
transform -1 0 18592 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0789_
timestamp 1698175906
transform -1 0 24864 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0790_
timestamp 1698175906
transform -1 0 19040 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0791_
timestamp 1698175906
transform 1 0 19712 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0792_
timestamp 1698175906
transform -1 0 21840 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0793_
timestamp 1698175906
transform -1 0 15568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0794_
timestamp 1698175906
transform -1 0 20832 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0795_
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0796_
timestamp 1698175906
transform 1 0 7952 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0797_
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0798_
timestamp 1698175906
transform 1 0 15456 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0799_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0800_
timestamp 1698175906
transform 1 0 19152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0801_
timestamp 1698175906
transform -1 0 20944 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0802_
timestamp 1698175906
transform 1 0 18592 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0803_
timestamp 1698175906
transform -1 0 18368 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0804_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20272 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0805_
timestamp 1698175906
transform -1 0 14672 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0806_
timestamp 1698175906
transform 1 0 11088 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0807_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19376 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0808_
timestamp 1698175906
transform 1 0 13216 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0809_
timestamp 1698175906
transform 1 0 16912 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0810_
timestamp 1698175906
transform 1 0 18816 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0811_
timestamp 1698175906
transform -1 0 11760 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0812_
timestamp 1698175906
transform 1 0 8064 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0813_
timestamp 1698175906
transform -1 0 19600 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0814_
timestamp 1698175906
transform -1 0 20496 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0815_
timestamp 1698175906
transform -1 0 18704 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0816_
timestamp 1698175906
transform 1 0 16576 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0817_
timestamp 1698175906
transform -1 0 14672 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0818_
timestamp 1698175906
transform 1 0 11424 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0819_
timestamp 1698175906
transform 1 0 26544 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0820_
timestamp 1698175906
transform -1 0 11872 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0821_
timestamp 1698175906
transform 1 0 15904 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0822_
timestamp 1698175906
transform 1 0 26096 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0823_
timestamp 1698175906
transform 1 0 17248 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0824_
timestamp 1698175906
transform -1 0 20384 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0825_
timestamp 1698175906
transform -1 0 18368 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0826_
timestamp 1698175906
transform -1 0 26432 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0827_
timestamp 1698175906
transform -1 0 33376 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0828_
timestamp 1698175906
transform 1 0 22064 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0829_
timestamp 1698175906
transform 1 0 22624 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0830_
timestamp 1698175906
transform -1 0 21840 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0831_
timestamp 1698175906
transform 1 0 29232 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0832_
timestamp 1698175906
transform -1 0 20944 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0833_
timestamp 1698175906
transform -1 0 19712 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0834_
timestamp 1698175906
transform 1 0 15344 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0835_
timestamp 1698175906
transform -1 0 15120 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0836_
timestamp 1698175906
transform -1 0 11088 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0837_
timestamp 1698175906
transform 1 0 10416 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0838_
timestamp 1698175906
transform 1 0 10080 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0839_
timestamp 1698175906
transform -1 0 7392 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0840_
timestamp 1698175906
transform 1 0 7392 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0841_
timestamp 1698175906
transform -1 0 8848 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0842_
timestamp 1698175906
transform -1 0 8288 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0843_
timestamp 1698175906
transform 1 0 6160 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0844_
timestamp 1698175906
transform -1 0 8512 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0845_
timestamp 1698175906
transform 1 0 6496 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0846_
timestamp 1698175906
transform -1 0 6944 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0847_
timestamp 1698175906
transform -1 0 7280 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0848_
timestamp 1698175906
transform -1 0 7280 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0849_
timestamp 1698175906
transform -1 0 6384 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0850_
timestamp 1698175906
transform -1 0 5600 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0851_
timestamp 1698175906
transform -1 0 6160 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0852_
timestamp 1698175906
transform 1 0 3696 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0853_
timestamp 1698175906
transform 1 0 4256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0854_
timestamp 1698175906
transform -1 0 6496 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0855_
timestamp 1698175906
transform -1 0 3920 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0856_
timestamp 1698175906
transform -1 0 5488 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0857_
timestamp 1698175906
transform -1 0 4928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0858_
timestamp 1698175906
transform -1 0 5376 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0859_
timestamp 1698175906
transform 1 0 2800 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0860_
timestamp 1698175906
transform 1 0 3920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0861_
timestamp 1698175906
transform -1 0 4816 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0862_
timestamp 1698175906
transform -1 0 6048 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0863_
timestamp 1698175906
transform -1 0 7952 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0864_
timestamp 1698175906
transform 1 0 3920 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0865_
timestamp 1698175906
transform 1 0 6496 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0866_
timestamp 1698175906
transform 1 0 4928 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0867_
timestamp 1698175906
transform -1 0 6048 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0868_
timestamp 1698175906
transform -1 0 5712 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0869_
timestamp 1698175906
transform -1 0 8736 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0870_
timestamp 1698175906
transform -1 0 7840 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0871_
timestamp 1698175906
transform 1 0 5936 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0872_
timestamp 1698175906
transform 1 0 6160 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0873_
timestamp 1698175906
transform -1 0 9296 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0874_
timestamp 1698175906
transform -1 0 8400 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0875_
timestamp 1698175906
transform 1 0 7840 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0876_
timestamp 1698175906
transform -1 0 11200 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0877_
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0878_
timestamp 1698175906
transform 1 0 10416 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0879_
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0880_
timestamp 1698175906
transform 1 0 11536 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0881_
timestamp 1698175906
transform -1 0 12880 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0882_
timestamp 1698175906
transform -1 0 11760 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0883_
timestamp 1698175906
transform -1 0 11536 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0884_
timestamp 1698175906
transform -1 0 16352 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0885_
timestamp 1698175906
transform 1 0 12880 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0886_
timestamp 1698175906
transform 1 0 13440 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0887_
timestamp 1698175906
transform -1 0 15792 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0888_
timestamp 1698175906
transform 1 0 13440 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0889_
timestamp 1698175906
transform -1 0 15232 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0890_
timestamp 1698175906
transform -1 0 15568 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0891_
timestamp 1698175906
transform 1 0 13440 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0892_
timestamp 1698175906
transform 1 0 13888 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0893_
timestamp 1698175906
transform 1 0 14000 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0894_
timestamp 1698175906
transform -1 0 24304 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0895_
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0896_
timestamp 1698175906
transform -1 0 13104 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0897_
timestamp 1698175906
transform -1 0 7504 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0898_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0899_
timestamp 1698175906
transform -1 0 14448 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0900_
timestamp 1698175906
transform 1 0 8176 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0901_
timestamp 1698175906
transform 1 0 7056 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0902_
timestamp 1698175906
transform -1 0 12432 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0903_
timestamp 1698175906
transform -1 0 12320 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0904_
timestamp 1698175906
transform 1 0 5152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0905_
timestamp 1698175906
transform -1 0 5712 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0906_
timestamp 1698175906
transform -1 0 7952 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0907_
timestamp 1698175906
transform -1 0 8960 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0908_
timestamp 1698175906
transform -1 0 8960 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0909_
timestamp 1698175906
transform 1 0 7728 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0910_
timestamp 1698175906
transform 1 0 7504 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0911_
timestamp 1698175906
transform 1 0 7168 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0912_
timestamp 1698175906
transform 1 0 7392 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0913_
timestamp 1698175906
transform -1 0 10304 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0914_
timestamp 1698175906
transform -1 0 14896 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0915_
timestamp 1698175906
transform 1 0 4704 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0916_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4368 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0917_
timestamp 1698175906
transform 1 0 6160 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0918_
timestamp 1698175906
transform -1 0 11088 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0919_
timestamp 1698175906
transform 1 0 6160 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0920_
timestamp 1698175906
transform 1 0 7728 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0921_
timestamp 1698175906
transform -1 0 3136 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0922_
timestamp 1698175906
transform -1 0 7840 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0923_
timestamp 1698175906
transform -1 0 17136 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0924_
timestamp 1698175906
transform -1 0 7168 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0925_
timestamp 1698175906
transform -1 0 11872 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0926_
timestamp 1698175906
transform -1 0 6160 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0927_
timestamp 1698175906
transform -1 0 6608 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0928_
timestamp 1698175906
transform -1 0 7056 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0929_
timestamp 1698175906
transform -1 0 4256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0930_
timestamp 1698175906
transform 1 0 5600 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0931_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5936 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0932_
timestamp 1698175906
transform -1 0 7840 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0933_
timestamp 1698175906
transform -1 0 7728 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0934_
timestamp 1698175906
transform -1 0 7056 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0935_
timestamp 1698175906
transform -1 0 3584 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0936_
timestamp 1698175906
transform -1 0 10080 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0937_
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0938_
timestamp 1698175906
transform -1 0 9072 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0939_
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0940_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5712 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0941_
timestamp 1698175906
transform 1 0 4368 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0942_
timestamp 1698175906
transform -1 0 4368 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0943_
timestamp 1698175906
transform -1 0 9184 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0944_
timestamp 1698175906
transform 1 0 10528 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0945_
timestamp 1698175906
transform -1 0 10640 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0946_
timestamp 1698175906
transform -1 0 11200 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0947_
timestamp 1698175906
transform 1 0 11200 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0948_
timestamp 1698175906
transform -1 0 9856 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0949_
timestamp 1698175906
transform 1 0 9408 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0950_
timestamp 1698175906
transform 1 0 9856 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0951_
timestamp 1698175906
transform 1 0 10864 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0952_
timestamp 1698175906
transform -1 0 11648 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0953_
timestamp 1698175906
transform -1 0 11536 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0954_
timestamp 1698175906
transform -1 0 11424 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0955_
timestamp 1698175906
transform -1 0 10192 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0956_
timestamp 1698175906
transform -1 0 17136 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0957_
timestamp 1698175906
transform 1 0 6496 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0958_
timestamp 1698175906
transform 1 0 12208 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0959_
timestamp 1698175906
transform 1 0 15792 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0960_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14000 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0961_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15792 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0962_
timestamp 1698175906
transform -1 0 17472 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0963_
timestamp 1698175906
transform 1 0 10528 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0964_
timestamp 1698175906
transform 1 0 15792 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0965_
timestamp 1698175906
transform 1 0 12992 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0966_
timestamp 1698175906
transform 1 0 10752 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0967_
timestamp 1698175906
transform -1 0 15792 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0968_
timestamp 1698175906
transform -1 0 15344 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0969_
timestamp 1698175906
transform 1 0 13552 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0970_
timestamp 1698175906
transform 1 0 11648 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0971_
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0972_
timestamp 1698175906
transform -1 0 12992 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0973_
timestamp 1698175906
transform 1 0 9968 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0974_
timestamp 1698175906
transform -1 0 13104 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0975_
timestamp 1698175906
transform -1 0 12880 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0976_
timestamp 1698175906
transform 1 0 9184 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0977_
timestamp 1698175906
transform 1 0 13776 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0978_
timestamp 1698175906
transform -1 0 17024 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0979_
timestamp 1698175906
transform 1 0 12768 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0980_
timestamp 1698175906
transform 1 0 13552 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0981_
timestamp 1698175906
transform 1 0 14784 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0982_
timestamp 1698175906
transform 1 0 17360 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0983_
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0984_
timestamp 1698175906
transform 1 0 20272 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0985_
timestamp 1698175906
transform 1 0 19040 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0986_
timestamp 1698175906
transform 1 0 18032 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0987_
timestamp 1698175906
transform 1 0 20160 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0988_
timestamp 1698175906
transform 1 0 19040 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0989_
timestamp 1698175906
transform 1 0 14672 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0990_
timestamp 1698175906
transform -1 0 16464 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0991_
timestamp 1698175906
transform 1 0 19936 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0992_
timestamp 1698175906
transform 1 0 18032 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0993_
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0994_
timestamp 1698175906
transform 1 0 19264 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0995_
timestamp 1698175906
transform 1 0 20048 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0996_
timestamp 1698175906
transform 1 0 18368 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0997_
timestamp 1698175906
transform 1 0 19488 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0998_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16912 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0999_
timestamp 1698175906
transform 1 0 16016 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1000_
timestamp 1698175906
transform -1 0 19264 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1001_
timestamp 1698175906
transform 1 0 17136 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1002_
timestamp 1698175906
transform -1 0 7840 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1003_
timestamp 1698175906
transform 1 0 7504 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1004_
timestamp 1698175906
transform 1 0 6608 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1005_
timestamp 1698175906
transform 1 0 8512 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1006_
timestamp 1698175906
transform 1 0 7504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1007_
timestamp 1698175906
transform 1 0 6944 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1008_
timestamp 1698175906
transform 1 0 4592 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1009_
timestamp 1698175906
transform -1 0 9968 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1010_
timestamp 1698175906
transform -1 0 5712 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1011_
timestamp 1698175906
transform -1 0 9072 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1012_
timestamp 1698175906
transform -1 0 9296 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1013_
timestamp 1698175906
transform 1 0 6608 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1014_
timestamp 1698175906
transform 1 0 4928 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1015_
timestamp 1698175906
transform -1 0 6048 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1016_
timestamp 1698175906
transform 1 0 8064 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1017_
timestamp 1698175906
transform -1 0 5488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1018_
timestamp 1698175906
transform 1 0 1680 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1019_
timestamp 1698175906
transform -1 0 2800 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1020_
timestamp 1698175906
transform 1 0 5600 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1021_
timestamp 1698175906
transform 1 0 1792 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1022_
timestamp 1698175906
transform -1 0 4592 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1023_
timestamp 1698175906
transform 1 0 5488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1024_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1025_
timestamp 1698175906
transform -1 0 4816 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1026_
timestamp 1698175906
transform 1 0 9072 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1027_
timestamp 1698175906
transform -1 0 12656 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1028_
timestamp 1698175906
transform 1 0 8848 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1029_
timestamp 1698175906
transform -1 0 12656 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1030_
timestamp 1698175906
transform -1 0 15792 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1031_
timestamp 1698175906
transform 1 0 13440 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1032_
timestamp 1698175906
transform 1 0 15680 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1033_
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1034_
timestamp 1698175906
transform 1 0 12096 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1035_
timestamp 1698175906
transform 1 0 13552 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1036_
timestamp 1698175906
transform 1 0 16352 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1037_
timestamp 1698175906
transform 1 0 18816 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1038_
timestamp 1698175906
transform 1 0 21616 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1039_
timestamp 1698175906
transform 1 0 25200 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1040_
timestamp 1698175906
transform 1 0 25760 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1041_
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1042_
timestamp 1698175906
transform 1 0 17696 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1043_
timestamp 1698175906
transform 1 0 18816 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1044_
timestamp 1698175906
transform 1 0 20720 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1045_
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1046_
timestamp 1698175906
transform 1 0 28336 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1047_
timestamp 1698175906
transform -1 0 33376 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1048_
timestamp 1698175906
transform -1 0 33376 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1049_
timestamp 1698175906
transform -1 0 33376 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1050_
timestamp 1698175906
transform 1 0 22512 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1051_
timestamp 1698175906
transform 1 0 24640 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1052_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18592 0 -1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1053_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19376 0 -1 12544
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1054_
timestamp 1698175906
transform 1 0 13552 0 -1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1055_
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1056_
timestamp 1698175906
transform -1 0 28784 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1057_
timestamp 1698175906
transform -1 0 32704 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1058_
timestamp 1698175906
transform -1 0 33376 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1059_
timestamp 1698175906
transform 1 0 29456 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1060_
timestamp 1698175906
transform 1 0 16912 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1061_
timestamp 1698175906
transform 1 0 9856 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1062_
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1063_
timestamp 1698175906
transform 1 0 21840 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1064_
timestamp 1698175906
transform 1 0 23296 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1065_
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1066_
timestamp 1698175906
transform 1 0 26432 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1067_
timestamp 1698175906
transform 1 0 28224 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1068_
timestamp 1698175906
transform 1 0 30128 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1069_
timestamp 1698175906
transform 1 0 25088 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1070_
timestamp 1698175906
transform 1 0 30128 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1071_
timestamp 1698175906
transform 1 0 29456 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1072_
timestamp 1698175906
transform 1 0 30128 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1073_
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1074_
timestamp 1698175906
transform -1 0 12096 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1075_
timestamp 1698175906
transform 1 0 5936 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1076_
timestamp 1698175906
transform -1 0 8736 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1077_
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1078_
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1079_
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1080_
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1081_
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1082_
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1083_
timestamp 1698175906
transform 1 0 5600 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1084_
timestamp 1698175906
transform 1 0 7056 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1085_
timestamp 1698175906
transform 1 0 9520 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1086_
timestamp 1698175906
transform 1 0 8960 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1087_
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1088_
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1089_
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1090_
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1091_
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1092_
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1093_
timestamp 1698175906
transform 1 0 2016 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1094_
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1095_
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1096_
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1097_
timestamp 1698175906
transform 1 0 9632 0 1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1098_
timestamp 1698175906
transform 1 0 15232 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1099_
timestamp 1698175906
transform 1 0 15568 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1100_
timestamp 1698175906
transform 1 0 11872 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1101_
timestamp 1698175906
transform 1 0 18592 0 -1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1102_
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1103_
timestamp 1698175906
transform 1 0 20832 0 -1 28224
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1104_
timestamp 1698175906
transform 1 0 20944 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1105_
timestamp 1698175906
transform 1 0 21392 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1106_
timestamp 1698175906
transform 1 0 5936 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1107_
timestamp 1698175906
transform -1 0 9072 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1108_
timestamp 1698175906
transform -1 0 9072 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1109_
timestamp 1698175906
transform 1 0 4816 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1110_
timestamp 1698175906
transform -1 0 4816 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1111_
timestamp 1698175906
transform -1 0 4816 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0524__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0533__I
timestamp 1698175906
transform -1 0 20496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0537__I
timestamp 1698175906
transform -1 0 26880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0540__I
timestamp 1698175906
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0541__I
timestamp 1698175906
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0545__A1
timestamp 1698175906
transform -1 0 21616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0553__A1
timestamp 1698175906
transform 1 0 15456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0554__A2
timestamp 1698175906
transform -1 0 17472 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0556__I
timestamp 1698175906
transform -1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0557__I
timestamp 1698175906
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0560__I
timestamp 1698175906
transform -1 0 17696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0562__A3
timestamp 1698175906
transform 1 0 28336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0563__I
timestamp 1698175906
transform -1 0 7840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0566__A1
timestamp 1698175906
transform 1 0 29232 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0566__A2
timestamp 1698175906
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0567__A2
timestamp 1698175906
transform -1 0 3808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0569__B
timestamp 1698175906
transform 1 0 18368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0572__A1
timestamp 1698175906
transform 1 0 21952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0573__A3
timestamp 1698175906
transform 1 0 17920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0574__A1
timestamp 1698175906
transform -1 0 20048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0576__A1
timestamp 1698175906
transform 1 0 21504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0578__A1
timestamp 1698175906
transform 1 0 22288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0580__A1
timestamp 1698175906
transform 1 0 21840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0582__A1
timestamp 1698175906
transform 1 0 9184 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0582__B
timestamp 1698175906
transform -1 0 12320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0584__B
timestamp 1698175906
transform -1 0 26768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0584__C
timestamp 1698175906
transform 1 0 32816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0588__I
timestamp 1698175906
transform -1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0590__I
timestamp 1698175906
transform -1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0592__B
timestamp 1698175906
transform -1 0 17920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0599__I
timestamp 1698175906
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0600__A1
timestamp 1698175906
transform -1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0607__A1
timestamp 1698175906
transform 1 0 18144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0611__A1
timestamp 1698175906
transform 1 0 22288 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0611__A2
timestamp 1698175906
transform 1 0 24640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0614__I
timestamp 1698175906
transform -1 0 17696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0617__A1
timestamp 1698175906
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0618__A1
timestamp 1698175906
transform 1 0 29568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0618__A2
timestamp 1698175906
transform 1 0 20272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0619__A1
timestamp 1698175906
transform -1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0622__A1
timestamp 1698175906
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0622__A2
timestamp 1698175906
transform 1 0 29232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0626__A2
timestamp 1698175906
transform -1 0 16464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0630__A1
timestamp 1698175906
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0631__A2
timestamp 1698175906
transform -1 0 19152 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0636__A1
timestamp 1698175906
transform 1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0636__C
timestamp 1698175906
transform 1 0 20496 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0641__A1
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0642__A1
timestamp 1698175906
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0643__I
timestamp 1698175906
transform 1 0 6384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0644__I
timestamp 1698175906
transform 1 0 9632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0646__I
timestamp 1698175906
transform 1 0 5936 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0647__B
timestamp 1698175906
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0650__B
timestamp 1698175906
transform 1 0 4816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0653__A2
timestamp 1698175906
transform -1 0 19152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0654__A3
timestamp 1698175906
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0655__I
timestamp 1698175906
transform -1 0 10528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0657__A2
timestamp 1698175906
transform 1 0 12544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0658__A1
timestamp 1698175906
transform 1 0 11424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0660__A3
timestamp 1698175906
transform 1 0 27664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0661__I
timestamp 1698175906
transform 1 0 14224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0664__I
timestamp 1698175906
transform -1 0 12096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0674__I
timestamp 1698175906
transform 1 0 13104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0677__I
timestamp 1698175906
transform 1 0 14784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0679__A2
timestamp 1698175906
transform 1 0 20272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0682__A2
timestamp 1698175906
transform 1 0 18368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0685__A2
timestamp 1698175906
transform 1 0 20272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0689__A2
timestamp 1698175906
transform 1 0 29120 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0737__I
timestamp 1698175906
transform 1 0 13328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0738__I
timestamp 1698175906
transform 1 0 22176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__A1
timestamp 1698175906
transform 1 0 33152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__A3
timestamp 1698175906
transform -1 0 30128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0763__I
timestamp 1698175906
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__I
timestamp 1698175906
transform 1 0 10864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0784__B
timestamp 1698175906
transform 1 0 23184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0794__A1
timestamp 1698175906
transform 1 0 18592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0816__I0
timestamp 1698175906
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0818__A1
timestamp 1698175906
transform -1 0 12544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0823__I
timestamp 1698175906
transform -1 0 18368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__A1
timestamp 1698175906
transform -1 0 9072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__A2
timestamp 1698175906
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A1
timestamp 1698175906
transform -1 0 7280 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A2
timestamp 1698175906
transform -1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0830__A1
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0832__A1
timestamp 1698175906
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0834__I0
timestamp 1698175906
transform -1 0 17248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0837__B
timestamp 1698175906
transform 1 0 10192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__A1
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0839__I
timestamp 1698175906
transform -1 0 7616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0854__I
timestamp 1698175906
transform 1 0 6720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__I
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__I
timestamp 1698175906
transform 1 0 13664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0895__I
timestamp 1698175906
transform 1 0 14784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__I
timestamp 1698175906
transform 1 0 9632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0920__C
timestamp 1698175906
transform 1 0 8064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__C
timestamp 1698175906
transform -1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__I
timestamp 1698175906
transform -1 0 9968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__I
timestamp 1698175906
transform 1 0 11536 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__C
timestamp 1698175906
transform 1 0 14672 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0968__A1
timestamp 1698175906
transform 1 0 8512 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1000__B
timestamp 1698175906
transform -1 0 17696 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__C
timestamp 1698175906
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__A1
timestamp 1698175906
transform 1 0 8064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__B
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1006__B
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1008__I
timestamp 1698175906
transform -1 0 4592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__I
timestamp 1698175906
transform -1 0 5936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1011__I
timestamp 1698175906
transform 1 0 9408 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__I
timestamp 1698175906
transform -1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__CLK
timestamp 1698175906
transform 1 0 22288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__CLK
timestamp 1698175906
transform 1 0 25312 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__CLK
timestamp 1698175906
transform 1 0 21840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__CLK
timestamp 1698175906
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__CLK
timestamp 1698175906
transform -1 0 25648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1062__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__CLK
timestamp 1698175906
transform -1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__CLK
timestamp 1698175906
transform 1 0 5824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__CLK
timestamp 1698175906
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__CLK
timestamp 1698175906
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__CLK
timestamp 1698175906
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__CLK
timestamp 1698175906
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__CLK
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__CLK
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__CLK
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__CLK
timestamp 1698175906
transform -1 0 12432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__CLK
timestamp 1698175906
transform 1 0 16800 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__CLK
timestamp 1698175906
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1089__CLK
timestamp 1698175906
transform 1 0 16800 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__CLK
timestamp 1698175906
transform 1 0 4816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__CLK
timestamp 1698175906
transform 1 0 5712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__CLK
timestamp 1698175906
transform 1 0 5040 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__CLK
timestamp 1698175906
transform 1 0 4480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__CLK
timestamp 1698175906
transform 1 0 5488 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__CLK
timestamp 1698175906
transform 1 0 5712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__CLK
timestamp 1698175906
transform 1 0 11648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__CLK
timestamp 1698175906
transform -1 0 6832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__CLK
timestamp 1698175906
transform 1 0 9296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__CLK
timestamp 1698175906
transform 1 0 8400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__CLK
timestamp 1698175906
transform 1 0 9632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_i_I
timestamp 1698175906
transform -1 0 22960 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_clk_i_I
timestamp 1698175906
transform -1 0 12544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_clk_i_I
timestamp 1698175906
transform 1 0 19824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_clk_i_I
timestamp 1698175906
transform 1 0 11984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_clk_i_I
timestamp 1698175906
transform 1 0 15792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_clk_i_I
timestamp 1698175906
transform 1 0 22288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_clk_i_I
timestamp 1698175906
transform 1 0 26208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_clk_i_I
timestamp 1698175906
transform 1 0 20944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_clk_i_I
timestamp 1698175906
transform 1 0 13552 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform -1 0 33376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698175906
transform -1 0 9296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698175906
transform -1 0 22848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698175906
transform -1 0 21952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698175906
transform -1 0 22400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698175906
transform -1 0 28448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698175906
transform -1 0 21616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698175906
transform -1 0 27328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698175906
transform -1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698175906
transform -1 0 5152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698175906
transform -1 0 25984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698175906
transform 1 0 25872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698175906
transform 1 0 26992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698175906
transform 1 0 27440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698175906
transform -1 0 21392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698175906
transform -1 0 24416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698175906
transform -1 0 26544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698175906
transform -1 0 22960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698175906
transform -1 0 25200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output33_I
timestamp 1698175906
transform -1 0 20048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1698175906
transform -1 0 5600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1698175906
transform 1 0 19376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1698175906
transform -1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output39_I
timestamp 1698175906
transform -1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23072 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_clk_i
timestamp 1698175906
transform -1 0 12096 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_clk_i
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_clk_i
timestamp 1698175906
transform -1 0 11088 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_clk_i
timestamp 1698175906
transform 1 0 10192 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_clk_i
timestamp 1698175906
transform -1 0 28112 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_clk_i
timestamp 1698175906
transform 1 0 26992 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_clk_i
timestamp 1698175906
transform -1 0 26768 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_clk_i
timestamp 1698175906
transform 1 0 27104 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout58
timestamp 1698175906
transform -1 0 14000 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout59
timestamp 1698175906
transform -1 0 15232 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout60
timestamp 1698175906
transform -1 0 6384 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout61
timestamp 1698175906
transform -1 0 7952 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout62
timestamp 1698175906
transform -1 0 14224 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout63
timestamp 1698175906
transform 1 0 28112 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout64
timestamp 1698175906
transform -1 0 30576 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout65
timestamp 1698175906
transform 1 0 26432 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout66
timestamp 1698175906
transform 1 0 14672 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698175906
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_213
timestamp 1698175906
transform 1 0 25200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_217
timestamp 1698175906
transform 1 0 25648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_227
timestamp 1698175906
transform 1 0 26768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_231
timestamp 1698175906
transform 1 0 27216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_235
timestamp 1698175906
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_246
timestamp 1698175906
transform 1 0 28896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_248
timestamp 1698175906
transform 1 0 29120 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_255
timestamp 1698175906
transform 1 0 29904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_269
timestamp 1698175906
transform 1 0 31472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698175906
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_68
timestamp 1698175906
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_129
timestamp 1698175906
transform 1 0 15792 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_131
timestamp 1698175906
transform 1 0 16016 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_171
timestamp 1698175906
transform 1 0 20496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698175906
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_167
timestamp 1698175906
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_230
timestamp 1698175906
transform 1 0 27104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_232
timestamp 1698175906
transform 1 0 27328 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_255
timestamp 1698175906
transform 1 0 29904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_31
timestamp 1698175906
transform 1 0 4816 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698175906
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_78
timestamp 1698175906
transform 1 0 10080 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698175906
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_154
timestamp 1698175906
transform 1 0 18592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698175906
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_228
timestamp 1698175906
transform 1 0 26880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_235
timestamp 1698175906
transform 1 0 27664 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698175906
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_28
timestamp 1698175906
transform 1 0 4480 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_77
timestamp 1698175906
transform 1 0 9968 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_96
timestamp 1698175906
transform 1 0 12096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_145
timestamp 1698175906
transform 1 0 17584 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_179
timestamp 1698175906
transform 1 0 21392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_209
timestamp 1698175906
transform 1 0 24752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_225
timestamp 1698175906
transform 1 0 26544 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_238
timestamp 1698175906
transform 1 0 28000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_249
timestamp 1698175906
transform 1 0 29232 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_272
timestamp 1698175906
transform 1 0 31808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_4
timestamp 1698175906
transform 1 0 1792 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_45
timestamp 1698175906
transform 1 0 6384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698175906
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_101
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_103
timestamp 1698175906
transform 1 0 12880 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_163
timestamp 1698175906
transform 1 0 19600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_167
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_171 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_175
timestamp 1698175906
transform 1 0 20944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_192
timestamp 1698175906
transform 1 0 22848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_199
timestamp 1698175906
transform 1 0 23632 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_203
timestamp 1698175906
transform 1 0 24080 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_218
timestamp 1698175906
transform 1 0 25760 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_222
timestamp 1698175906
transform 1 0 26208 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_231
timestamp 1698175906
transform 1 0 27216 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_238
timestamp 1698175906
transform 1 0 28000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_253
timestamp 1698175906
transform 1 0 29680 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_277
timestamp 1698175906
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698175906
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_31
timestamp 1698175906
transform 1 0 4816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_96
timestamp 1698175906
transform 1 0 12096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_98
timestamp 1698175906
transform 1 0 12320 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_157
timestamp 1698175906
transform 1 0 18928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_159
timestamp 1698175906
transform 1 0 19152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698175906
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_181
timestamp 1698175906
transform 1 0 21616 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_184
timestamp 1698175906
transform 1 0 21952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_188
timestamp 1698175906
transform 1 0 22400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_212
timestamp 1698175906
transform 1 0 25088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_216
timestamp 1698175906
transform 1 0 25536 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_220
timestamp 1698175906
transform 1 0 25984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_224
timestamp 1698175906
transform 1 0 26432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_228
timestamp 1698175906
transform 1 0 26880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_253
timestamp 1698175906
transform 1 0 29680 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_39
timestamp 1698175906
transform 1 0 5712 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_101
timestamp 1698175906
transform 1 0 12656 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_107
timestamp 1698175906
transform 1 0 13328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698175906
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_155
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_185
timestamp 1698175906
transform 1 0 22064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_189
timestamp 1698175906
transform 1 0 22512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_193
timestamp 1698175906
transform 1 0 22960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698175906
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_255
timestamp 1698175906
transform 1 0 29904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698175906
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_31
timestamp 1698175906
transform 1 0 4816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_98
timestamp 1698175906
transform 1 0 12320 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_102
timestamp 1698175906
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698175906
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_109
timestamp 1698175906
transform 1 0 13552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_163
timestamp 1698175906
transform 1 0 19600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698175906
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_185
timestamp 1698175906
transform 1 0 22064 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_194
timestamp 1698175906
transform 1 0 23072 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_211
timestamp 1698175906
transform 1 0 24976 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698175906
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_255
timestamp 1698175906
transform 1 0 29904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_23
timestamp 1698175906
transform 1 0 3920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_29
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_33
timestamp 1698175906
transform 1 0 5040 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_39
timestamp 1698175906
transform 1 0 5712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_43
timestamp 1698175906
transform 1 0 6160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_63
timestamp 1698175906
transform 1 0 8400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_67
timestamp 1698175906
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698175906
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_76
timestamp 1698175906
transform 1 0 9856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_133
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698175906
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698175906
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_150
timestamp 1698175906
transform 1 0 18144 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_158
timestamp 1698175906
transform 1 0 19040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_180
timestamp 1698175906
transform 1 0 21504 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_228
timestamp 1698175906
transform 1 0 26880 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698175906
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_70
timestamp 1698175906
transform 1 0 9184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_74
timestamp 1698175906
transform 1 0 9632 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_83
timestamp 1698175906
transform 1 0 10640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_87
timestamp 1698175906
transform 1 0 11088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_89
timestamp 1698175906
transform 1 0 11312 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_92
timestamp 1698175906
transform 1 0 11648 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_96
timestamp 1698175906
transform 1 0 12096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_98
timestamp 1698175906
transform 1 0 12320 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_113
timestamp 1698175906
transform 1 0 14000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_117
timestamp 1698175906
transform 1 0 14448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_119
timestamp 1698175906
transform 1 0 14672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_122
timestamp 1698175906
transform 1 0 15008 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_138
timestamp 1698175906
transform 1 0 16800 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_168
timestamp 1698175906
transform 1 0 20160 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_172
timestamp 1698175906
transform 1 0 20608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698175906
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_181
timestamp 1698175906
transform 1 0 21616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_185
timestamp 1698175906
transform 1 0 22064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_282
timestamp 1698175906
transform 1 0 32928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_34
timestamp 1698175906
transform 1 0 5152 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_50
timestamp 1698175906
transform 1 0 6944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_52
timestamp 1698175906
transform 1 0 7168 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_58
timestamp 1698175906
transform 1 0 7840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_62
timestamp 1698175906
transform 1 0 8288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_88
timestamp 1698175906
transform 1 0 11200 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_92
timestamp 1698175906
transform 1 0 11648 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_105
timestamp 1698175906
transform 1 0 13104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_115
timestamp 1698175906
transform 1 0 14224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_123
timestamp 1698175906
transform 1 0 15120 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1698175906
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_158
timestamp 1698175906
transform 1 0 19040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_160
timestamp 1698175906
transform 1 0 19264 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_191
timestamp 1698175906
transform 1 0 22736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_193
timestamp 1698175906
transform 1 0 22960 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_250
timestamp 1698175906
transform 1 0 29344 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_66
timestamp 1698175906
transform 1 0 8736 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_74
timestamp 1698175906
transform 1 0 9632 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_136
timestamp 1698175906
transform 1 0 16576 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_142
timestamp 1698175906
transform 1 0 17248 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_146
timestamp 1698175906
transform 1 0 17696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_155
timestamp 1698175906
transform 1 0 18704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_159
timestamp 1698175906
transform 1 0 19152 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_167
timestamp 1698175906
transform 1 0 20048 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_181
timestamp 1698175906
transform 1 0 21616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_185
timestamp 1698175906
transform 1 0 22064 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_190
timestamp 1698175906
transform 1 0 22624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_192
timestamp 1698175906
transform 1 0 22848 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_233
timestamp 1698175906
transform 1 0 27440 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_251
timestamp 1698175906
transform 1 0 29456 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_283
timestamp 1698175906
transform 1 0 33040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_285
timestamp 1698175906
transform 1 0 33264 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_34
timestamp 1698175906
transform 1 0 5152 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_38
timestamp 1698175906
transform 1 0 5600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_40
timestamp 1698175906
transform 1 0 5824 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_76
timestamp 1698175906
transform 1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_78
timestamp 1698175906
transform 1 0 10080 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_89
timestamp 1698175906
transform 1 0 11312 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_96
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_100
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_108
timestamp 1698175906
transform 1 0 13440 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_112
timestamp 1698175906
transform 1 0 13888 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_172
timestamp 1698175906
transform 1 0 20608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_174
timestamp 1698175906
transform 1 0 20832 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_188
timestamp 1698175906
transform 1 0 22400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_218
timestamp 1698175906
transform 1 0 25760 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_250
timestamp 1698175906
transform 1 0 29344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_31
timestamp 1698175906
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_45
timestamp 1698175906
transform 1 0 6384 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_102
timestamp 1698175906
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698175906
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_164
timestamp 1698175906
transform 1 0 19712 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_181
timestamp 1698175906
transform 1 0 21616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_183
timestamp 1698175906
transform 1 0 21840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_255
timestamp 1698175906
transform 1 0 29904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_31
timestamp 1698175906
transform 1 0 4816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_38
timestamp 1698175906
transform 1 0 5600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_42
timestamp 1698175906
transform 1 0 6048 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_53
timestamp 1698175906
transform 1 0 7280 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_64
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698175906
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_76
timestamp 1698175906
transform 1 0 9856 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_86
timestamp 1698175906
transform 1 0 10976 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_90
timestamp 1698175906
transform 1 0 11424 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_100
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_102
timestamp 1698175906
transform 1 0 12768 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_157
timestamp 1698175906
transform 1 0 18928 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_222
timestamp 1698175906
transform 1 0 26208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_230
timestamp 1698175906
transform 1 0 27104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_232
timestamp 1698175906
transform 1 0 27328 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_246
timestamp 1698175906
transform 1 0 28896 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_250
timestamp 1698175906
transform 1 0 29344 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_18
timestamp 1698175906
transform 1 0 3360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_20
timestamp 1698175906
transform 1 0 3584 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_50
timestamp 1698175906
transform 1 0 6944 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_56
timestamp 1698175906
transform 1 0 7616 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_72
timestamp 1698175906
transform 1 0 9408 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_80
timestamp 1698175906
transform 1 0 10304 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_87
timestamp 1698175906
transform 1 0 11088 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_94
timestamp 1698175906
transform 1 0 11872 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_102
timestamp 1698175906
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698175906
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_123
timestamp 1698175906
transform 1 0 15120 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_131
timestamp 1698175906
transform 1 0 16016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_183
timestamp 1698175906
transform 1 0 21840 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_213
timestamp 1698175906
transform 1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_223
timestamp 1698175906
transform 1 0 26320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_276
timestamp 1698175906
transform 1 0 32256 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_285
timestamp 1698175906
transform 1 0 33264 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_18
timestamp 1698175906
transform 1 0 3360 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_22
timestamp 1698175906
transform 1 0 3808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_37
timestamp 1698175906
transform 1 0 5488 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_54
timestamp 1698175906
transform 1 0 7392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_56
timestamp 1698175906
transform 1 0 7616 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_76
timestamp 1698175906
transform 1 0 9856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_80
timestamp 1698175906
transform 1 0 10304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_93
timestamp 1698175906
transform 1 0 11760 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_99
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_107
timestamp 1698175906
transform 1 0 13328 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_117
timestamp 1698175906
transform 1 0 14448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1698175906
transform 1 0 16240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_194
timestamp 1698175906
transform 1 0 23072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_196
timestamp 1698175906
transform 1 0 23296 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_214
timestamp 1698175906
transform 1 0 25312 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_239
timestamp 1698175906
transform 1 0 28112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_243
timestamp 1698175906
transform 1 0 28560 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_252
timestamp 1698175906
transform 1 0 29568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_254
timestamp 1698175906
transform 1 0 29792 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_31
timestamp 1698175906
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_43
timestamp 1698175906
transform 1 0 6160 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_58
timestamp 1698175906
transform 1 0 7840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_66
timestamp 1698175906
transform 1 0 8736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698175906
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_136
timestamp 1698175906
transform 1 0 16576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_140
timestamp 1698175906
transform 1 0 17024 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_170
timestamp 1698175906
transform 1 0 20384 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_200
timestamp 1698175906
transform 1 0 23744 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_241
timestamp 1698175906
transform 1 0 28336 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_10
timestamp 1698175906
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_12
timestamp 1698175906
transform 1 0 2688 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_36
timestamp 1698175906
transform 1 0 5376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_46
timestamp 1698175906
transform 1 0 6496 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_50
timestamp 1698175906
transform 1 0 6944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_52
timestamp 1698175906
transform 1 0 7168 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_59
timestamp 1698175906
transform 1 0 7952 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_80
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_82
timestamp 1698175906
transform 1 0 10528 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_96
timestamp 1698175906
transform 1 0 12096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_100
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_102
timestamp 1698175906
transform 1 0 12768 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_134
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_169
timestamp 1698175906
transform 1 0 20272 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_173
timestamp 1698175906
transform 1 0 20720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_187
timestamp 1698175906
transform 1 0 22288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_189
timestamp 1698175906
transform 1 0 22512 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_31
timestamp 1698175906
transform 1 0 4816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_42
timestamp 1698175906
transform 1 0 6048 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_63
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_65
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_71
timestamp 1698175906
transform 1 0 9296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_75
timestamp 1698175906
transform 1 0 9744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_79
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_93
timestamp 1698175906
transform 1 0 11760 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_148
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_152
timestamp 1698175906
transform 1 0 18368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_156
timestamp 1698175906
transform 1 0 18816 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_159
timestamp 1698175906
transform 1 0 19152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_163
timestamp 1698175906
transform 1 0 19600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_167
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_181
timestamp 1698175906
transform 1 0 21616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_185
timestamp 1698175906
transform 1 0 22064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_189
timestamp 1698175906
transform 1 0 22512 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_217
timestamp 1698175906
transform 1 0 25648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_229
timestamp 1698175906
transform 1 0 26992 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_279
timestamp 1698175906
transform 1 0 32592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_283
timestamp 1698175906
transform 1 0 33040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_285
timestamp 1698175906
transform 1 0 33264 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_18
timestamp 1698175906
transform 1 0 3360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_31
timestamp 1698175906
transform 1 0 4816 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698175906
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698175906
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_102
timestamp 1698175906
transform 1 0 12768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_106
timestamp 1698175906
transform 1 0 13216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_121
timestamp 1698175906
transform 1 0 14896 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_127
timestamp 1698175906
transform 1 0 15568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_129
timestamp 1698175906
transform 1 0 15792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_135
timestamp 1698175906
transform 1 0 16464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_137
timestamp 1698175906
transform 1 0 16688 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_171
timestamp 1698175906
transform 1 0 20496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_177
timestamp 1698175906
transform 1 0 21168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_179
timestamp 1698175906
transform 1 0 21392 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_182
timestamp 1698175906
transform 1 0 21728 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698175906
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_262
timestamp 1698175906
transform 1 0 30688 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_18
timestamp 1698175906
transform 1 0 3360 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_22
timestamp 1698175906
transform 1 0 3808 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_31
timestamp 1698175906
transform 1 0 4816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_42
timestamp 1698175906
transform 1 0 6048 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_80
timestamp 1698175906
transform 1 0 10304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_82
timestamp 1698175906
transform 1 0 10528 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_88
timestamp 1698175906
transform 1 0 11200 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_90
timestamp 1698175906
transform 1 0 11424 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_93
timestamp 1698175906
transform 1 0 11760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_97
timestamp 1698175906
transform 1 0 12208 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_136
timestamp 1698175906
transform 1 0 16576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_140
timestamp 1698175906
transform 1 0 17024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_152
timestamp 1698175906
transform 1 0 18368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_154
timestamp 1698175906
transform 1 0 18592 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_170
timestamp 1698175906
transform 1 0 20384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_172
timestamp 1698175906
transform 1 0 20608 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_206
timestamp 1698175906
transform 1 0 24416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_39
timestamp 1698175906
transform 1 0 5712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_51
timestamp 1698175906
transform 1 0 7056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_77
timestamp 1698175906
transform 1 0 9968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_79
timestamp 1698175906
transform 1 0 10192 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_82
timestamp 1698175906
transform 1 0 10528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_84
timestamp 1698175906
transform 1 0 10752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_91
timestamp 1698175906
transform 1 0 11536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_93
timestamp 1698175906
transform 1 0 11760 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_107
timestamp 1698175906
transform 1 0 13328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_109
timestamp 1698175906
transform 1 0 13552 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_118
timestamp 1698175906
transform 1 0 14560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_122
timestamp 1698175906
transform 1 0 15008 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_128
timestamp 1698175906
transform 1 0 15680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_132
timestamp 1698175906
transform 1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_146
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698175906
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_185
timestamp 1698175906
transform 1 0 22064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_256
timestamp 1698175906
transform 1 0 30016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_31
timestamp 1698175906
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_98
timestamp 1698175906
transform 1 0 12320 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_127
timestamp 1698175906
transform 1 0 15568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_145
timestamp 1698175906
transform 1 0 17584 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_149
timestamp 1698175906
transform 1 0 18032 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_152
timestamp 1698175906
transform 1 0 18368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_163
timestamp 1698175906
transform 1 0 19600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_167
timestamp 1698175906
transform 1 0 20048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_18
timestamp 1698175906
transform 1 0 3360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_26
timestamp 1698175906
transform 1 0 4256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_30
timestamp 1698175906
transform 1 0 4704 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_45
timestamp 1698175906
transform 1 0 6384 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_59
timestamp 1698175906
transform 1 0 7952 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_63
timestamp 1698175906
transform 1 0 8400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_78
timestamp 1698175906
transform 1 0 10080 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698175906
transform 1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698175906
transform 1 0 17920 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_175
timestamp 1698175906
transform 1 0 20944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_177
timestamp 1698175906
transform 1 0 21168 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_198
timestamp 1698175906
transform 1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698175906
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_33
timestamp 1698175906
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_68
timestamp 1698175906
transform 1 0 8960 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_72
timestamp 1698175906
transform 1 0 9408 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_74
timestamp 1698175906
transform 1 0 9632 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_117
timestamp 1698175906
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_141
timestamp 1698175906
transform 1 0 17136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_143
timestamp 1698175906
transform 1 0 17360 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_183
timestamp 1698175906
transform 1 0 21840 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_236
timestamp 1698175906
transform 1 0 27776 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_31
timestamp 1698175906
transform 1 0 4816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_33
timestamp 1698175906
transform 1 0 5040 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_42
timestamp 1698175906
transform 1 0 6048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698175906
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_87
timestamp 1698175906
transform 1 0 11088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_91
timestamp 1698175906
transform 1 0 11536 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_94
timestamp 1698175906
transform 1 0 11872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_114
timestamp 1698175906
transform 1 0 14112 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_147
timestamp 1698175906
transform 1 0 17808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_149
timestamp 1698175906
transform 1 0 18032 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_218
timestamp 1698175906
transform 1 0 25760 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_271
timestamp 1698175906
transform 1 0 31696 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_18
timestamp 1698175906
transform 1 0 3360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_20
timestamp 1698175906
transform 1 0 3584 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_58
timestamp 1698175906
transform 1 0 7840 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_66
timestamp 1698175906
transform 1 0 8736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_68
timestamp 1698175906
transform 1 0 8960 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_93
timestamp 1698175906
transform 1 0 11760 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_151
timestamp 1698175906
transform 1 0 18256 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_168
timestamp 1698175906
transform 1 0 20160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_18
timestamp 1698175906
transform 1 0 3360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_26
timestamp 1698175906
transform 1 0 4256 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_39
timestamp 1698175906
transform 1 0 5712 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_59
timestamp 1698175906
transform 1 0 7952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698175906
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_91
timestamp 1698175906
transform 1 0 11536 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_176
timestamp 1698175906
transform 1 0 21056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_178
timestamp 1698175906
transform 1 0 21280 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_239
timestamp 1698175906
transform 1 0 28112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_10
timestamp 1698175906
transform 1 0 2464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_20
timestamp 1698175906
transform 1 0 3584 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_67
timestamp 1698175906
transform 1 0 8848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_69
timestamp 1698175906
transform 1 0 9072 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_90
timestamp 1698175906
transform 1 0 11424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_209
timestamp 1698175906
transform 1 0 24752 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_211
timestamp 1698175906
transform 1 0 24976 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_31
timestamp 1698175906
transform 1 0 4816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_35
timestamp 1698175906
transform 1 0 5264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_39
timestamp 1698175906
transform 1 0 5712 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_54
timestamp 1698175906
transform 1 0 7392 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_58
timestamp 1698175906
transform 1 0 7840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_62
timestamp 1698175906
transform 1 0 8288 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_31
timestamp 1698175906
transform 1 0 4816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_51
timestamp 1698175906
transform 1 0 7056 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_53
timestamp 1698175906
transform 1 0 7280 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_60
timestamp 1698175906
transform 1 0 8064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_62
timestamp 1698175906
transform 1 0 8288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_65
timestamp 1698175906
transform 1 0 8624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_69
timestamp 1698175906
transform 1 0 9072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_18
timestamp 1698175906
transform 1 0 3360 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_26
timestamp 1698175906
transform 1 0 4256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_30
timestamp 1698175906
transform 1 0 4704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_34
timestamp 1698175906
transform 1 0 5152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_44
timestamp 1698175906
transform 1 0 6272 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_46
timestamp 1698175906
transform 1 0 6496 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_49
timestamp 1698175906
transform 1 0 6832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_82
timestamp 1698175906
transform 1 0 10528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_123
timestamp 1698175906
transform 1 0 15120 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_125
timestamp 1698175906
transform 1 0 15344 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_137
timestamp 1698175906
transform 1 0 16688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698175906
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698175906
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_125
timestamp 1698175906
transform 1 0 15344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_156
timestamp 1698175906
transform 1 0 18816 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_243
timestamp 1698175906
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_11
timestamp 1698175906
transform 1 0 2576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_17
timestamp 1698175906
transform 1 0 3248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_19
timestamp 1698175906
transform 1 0 3472 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_36
timestamp 1698175906
transform 1 0 5376 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_101
timestamp 1698175906
transform 1 0 12656 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_104
timestamp 1698175906
transform 1 0 12992 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_269
timestamp 1698175906
transform 1 0 31472 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_271
timestamp 1698175906
transform 1 0 31696 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_285
timestamp 1698175906
transform 1 0 33264 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698175906
transform 1 0 30016 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698175906
transform -1 0 24192 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698175906
transform -1 0 30016 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698175906
transform -1 0 32704 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698175906
transform -1 0 33376 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698175906
transform 1 0 27440 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698175906
transform -1 0 32928 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698175906
transform 1 0 25424 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698175906
transform -1 0 19824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698175906
transform -1 0 33376 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698175906
transform -1 0 24192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698175906
transform -1 0 25200 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698175906
transform -1 0 26768 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698175906
transform -1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698175906
transform -1 0 29904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698175906
transform 1 0 30800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698175906
transform 1 0 30128 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11088 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 12880 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 14000 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 13664 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 17360 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 17472 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698175906
transform 1 0 20608 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output29
timestamp 1698175906
transform -1 0 24752 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output30
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output31
timestamp 1698175906
transform 1 0 25760 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output32
timestamp 1698175906
transform 1 0 25200 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output33
timestamp 1698175906
transform 1 0 29680 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output34
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output35
timestamp 1698175906
transform -1 0 32592 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output36
timestamp 1698175906
transform 1 0 29680 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output37
timestamp 1698175906
transform -1 0 32704 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output38
timestamp 1698175906
transform 1 0 29792 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output39
timestamp 1698175906
transform 1 0 30464 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output40
timestamp 1698175906
transform 1 0 28784 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output41
timestamp 1698175906
transform 1 0 6048 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output42
timestamp 1698175906
transform 1 0 10192 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output43
timestamp 1698175906
transform -1 0 4480 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output44
timestamp 1698175906
transform -1 0 5264 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output45
timestamp 1698175906
transform 1 0 2240 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output46
timestamp 1698175906
transform 1 0 5712 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output47
timestamp 1698175906
transform -1 0 8848 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output48
timestamp 1698175906
transform 1 0 6048 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49
timestamp 1698175906
transform -1 0 28784 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698175906
transform -1 0 12544 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698175906
transform 1 0 11200 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698175906
transform 1 0 13552 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698175906
transform 1 0 14112 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698175906
transform 1 0 13664 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698175906
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output57
timestamp 1698175906
transform 1 0 21392 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 33600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_37
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 33600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_38
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 33600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_39
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 33600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_40
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 33600 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_41
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 33600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_42
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 33600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_43
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 33600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_44
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 33600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_45
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 33600 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_46
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 33600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_47
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 33600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_48
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 33600 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_49
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 33600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_50
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 33600 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_51
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 33600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_52
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 33600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_53
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 33600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_54
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 33600 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_55
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 33600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_56
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 33600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_57
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 33600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_58
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 33600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_59
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 33600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_60
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 33600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_61
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 33600 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_62
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 33600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_63
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 33600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_64
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 33600 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_65
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 33600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_66
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 33600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_67
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 33600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_68
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 33600 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_69
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 33600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_70
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 33600 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_71
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 33600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_72 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_73
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_74
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_75
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_76
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_77
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_78
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_79
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_80
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_81
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_82
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_83
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_84
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_85
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_86
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_87
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_88
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_89
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_90
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_91
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_92
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_93
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_94
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_95
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_96
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_97
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_98
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_99
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_100
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_101
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_102
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_103
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_104
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_105
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_106
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_107
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_108
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_109
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_110
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_111
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_112
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_113
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_114
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_115
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_116
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_117
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_118
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_119
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_120
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_121
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_122
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_123
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_124
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_125
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_127
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_128
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_129
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_131
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_132
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_133
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_134
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_135
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_136
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_137
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_138
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_139
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_140
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_141
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_142
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_143
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_144
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_145
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_146
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_147
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_148
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_149
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_150
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_151
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_152
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_153
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_154
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_155
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_156
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_157
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_158
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_159
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_160
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_161
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_162
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_163
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_164
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_165
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_166
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_167
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_168
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_169
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_170
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_171
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_172
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_173
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_174
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_175
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_176
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_177
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_178
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_179
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_180
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_181
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_182
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_183
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_184
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_185
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_186
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_187
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_188
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_189
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_190
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_191
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_192
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_193
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_194
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_195
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_196
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_197
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_198
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_199
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_200
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_201
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_202
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_203
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_204
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_205
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_206
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_207
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_208
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_209
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_210
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_211
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_212
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_213
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_214
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_215
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_216
timestamp 1698175906
transform 1 0 5152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_217
timestamp 1698175906
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_218
timestamp 1698175906
transform 1 0 12768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_219
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_220
timestamp 1698175906
transform 1 0 20384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_221
timestamp 1698175906
transform 1 0 24192 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_222
timestamp 1698175906
transform 1 0 28000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_223
timestamp 1698175906
transform 1 0 31808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_67 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 2576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_68
timestamp 1698175906
transform -1 0 2128 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_69
timestamp 1698175906
transform -1 0 3248 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_70
timestamp 1698175906
transform -1 0 4256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_71
timestamp 1698175906
transform 1 0 4256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_72
timestamp 1698175906
transform 1 0 4704 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_73
timestamp 1698175906
transform 1 0 5600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_mc14500_74
timestamp 1698175906
transform -1 0 9184 0 1 29792
box -86 -86 534 870
<< labels >>
flabel metal3 s 34200 28000 35000 28112 0 FreeSans 448 0 0 0 SDI
port 0 nsew signal input
flabel metal3 s 34200 1120 35000 1232 0 FreeSans 448 0 0 0 clk_i
port 1 nsew signal input
flabel metal3 s 34200 33376 35000 33488 0 FreeSans 448 0 0 0 custom_setting
port 2 nsew signal input
flabel metal3 s 34200 6496 35000 6608 0 FreeSans 448 0 0 0 io_in[0]
port 3 nsew signal input
flabel metal3 s 34200 9184 35000 9296 0 FreeSans 448 0 0 0 io_in[1]
port 4 nsew signal input
flabel metal3 s 34200 11872 35000 11984 0 FreeSans 448 0 0 0 io_in[2]
port 5 nsew signal input
flabel metal3 s 34200 14560 35000 14672 0 FreeSans 448 0 0 0 io_in[3]
port 6 nsew signal input
flabel metal3 s 34200 17248 35000 17360 0 FreeSans 448 0 0 0 io_in[4]
port 7 nsew signal input
flabel metal3 s 34200 19936 35000 20048 0 FreeSans 448 0 0 0 io_in[5]
port 8 nsew signal input
flabel metal3 s 34200 22624 35000 22736 0 FreeSans 448 0 0 0 io_in[6]
port 9 nsew signal input
flabel metal3 s 34200 25312 35000 25424 0 FreeSans 448 0 0 0 io_in[7]
port 10 nsew signal input
flabel metal2 s 448 34200 560 35000 0 FreeSans 448 90 0 0 io_out[0]
port 11 nsew signal tristate
flabel metal2 s 11648 34200 11760 35000 0 FreeSans 448 90 0 0 io_out[10]
port 12 nsew signal tristate
flabel metal2 s 12768 34200 12880 35000 0 FreeSans 448 90 0 0 io_out[11]
port 13 nsew signal tristate
flabel metal2 s 13888 34200 14000 35000 0 FreeSans 448 90 0 0 io_out[12]
port 14 nsew signal tristate
flabel metal2 s 15008 34200 15120 35000 0 FreeSans 448 90 0 0 io_out[13]
port 15 nsew signal tristate
flabel metal2 s 16128 34200 16240 35000 0 FreeSans 448 90 0 0 io_out[14]
port 16 nsew signal tristate
flabel metal2 s 17248 34200 17360 35000 0 FreeSans 448 90 0 0 io_out[15]
port 17 nsew signal tristate
flabel metal2 s 18368 34200 18480 35000 0 FreeSans 448 90 0 0 io_out[16]
port 18 nsew signal tristate
flabel metal2 s 19488 34200 19600 35000 0 FreeSans 448 90 0 0 io_out[17]
port 19 nsew signal tristate
flabel metal2 s 20608 34200 20720 35000 0 FreeSans 448 90 0 0 io_out[18]
port 20 nsew signal tristate
flabel metal2 s 21728 34200 21840 35000 0 FreeSans 448 90 0 0 io_out[19]
port 21 nsew signal tristate
flabel metal2 s 1568 34200 1680 35000 0 FreeSans 448 90 0 0 io_out[1]
port 22 nsew signal tristate
flabel metal2 s 22848 34200 22960 35000 0 FreeSans 448 90 0 0 io_out[20]
port 23 nsew signal tristate
flabel metal2 s 23968 34200 24080 35000 0 FreeSans 448 90 0 0 io_out[21]
port 24 nsew signal tristate
flabel metal2 s 25088 34200 25200 35000 0 FreeSans 448 90 0 0 io_out[22]
port 25 nsew signal tristate
flabel metal2 s 26208 34200 26320 35000 0 FreeSans 448 90 0 0 io_out[23]
port 26 nsew signal tristate
flabel metal2 s 27328 34200 27440 35000 0 FreeSans 448 90 0 0 io_out[24]
port 27 nsew signal tristate
flabel metal2 s 28448 34200 28560 35000 0 FreeSans 448 90 0 0 io_out[25]
port 28 nsew signal tristate
flabel metal2 s 29568 34200 29680 35000 0 FreeSans 448 90 0 0 io_out[26]
port 29 nsew signal tristate
flabel metal2 s 30688 34200 30800 35000 0 FreeSans 448 90 0 0 io_out[27]
port 30 nsew signal tristate
flabel metal2 s 31808 34200 31920 35000 0 FreeSans 448 90 0 0 io_out[28]
port 31 nsew signal tristate
flabel metal2 s 32928 34200 33040 35000 0 FreeSans 448 90 0 0 io_out[29]
port 32 nsew signal tristate
flabel metal2 s 2688 34200 2800 35000 0 FreeSans 448 90 0 0 io_out[2]
port 33 nsew signal tristate
flabel metal2 s 34048 34200 34160 35000 0 FreeSans 448 90 0 0 io_out[30]
port 34 nsew signal tristate
flabel metal2 s 3808 34200 3920 35000 0 FreeSans 448 90 0 0 io_out[3]
port 35 nsew signal tristate
flabel metal2 s 4928 34200 5040 35000 0 FreeSans 448 90 0 0 io_out[4]
port 36 nsew signal tristate
flabel metal2 s 6048 34200 6160 35000 0 FreeSans 448 90 0 0 io_out[5]
port 37 nsew signal tristate
flabel metal2 s 7168 34200 7280 35000 0 FreeSans 448 90 0 0 io_out[6]
port 38 nsew signal tristate
flabel metal2 s 8288 34200 8400 35000 0 FreeSans 448 90 0 0 io_out[7]
port 39 nsew signal tristate
flabel metal2 s 9408 34200 9520 35000 0 FreeSans 448 90 0 0 io_out[8]
port 40 nsew signal tristate
flabel metal2 s 10528 34200 10640 35000 0 FreeSans 448 90 0 0 io_out[9]
port 41 nsew signal tristate
flabel metal3 s 34200 3808 35000 3920 0 FreeSans 448 0 0 0 rst_n
port 42 nsew signal input
flabel metal2 s 896 0 1008 800 0 FreeSans 448 90 0 0 sram_addr[0]
port 43 nsew signal tristate
flabel metal2 s 2464 0 2576 800 0 FreeSans 448 90 0 0 sram_addr[1]
port 44 nsew signal tristate
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 sram_addr[2]
port 45 nsew signal tristate
flabel metal2 s 5600 0 5712 800 0 FreeSans 448 90 0 0 sram_addr[3]
port 46 nsew signal tristate
flabel metal2 s 7168 0 7280 800 0 FreeSans 448 90 0 0 sram_addr[4]
port 47 nsew signal tristate
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 sram_addr[5]
port 48 nsew signal tristate
flabel metal3 s 34200 30688 35000 30800 0 FreeSans 448 0 0 0 sram_gwe
port 49 nsew signal tristate
flabel metal2 s 10304 0 10416 800 0 FreeSans 448 90 0 0 sram_in[0]
port 50 nsew signal tristate
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 sram_in[1]
port 51 nsew signal tristate
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 sram_in[2]
port 52 nsew signal tristate
flabel metal2 s 15008 0 15120 800 0 FreeSans 448 90 0 0 sram_in[3]
port 53 nsew signal tristate
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 sram_in[4]
port 54 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 sram_in[5]
port 55 nsew signal tristate
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 sram_in[6]
port 56 nsew signal tristate
flabel metal2 s 21280 0 21392 800 0 FreeSans 448 90 0 0 sram_in[7]
port 57 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 sram_out[0]
port 58 nsew signal input
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 sram_out[1]
port 59 nsew signal input
flabel metal2 s 25984 0 26096 800 0 FreeSans 448 90 0 0 sram_out[2]
port 60 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 sram_out[3]
port 61 nsew signal input
flabel metal2 s 29120 0 29232 800 0 FreeSans 448 90 0 0 sram_out[4]
port 62 nsew signal input
flabel metal2 s 30688 0 30800 800 0 FreeSans 448 90 0 0 sram_out[5]
port 63 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 sram_out[6]
port 64 nsew signal input
flabel metal2 s 33824 0 33936 800 0 FreeSans 448 90 0 0 sram_out[7]
port 65 nsew signal input
flabel metal4 s 5216 3076 5536 31420 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 13280 3076 13600 31420 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 21344 3076 21664 31420 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 29408 3076 29728 31420 0 FreeSans 1280 90 0 0 vdd
port 66 nsew power bidirectional
flabel metal4 s 9248 3076 9568 31420 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
flabel metal4 s 17312 3076 17632 31420 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
flabel metal4 s 25376 3076 25696 31420 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
flabel metal4 s 33440 3076 33760 31420 0 FreeSans 1280 90 0 0 vss
port 67 nsew ground bidirectional
rlabel metal1 17472 30576 17472 30576 0 vdd
rlabel via1 17552 31360 17552 31360 0 vss
rlabel metal2 30296 20048 30296 20048 0 SDI
rlabel metal2 14504 14896 14504 14896 0 _0000_
rlabel metal2 17864 12712 17864 12712 0 _0001_
rlabel metal2 20216 12824 20216 12824 0 _0002_
rlabel metal2 23016 19656 23016 19656 0 _0003_
rlabel metal3 23296 21784 23296 21784 0 _0004_
rlabel metal3 25760 23800 25760 23800 0 _0005_
rlabel metal2 26040 27944 26040 27944 0 _0006_
rlabel metal2 31080 25816 31080 25816 0 _0007_
rlabel metal2 31136 27160 31136 27160 0 _0008_
rlabel metal2 28504 23296 28504 23296 0 _0009_
rlabel metal2 27440 29288 27440 29288 0 _0010_
rlabel metal2 3080 7896 3080 7896 0 _0011_
rlabel metal2 3416 9352 3416 9352 0 _0012_
rlabel metal2 10024 10192 10024 10192 0 _0013_
rlabel metal2 10920 7056 10920 7056 0 _0014_
rlabel metal3 10192 5208 10192 5208 0 _0015_
rlabel metal2 11704 4368 11704 4368 0 _0016_
rlabel metal2 14840 4480 14840 4480 0 _0017_
rlabel metal2 14392 6216 14392 6216 0 _0018_
rlabel metal2 16632 4760 16632 4760 0 _0019_
rlabel metal2 18200 5208 18200 5208 0 _0020_
rlabel metal3 13496 9912 13496 9912 0 _0021_
rlabel metal2 14392 9128 14392 9128 0 _0022_
rlabel metal2 17304 9968 17304 9968 0 _0023_
rlabel metal2 19768 9688 19768 9688 0 _0024_
rlabel metal2 23464 10192 23464 10192 0 _0025_
rlabel metal2 26264 11424 26264 11424 0 _0026_
rlabel metal2 26712 9352 26712 9352 0 _0027_
rlabel metal2 28392 10584 28392 10584 0 _0028_
rlabel metal3 20216 6440 20216 6440 0 _0029_
rlabel metal3 21224 5992 21224 5992 0 _0030_
rlabel metal2 21672 4760 21672 4760 0 _0031_
rlabel metal2 25984 4424 25984 4424 0 _0032_
rlabel metal2 29288 4648 29288 4648 0 _0033_
rlabel metal2 31864 4816 31864 4816 0 _0034_
rlabel metal2 32088 7784 32088 7784 0 _0035_
rlabel metal2 32312 9464 32312 9464 0 _0036_
rlabel metal2 23464 28952 23464 28952 0 _0037_
rlabel metal2 18760 29456 18760 29456 0 _0038_
rlabel metal2 19320 21168 19320 21168 0 _0039_
rlabel metal2 14224 13944 14224 13944 0 _0040_
rlabel metal2 10808 13272 10808 13272 0 _0041_
rlabel metal2 18144 20104 18144 20104 0 _0042_
rlabel metal3 22904 29456 22904 29456 0 _0043_
rlabel metal2 31080 29512 31080 29512 0 _0044_
rlabel metal2 14616 12600 14616 12600 0 _0045_
rlabel metal2 10808 15512 10808 15512 0 _0046_
rlabel metal2 6888 14000 6888 14000 0 _0047_
rlabel metal3 7280 12824 7280 12824 0 _0048_
rlabel metal2 2520 14896 2520 14896 0 _0049_
rlabel metal2 2520 15624 2520 15624 0 _0050_
rlabel metal2 4536 17304 4536 17304 0 _0051_
rlabel metal2 2520 18704 2520 18704 0 _0052_
rlabel metal2 4200 21168 4200 21168 0 _0053_
rlabel metal2 2520 22008 2520 22008 0 _0054_
rlabel metal2 6552 20328 6552 20328 0 _0055_
rlabel metal2 8064 20888 8064 20888 0 _0056_
rlabel metal2 10528 19320 10528 19320 0 _0057_
rlabel metal2 9912 18032 9912 18032 0 _0058_
rlabel metal2 14280 17864 14280 17864 0 _0059_
rlabel metal2 14952 18872 14952 18872 0 _0060_
rlabel metal2 14392 20440 14392 20440 0 _0061_
rlabel metal2 2520 23576 2520 23576 0 _0062_
rlabel metal2 7672 29400 7672 29400 0 _0063_
rlabel metal2 2856 27496 2856 27496 0 _0064_
rlabel metal2 3976 29848 3976 29848 0 _0065_
rlabel metal2 3304 27888 3304 27888 0 _0066_
rlabel metal2 2520 25032 2520 25032 0 _0067_
rlabel metal2 10136 30240 10136 30240 0 _0068_
rlabel metal2 9632 28840 9632 28840 0 _0069_
rlabel metal2 16240 26488 16240 26488 0 _0070_
rlabel metal2 16520 30296 16520 30296 0 _0071_
rlabel metal2 12768 29512 12768 29512 0 _0072_
rlabel metal3 18704 29288 18704 29288 0 _0073_
rlabel metal3 21056 26488 21056 26488 0 _0074_
rlabel metal3 20384 27720 20384 27720 0 _0075_
rlabel metal3 21000 23688 21000 23688 0 _0076_
rlabel metal2 18088 25648 18088 25648 0 _0077_
rlabel metal2 6888 11032 6888 11032 0 _0078_
rlabel metal2 8120 9240 8120 9240 0 _0079_
rlabel metal2 8120 6104 8120 6104 0 _0080_
rlabel metal2 5768 5264 5768 5264 0 _0081_
rlabel metal2 3864 5040 3864 5040 0 _0082_
rlabel metal2 3864 6216 3864 6216 0 _0083_
rlabel metal2 23800 13104 23800 13104 0 _0084_
rlabel metal3 30184 14280 30184 14280 0 _0085_
rlabel metal2 23464 14168 23464 14168 0 _0086_
rlabel metal2 24360 13440 24360 13440 0 _0087_
rlabel metal3 22960 15288 22960 15288 0 _0088_
rlabel metal2 26040 15456 26040 15456 0 _0089_
rlabel metal3 25872 15400 25872 15400 0 _0090_
rlabel metal2 24136 15568 24136 15568 0 _0091_
rlabel metal3 25200 15288 25200 15288 0 _0092_
rlabel metal3 24864 13944 24864 13944 0 _0093_
rlabel metal2 24696 15680 24696 15680 0 _0094_
rlabel metal2 20664 17248 20664 17248 0 _0095_
rlabel metal2 20776 17920 20776 17920 0 _0096_
rlabel metal2 23128 13776 23128 13776 0 _0097_
rlabel metal2 22904 14224 22904 14224 0 _0098_
rlabel metal2 18984 13496 18984 13496 0 _0099_
rlabel metal2 20664 15008 20664 15008 0 _0100_
rlabel metal2 23912 15792 23912 15792 0 _0101_
rlabel metal3 20776 18424 20776 18424 0 _0102_
rlabel metal3 23576 18424 23576 18424 0 _0103_
rlabel metal2 23912 22848 23912 22848 0 _0104_
rlabel metal2 26376 29288 26376 29288 0 _0105_
rlabel metal3 33264 24696 33264 24696 0 _0106_
rlabel metal2 22680 23912 22680 23912 0 _0107_
rlabel metal2 25480 22736 25480 22736 0 _0108_
rlabel via2 22232 26152 22232 26152 0 _0109_
rlabel metal2 25256 21504 25256 21504 0 _0110_
rlabel metal3 24920 21672 24920 21672 0 _0111_
rlabel metal2 29288 18928 29288 18928 0 _0112_
rlabel metal3 28056 23912 28056 23912 0 _0113_
rlabel metal2 24472 15624 24472 15624 0 _0114_
rlabel metal2 23240 18200 23240 18200 0 _0115_
rlabel metal2 23912 17248 23912 17248 0 _0116_
rlabel metal2 23072 12936 23072 12936 0 _0117_
rlabel metal2 24136 16632 24136 16632 0 _0118_
rlabel metal2 24640 17080 24640 17080 0 _0119_
rlabel metal2 26488 18592 26488 18592 0 _0120_
rlabel metal3 24584 23688 24584 23688 0 _0121_
rlabel metal2 22456 23912 22456 23912 0 _0122_
rlabel metal2 26488 28224 26488 28224 0 _0123_
rlabel metal2 29624 26628 29624 26628 0 _0124_
rlabel metal2 21896 19376 21896 19376 0 _0125_
rlabel metal2 26264 19208 26264 19208 0 _0126_
rlabel metal3 23576 19152 23576 19152 0 _0127_
rlabel metal2 25032 19152 25032 19152 0 _0128_
rlabel metal3 26040 22232 26040 22232 0 _0129_
rlabel metal2 28448 20104 28448 20104 0 _0130_
rlabel metal2 12152 15176 12152 15176 0 _0131_
rlabel metal2 25592 22512 25592 22512 0 _0132_
rlabel metal2 25368 29400 25368 29400 0 _0133_
rlabel metal2 26264 28616 26264 28616 0 _0134_
rlabel metal2 21896 29736 21896 29736 0 _0135_
rlabel metal2 23016 23016 23016 23016 0 _0136_
rlabel metal2 27608 22680 27608 22680 0 _0137_
rlabel metal2 21560 19824 21560 19824 0 _0138_
rlabel metal2 22624 19768 22624 19768 0 _0139_
rlabel metal2 23912 21952 23912 21952 0 _0140_
rlabel metal2 23240 21840 23240 21840 0 _0141_
rlabel metal3 23744 19432 23744 19432 0 _0142_
rlabel via2 23912 20104 23912 20104 0 _0143_
rlabel metal2 23744 19432 23744 19432 0 _0144_
rlabel metal3 23016 19264 23016 19264 0 _0145_
rlabel metal2 24696 25144 24696 25144 0 _0146_
rlabel metal3 28560 26936 28560 26936 0 _0147_
rlabel metal2 27272 21280 27272 21280 0 _0148_
rlabel metal2 21224 12936 21224 12936 0 _0149_
rlabel metal2 19992 15624 19992 15624 0 _0150_
rlabel metal3 20272 15512 20272 15512 0 _0151_
rlabel metal2 19096 15680 19096 15680 0 _0152_
rlabel metal2 11592 11200 11592 11200 0 _0153_
rlabel metal2 11928 25816 11928 25816 0 _0154_
rlabel metal3 20664 15288 20664 15288 0 _0155_
rlabel metal3 18480 16072 18480 16072 0 _0156_
rlabel metal3 19096 13720 19096 13720 0 _0157_
rlabel metal3 25816 19880 25816 19880 0 _0158_
rlabel metal2 27720 21112 27720 21112 0 _0159_
rlabel metal2 32200 18592 32200 18592 0 _0160_
rlabel metal2 28000 20776 28000 20776 0 _0161_
rlabel metal2 28168 21056 28168 21056 0 _0162_
rlabel metal3 26488 13104 26488 13104 0 _0163_
rlabel metal2 27272 18088 27272 18088 0 _0164_
rlabel metal2 28448 20776 28448 20776 0 _0165_
rlabel metal2 30632 18424 30632 18424 0 _0166_
rlabel metal2 32312 21448 32312 21448 0 _0167_
rlabel metal2 22344 15400 22344 15400 0 _0168_
rlabel metal2 31752 19992 31752 19992 0 _0169_
rlabel metal2 32536 21448 32536 21448 0 _0170_
rlabel metal2 22904 21448 22904 21448 0 _0171_
rlabel metal2 23016 21168 23016 21168 0 _0172_
rlabel metal2 31864 20720 31864 20720 0 _0173_
rlabel metal2 30744 19600 30744 19600 0 _0174_
rlabel metal2 32088 17864 32088 17864 0 _0175_
rlabel metal2 31416 17528 31416 17528 0 _0176_
rlabel metal2 30016 16632 30016 16632 0 _0177_
rlabel metal2 28840 17640 28840 17640 0 _0178_
rlabel metal2 29624 18536 29624 18536 0 _0179_
rlabel metal2 31808 18088 31808 18088 0 _0180_
rlabel metal2 30408 17752 30408 17752 0 _0181_
rlabel metal2 31304 17304 31304 17304 0 _0182_
rlabel metal2 26152 17248 26152 17248 0 _0183_
rlabel metal3 30296 16800 30296 16800 0 _0184_
rlabel metal3 26880 14392 26880 14392 0 _0185_
rlabel metal3 17808 13944 17808 13944 0 _0186_
rlabel metal3 17808 14504 17808 14504 0 _0187_
rlabel metal2 18648 17640 18648 17640 0 _0188_
rlabel metal2 21672 15904 21672 15904 0 _0189_
rlabel metal3 19600 15960 19600 15960 0 _0190_
rlabel metal3 18312 15512 18312 15512 0 _0191_
rlabel metal2 18424 15848 18424 15848 0 _0192_
rlabel metal2 19320 17248 19320 17248 0 _0193_
rlabel metal2 18648 16856 18648 16856 0 _0194_
rlabel metal2 18760 16408 18760 16408 0 _0195_
rlabel metal2 17808 17752 17808 17752 0 _0196_
rlabel metal2 18984 14728 18984 14728 0 _0197_
rlabel metal3 23576 15960 23576 15960 0 _0198_
rlabel metal2 27720 17528 27720 17528 0 _0199_
rlabel metal4 27048 16688 27048 16688 0 _0200_
rlabel metal2 23464 17136 23464 17136 0 _0201_
rlabel metal2 22232 15512 22232 15512 0 _0202_
rlabel metal2 3304 8680 3304 8680 0 _0203_
rlabel metal2 2856 10192 2856 10192 0 _0204_
rlabel metal2 2856 7616 2856 7616 0 _0205_
rlabel metal2 7616 10584 7616 10584 0 _0206_
rlabel metal2 3528 8232 3528 8232 0 _0207_
rlabel metal2 3192 10192 3192 10192 0 _0208_
rlabel metal2 3976 9800 3976 9800 0 _0209_
rlabel metal2 24528 23016 24528 23016 0 _0210_
rlabel metal2 21560 23184 21560 23184 0 _0211_
rlabel metal2 26208 16632 26208 16632 0 _0212_
rlabel metal2 10248 6440 10248 6440 0 _0213_
rlabel metal2 16296 9520 16296 9520 0 _0214_
rlabel metal2 11480 9912 11480 9912 0 _0215_
rlabel metal2 26432 17528 26432 17528 0 _0216_
rlabel metal2 25872 16072 25872 16072 0 _0217_
rlabel metal2 12488 8960 12488 8960 0 _0218_
rlabel metal2 11144 6440 11144 6440 0 _0219_
rlabel metal2 10640 6664 10640 6664 0 _0220_
rlabel metal2 13160 16072 13160 16072 0 _0221_
rlabel metal2 11592 14056 11592 14056 0 _0222_
rlabel metal2 10808 6664 10808 6664 0 _0223_
rlabel metal2 10528 5992 10528 5992 0 _0224_
rlabel metal2 12600 5656 12600 5656 0 _0225_
rlabel metal2 12152 5376 12152 5376 0 _0226_
rlabel metal2 13664 3528 13664 3528 0 _0227_
rlabel metal2 19432 7392 19432 7392 0 _0228_
rlabel metal2 14168 5768 14168 5768 0 _0229_
rlabel metal2 17528 22904 17528 22904 0 _0230_
rlabel metal2 17976 6048 17976 6048 0 _0231_
rlabel metal2 17752 6608 17752 6608 0 _0232_
rlabel metal2 17304 5936 17304 5936 0 _0233_
rlabel metal2 16968 3696 16968 3696 0 _0234_
rlabel metal2 16968 5040 16968 5040 0 _0235_
rlabel metal2 18984 6384 18984 6384 0 _0236_
rlabel metal2 19936 5096 19936 5096 0 _0237_
rlabel metal3 23128 18536 23128 18536 0 _0238_
rlabel metal2 23800 18480 23800 18480 0 _0239_
rlabel metal2 23408 16408 23408 16408 0 _0240_
rlabel metal3 16688 10584 16688 10584 0 _0241_
rlabel metal2 24360 9128 24360 9128 0 _0242_
rlabel metal3 23744 7672 23744 7672 0 _0243_
rlabel metal2 17416 7392 17416 7392 0 _0244_
rlabel metal2 18200 9464 18200 9464 0 _0245_
rlabel metal3 19656 9800 19656 9800 0 _0246_
rlabel metal2 15176 10024 15176 10024 0 _0247_
rlabel metal2 24136 5040 24136 5040 0 _0248_
rlabel metal2 23744 8232 23744 8232 0 _0249_
rlabel metal3 17864 6440 17864 6440 0 _0250_
rlabel metal2 16912 6776 16912 6776 0 _0251_
rlabel metal2 15680 9912 15680 9912 0 _0252_
rlabel metal2 24472 6944 24472 6944 0 _0253_
rlabel metal2 18088 7952 18088 7952 0 _0254_
rlabel metal2 17360 7672 17360 7672 0 _0255_
rlabel metal2 17864 9912 17864 9912 0 _0256_
rlabel metal2 26376 5152 26376 5152 0 _0257_
rlabel metal3 21952 8008 21952 8008 0 _0258_
rlabel metal2 19544 7952 19544 7952 0 _0259_
rlabel metal2 20664 9912 20664 9912 0 _0260_
rlabel metal2 20160 9912 20160 9912 0 _0261_
rlabel metal2 23576 11032 23576 11032 0 _0262_
rlabel metal2 26152 9352 26152 9352 0 _0263_
rlabel metal2 24808 7728 24808 7728 0 _0264_
rlabel metal2 24808 9128 24808 9128 0 _0265_
rlabel metal3 23856 9688 23856 9688 0 _0266_
rlabel metal2 25256 10304 25256 10304 0 _0267_
rlabel metal2 23912 10136 23912 10136 0 _0268_
rlabel metal2 28616 5656 28616 5656 0 _0269_
rlabel metal2 26824 9352 26824 9352 0 _0270_
rlabel metal2 26208 9912 26208 9912 0 _0271_
rlabel metal2 26712 10248 26712 10248 0 _0272_
rlabel metal2 28056 5824 28056 5824 0 _0273_
rlabel metal2 29624 7728 29624 7728 0 _0274_
rlabel metal2 25816 9016 25816 9016 0 _0275_
rlabel metal3 27272 9688 27272 9688 0 _0276_
rlabel metal2 29176 6160 29176 6160 0 _0277_
rlabel metal2 29400 6496 29400 6496 0 _0278_
rlabel metal3 28952 9240 28952 9240 0 _0279_
rlabel metal2 22568 9856 22568 9856 0 _0280_
rlabel metal2 28672 12152 28672 12152 0 _0281_
rlabel metal2 28056 10920 28056 10920 0 _0282_
rlabel metal2 28056 19320 28056 19320 0 _0283_
rlabel metal2 27720 16464 27720 16464 0 _0284_
rlabel metal2 28112 16072 28112 16072 0 _0285_
rlabel metal3 26040 6664 26040 6664 0 _0286_
rlabel metal2 22792 6552 22792 6552 0 _0287_
rlabel metal2 27832 6776 27832 6776 0 _0288_
rlabel metal3 21952 7560 21952 7560 0 _0289_
rlabel metal2 21728 6664 21728 6664 0 _0290_
rlabel metal2 23464 6272 23464 6272 0 _0291_
rlabel metal2 22344 6328 22344 6328 0 _0292_
rlabel metal2 24584 7056 24584 7056 0 _0293_
rlabel metal3 22960 7448 22960 7448 0 _0294_
rlabel metal2 22456 6776 22456 6776 0 _0295_
rlabel metal2 23520 6776 23520 6776 0 _0296_
rlabel metal2 23576 6216 23576 6216 0 _0297_
rlabel metal3 23800 5096 23800 5096 0 _0298_
rlabel metal2 24920 4984 24920 4984 0 _0299_
rlabel metal2 26040 5152 26040 5152 0 _0300_
rlabel metal2 25480 5432 25480 5432 0 _0301_
rlabel metal2 25592 7000 25592 7000 0 _0302_
rlabel metal2 26040 5880 26040 5880 0 _0303_
rlabel metal2 31976 8232 31976 8232 0 _0304_
rlabel metal2 27832 7504 27832 7504 0 _0305_
rlabel metal2 27608 5488 27608 5488 0 _0306_
rlabel metal3 28560 5096 28560 5096 0 _0307_
rlabel metal2 31696 6552 31696 6552 0 _0308_
rlabel metal2 29792 5096 29792 5096 0 _0309_
rlabel metal3 29624 5880 29624 5880 0 _0310_
rlabel metal2 31640 4648 31640 4648 0 _0311_
rlabel metal2 32200 4368 32200 4368 0 _0312_
rlabel metal3 29176 6104 29176 6104 0 _0313_
rlabel metal2 30576 6664 30576 6664 0 _0314_
rlabel metal2 31584 6776 31584 6776 0 _0315_
rlabel metal2 28728 6776 28728 6776 0 _0316_
rlabel metal3 31360 7336 31360 7336 0 _0317_
rlabel metal2 23240 8848 23240 8848 0 _0318_
rlabel metal2 31864 9184 31864 9184 0 _0319_
rlabel metal4 22568 27944 22568 27944 0 _0320_
rlabel metal2 23464 29904 23464 29904 0 _0321_
rlabel metal2 24360 28168 24360 28168 0 _0322_
rlabel metal2 20664 22792 20664 22792 0 _0323_
rlabel metal2 17584 24808 17584 24808 0 _0324_
rlabel metal2 16184 22960 16184 22960 0 _0325_
rlabel metal3 18368 22904 18368 22904 0 _0326_
rlabel metal3 23184 28056 23184 28056 0 _0327_
rlabel metal2 15960 29568 15960 29568 0 _0328_
rlabel metal2 12600 28336 12600 28336 0 _0329_
rlabel metal2 16632 29120 16632 29120 0 _0330_
rlabel metal3 18760 24696 18760 24696 0 _0331_
rlabel metal2 19432 24528 19432 24528 0 _0332_
rlabel metal2 18760 24976 18760 24976 0 _0333_
rlabel metal2 18984 23128 18984 23128 0 _0334_
rlabel metal2 16520 22792 16520 22792 0 _0335_
rlabel metal2 19376 22904 19376 22904 0 _0336_
rlabel metal2 14168 23464 14168 23464 0 _0337_
rlabel metal3 18760 23128 18760 23128 0 _0338_
rlabel metal2 19208 21280 19208 21280 0 _0339_
rlabel metal2 19208 22456 19208 22456 0 _0340_
rlabel metal2 19208 26208 19208 26208 0 _0341_
rlabel metal2 19600 20776 19600 20776 0 _0342_
rlabel metal2 10864 16856 10864 16856 0 _0343_
rlabel metal2 17640 20608 17640 20608 0 _0344_
rlabel metal2 19544 14224 19544 14224 0 _0345_
rlabel metal2 17976 13832 17976 13832 0 _0346_
rlabel metal2 14504 14056 14504 14056 0 _0347_
rlabel metal3 20860 17080 20860 17080 0 _0348_
rlabel metal2 15960 18312 15960 18312 0 _0349_
rlabel metal2 16464 19992 16464 19992 0 _0350_
rlabel metal3 22512 18984 22512 18984 0 _0351_
rlabel metal3 19096 19096 19096 19096 0 _0352_
rlabel metal2 18312 20664 18312 20664 0 _0353_
rlabel metal2 21784 22120 21784 22120 0 _0354_
rlabel metal2 22232 29344 22232 29344 0 _0355_
rlabel metal2 22568 29680 22568 29680 0 _0356_
rlabel metal2 21336 23408 21336 23408 0 _0357_
rlabel metal2 20440 30240 20440 30240 0 _0358_
rlabel metal2 16744 13776 16744 13776 0 _0359_
rlabel metal2 14952 12880 14952 12880 0 _0360_
rlabel metal2 10248 15624 10248 15624 0 _0361_
rlabel metal2 10696 14616 10696 14616 0 _0362_
rlabel metal3 5880 15288 5880 15288 0 _0363_
rlabel metal2 7896 14896 7896 14896 0 _0364_
rlabel metal2 8232 14392 8232 14392 0 _0365_
rlabel metal2 6776 14504 6776 14504 0 _0366_
rlabel metal3 7280 15288 7280 15288 0 _0367_
rlabel metal2 5992 16128 5992 16128 0 _0368_
rlabel metal3 6496 15512 6496 15512 0 _0369_
rlabel metal2 4088 16968 4088 16968 0 _0370_
rlabel metal2 5096 15568 5096 15568 0 _0371_
rlabel metal2 3192 18256 3192 18256 0 _0372_
rlabel metal2 4312 15960 4312 15960 0 _0373_
rlabel metal3 5544 19992 5544 19992 0 _0374_
rlabel metal2 4424 17192 4424 17192 0 _0375_
rlabel metal2 4984 16912 4984 16912 0 _0376_
rlabel metal3 4648 18424 4648 18424 0 _0377_
rlabel metal3 3640 18424 3640 18424 0 _0378_
rlabel metal2 4312 20496 4312 20496 0 _0379_
rlabel metal3 4928 19432 4928 19432 0 _0380_
rlabel metal3 7672 20776 7672 20776 0 _0381_
rlabel metal3 6160 21560 6160 21560 0 _0382_
rlabel metal3 7840 21672 7840 21672 0 _0383_
rlabel metal2 5768 21280 5768 21280 0 _0384_
rlabel metal2 8232 18704 8232 18704 0 _0385_
rlabel metal2 6664 20888 6664 20888 0 _0386_
rlabel metal2 6216 21056 6216 21056 0 _0387_
rlabel metal2 8792 19684 8792 19684 0 _0388_
rlabel metal2 7896 20384 7896 20384 0 _0389_
rlabel metal2 10696 19880 10696 19880 0 _0390_
rlabel metal2 10360 19544 10360 19544 0 _0391_
rlabel metal2 10920 17752 10920 17752 0 _0392_
rlabel metal3 11592 18424 11592 18424 0 _0393_
rlabel metal2 13664 19208 13664 19208 0 _0394_
rlabel metal2 11312 18536 11312 18536 0 _0395_
rlabel metal3 15848 18368 15848 18368 0 _0396_
rlabel metal2 13384 18480 13384 18480 0 _0397_
rlabel metal3 15064 18424 15064 18424 0 _0398_
rlabel metal2 15064 18648 15064 18648 0 _0399_
rlabel metal3 14728 19992 14728 19992 0 _0400_
rlabel metal2 14056 19992 14056 19992 0 _0401_
rlabel metal3 10080 28392 10080 28392 0 _0402_
rlabel metal2 15176 18760 15176 18760 0 _0403_
rlabel metal3 15512 22456 15512 22456 0 _0404_
rlabel metal2 12656 22232 12656 22232 0 _0405_
rlabel metal2 7000 24080 7000 24080 0 _0406_
rlabel metal2 8344 25144 8344 25144 0 _0407_
rlabel metal2 12600 25816 12600 25816 0 _0408_
rlabel metal2 8008 23968 8008 23968 0 _0409_
rlabel metal2 5320 23184 5320 23184 0 _0410_
rlabel metal2 11928 24472 11928 24472 0 _0411_
rlabel metal2 11928 26152 11928 26152 0 _0412_
rlabel metal2 5600 23240 5600 23240 0 _0413_
rlabel metal2 7392 25480 7392 25480 0 _0414_
rlabel metal3 8064 23688 8064 23688 0 _0415_
rlabel metal2 6160 16968 6160 16968 0 _0416_
rlabel metal2 8288 17080 8288 17080 0 _0417_
rlabel metal2 7784 24080 7784 24080 0 _0418_
rlabel metal2 7672 26712 7672 26712 0 _0419_
rlabel metal2 17472 25480 17472 25480 0 _0420_
rlabel metal2 18536 24472 18536 24472 0 _0421_
rlabel metal2 5208 26544 5208 26544 0 _0422_
rlabel metal3 5936 26152 5936 26152 0 _0423_
rlabel metal3 5712 17080 5712 17080 0 _0424_
rlabel metal3 9632 25256 9632 25256 0 _0425_
rlabel metal3 7672 27048 7672 27048 0 _0426_
rlabel metal3 5488 27160 5488 27160 0 _0427_
rlabel metal2 6776 24584 6776 24584 0 _0428_
rlabel metal2 6664 23968 6664 23968 0 _0429_
rlabel metal2 6944 24920 6944 24920 0 _0430_
rlabel metal2 12376 27384 12376 27384 0 _0431_
rlabel metal2 5712 17080 5712 17080 0 _0432_
rlabel metal2 6440 27888 6440 27888 0 _0433_
rlabel metal3 5096 28728 5096 28728 0 _0434_
rlabel metal2 6272 27832 6272 27832 0 _0435_
rlabel metal2 7560 27328 7560 27328 0 _0436_
rlabel metal2 7336 17752 7336 17752 0 _0437_
rlabel metal2 6552 25396 6552 25396 0 _0438_
rlabel metal2 6384 25592 6384 25592 0 _0439_
rlabel metal2 9296 23240 9296 23240 0 _0440_
rlabel metal2 10024 25480 10024 25480 0 _0441_
rlabel metal2 9576 24808 9576 24808 0 _0442_
rlabel metal2 6440 24304 6440 24304 0 _0443_
rlabel metal2 3976 24640 3976 24640 0 _0444_
rlabel metal2 4424 25592 4424 25592 0 _0445_
rlabel metal2 8624 23352 8624 23352 0 _0446_
rlabel metal2 10584 26936 10584 26936 0 _0447_
rlabel metal2 11032 25760 11032 25760 0 _0448_
rlabel metal2 10584 25256 10584 25256 0 _0449_
rlabel metal3 10696 25368 10696 25368 0 _0450_
rlabel metal2 9744 26824 9744 26824 0 _0451_
rlabel metal2 10024 27720 10024 27720 0 _0452_
rlabel metal3 16744 23184 16744 23184 0 _0453_
rlabel metal2 11256 24808 11256 24808 0 _0454_
rlabel metal2 11144 26600 11144 26600 0 _0455_
rlabel metal2 10696 27272 10696 27272 0 _0456_
rlabel metal2 16856 25984 16856 25984 0 _0457_
rlabel metal4 16184 24696 16184 24696 0 _0458_
rlabel metal2 15848 26208 15848 26208 0 _0459_
rlabel metal2 16016 25256 16016 25256 0 _0460_
rlabel metal2 15960 26544 15960 26544 0 _0461_
rlabel metal2 17024 31080 17024 31080 0 _0462_
rlabel metal2 11032 24360 11032 24360 0 _0463_
rlabel metal2 18872 25648 18872 25648 0 _0464_
rlabel metal4 14952 27608 14952 27608 0 _0465_
rlabel metal3 12768 26824 12768 26824 0 _0466_
rlabel metal2 15568 24920 15568 24920 0 _0467_
rlabel metal2 13832 29960 13832 29960 0 _0468_
rlabel metal2 17416 24864 17416 24864 0 _0469_
rlabel metal2 16856 25088 16856 25088 0 _0470_
rlabel metal2 12712 25088 12712 25088 0 _0471_
rlabel metal2 10472 24024 10472 24024 0 _0472_
rlabel metal2 12152 25928 12152 25928 0 _0473_
rlabel metal3 10752 26488 10752 26488 0 _0474_
rlabel metal3 17416 26488 17416 26488 0 _0475_
rlabel metal2 16520 25032 16520 25032 0 _0476_
rlabel metal2 13216 21784 13216 21784 0 _0477_
rlabel metal3 14840 25368 14840 25368 0 _0478_
rlabel metal2 15512 25816 15512 25816 0 _0479_
rlabel metal3 18480 28392 18480 28392 0 _0480_
rlabel metal2 18984 26264 18984 26264 0 _0481_
rlabel metal2 18368 26488 18368 26488 0 _0482_
rlabel metal3 19768 26264 19768 26264 0 _0483_
rlabel metal3 20048 26152 20048 26152 0 _0484_
rlabel metal2 15456 22568 15456 22568 0 _0485_
rlabel metal3 17080 23800 17080 23800 0 _0486_
rlabel metal3 19488 27272 19488 27272 0 _0487_
rlabel metal2 19656 25088 19656 25088 0 _0488_
rlabel metal2 19544 25200 19544 25200 0 _0489_
rlabel metal2 19096 24360 19096 24360 0 _0490_
rlabel metal2 19320 23800 19320 23800 0 _0491_
rlabel metal2 16744 22512 16744 22512 0 _0492_
rlabel metal3 16800 23688 16800 23688 0 _0493_
rlabel metal3 18368 25592 18368 25592 0 _0494_
rlabel metal2 6776 11424 6776 11424 0 _0495_
rlabel metal2 7336 10752 7336 10752 0 _0496_
rlabel metal2 8792 9912 8792 9912 0 _0497_
rlabel metal2 7728 7672 7728 7672 0 _0498_
rlabel metal2 5992 7896 5992 7896 0 _0499_
rlabel metal2 1848 3472 1848 3472 0 _0500_
rlabel metal4 5096 8176 5096 8176 0 _0501_
rlabel metal2 2632 7336 2632 7336 0 _0502_
rlabel metal2 2072 7672 2072 7672 0 _0503_
rlabel metal2 5544 6328 5544 6328 0 _0504_
rlabel metal3 5712 3304 5712 3304 0 _0505_
rlabel metal2 8344 4928 8344 4928 0 _0506_
rlabel metal3 2688 3304 2688 3304 0 _0507_
rlabel metal2 6328 7840 6328 7840 0 _0508_
rlabel metal2 2296 5208 2296 5208 0 _0509_
rlabel metal3 5208 7448 5208 7448 0 _0510_
rlabel metal2 22792 17360 22792 17360 0 clk_i
rlabel metal2 26600 25592 26600 25592 0 clknet_0_clk_i
rlabel metal3 9296 12936 9296 12936 0 clknet_3_0__leaf_clk_i
rlabel metal2 17864 7392 17864 7392 0 clknet_3_1__leaf_clk_i
rlabel metal2 2296 29736 2296 29736 0 clknet_3_2__leaf_clk_i
rlabel metal2 16856 19152 16856 19152 0 clknet_3_3__leaf_clk_i
rlabel metal2 21448 20496 21448 20496 0 clknet_3_4__leaf_clk_i
rlabel metal2 26040 9744 26040 9744 0 clknet_3_5__leaf_clk_i
rlabel metal2 18760 20888 18760 20888 0 clknet_3_6__leaf_clk_i
rlabel metal2 24920 29680 24920 29680 0 clknet_3_7__leaf_clk_i
rlabel metal2 23912 31304 23912 31304 0 custom_setting
rlabel metal2 7392 17416 7392 17416 0 dest\[0\]
rlabel metal3 9576 20888 9576 20888 0 dest\[10\]
rlabel via2 12600 20104 12600 20104 0 dest\[11\]
rlabel metal2 21000 22120 21000 22120 0 dest\[12\]
rlabel metal2 16072 18480 16072 18480 0 dest\[13\]
rlabel metal2 17136 19320 17136 19320 0 dest\[14\]
rlabel metal2 16408 21504 16408 21504 0 dest\[15\]
rlabel metal2 19992 21336 19992 21336 0 dest\[16\]
rlabel metal2 8176 15512 8176 15512 0 dest\[1\]
rlabel metal2 6440 15624 6440 15624 0 dest\[2\]
rlabel metal3 6664 15792 6664 15792 0 dest\[3\]
rlabel metal2 5208 17136 5208 17136 0 dest\[4\]
rlabel metal3 3220 18648 3220 18648 0 dest\[5\]
rlabel metal3 7336 18984 7336 18984 0 dest\[6\]
rlabel metal3 8512 20552 8512 20552 0 dest\[7\]
rlabel metal2 6776 22512 6776 22512 0 dest\[8\]
rlabel metal3 9744 19880 9744 19880 0 dest\[9\]
rlabel metal2 15064 8120 15064 8120 0 dia\[0\]
rlabel metal2 16632 8288 16632 8288 0 dia\[1\]
rlabel metal2 19544 9912 19544 9912 0 dia\[2\]
rlabel metal2 21896 9352 21896 9352 0 dia\[3\]
rlabel metal3 25928 10584 25928 10584 0 dia\[4\]
rlabel metal2 27272 10640 27272 10640 0 dia\[5\]
rlabel metal2 29400 9408 29400 9408 0 dia\[6\]
rlabel metal2 32088 11816 32088 11816 0 dia\[7\]
rlabel metal2 22512 6104 22512 6104 0 dib\[0\]
rlabel metal2 23352 5824 23352 5824 0 dib\[1\]
rlabel metal2 24192 5880 24192 5880 0 dib\[2\]
rlabel metal2 27888 4984 27888 4984 0 dib\[3\]
rlabel metal2 30856 5376 30856 5376 0 dib\[4\]
rlabel metal2 30520 5824 30520 5824 0 dib\[5\]
rlabel metal3 30688 7672 30688 7672 0 dib\[6\]
rlabel metal2 30688 16744 30688 16744 0 dib\[7\]
rlabel metal3 22680 6608 22680 6608 0 io_in[0]
rlabel metal2 32536 7896 32536 7896 0 io_in[1]
rlabel metal3 23968 8344 23968 8344 0 io_in[2]
rlabel metal3 28224 14840 28224 14840 0 io_in[3]
rlabel metal3 31864 17080 31864 17080 0 io_in[4]
rlabel metal2 27328 9576 27328 9576 0 io_in[5]
rlabel metal2 21280 25704 21280 25704 0 io_in[6]
rlabel metal2 19656 31080 19656 31080 0 io_in[7]
rlabel metal2 11704 33418 11704 33418 0 io_out[10]
rlabel metal3 13608 28504 13608 28504 0 io_out[11]
rlabel metal3 15148 28056 15148 28056 0 io_out[12]
rlabel metal2 16856 27832 16856 27832 0 io_out[13]
rlabel metal2 16184 32578 16184 32578 0 io_out[14]
rlabel metal2 17304 32914 17304 32914 0 io_out[15]
rlabel metal2 18424 32746 18424 32746 0 io_out[16]
rlabel metal2 19544 32746 19544 32746 0 io_out[17]
rlabel metal2 20664 33698 20664 33698 0 io_out[18]
rlabel metal2 22344 27776 22344 27776 0 io_out[19]
rlabel metal3 24584 31192 24584 31192 0 io_out[20]
rlabel metal2 24024 31570 24024 31570 0 io_out[21]
rlabel metal2 25144 30898 25144 30898 0 io_out[22]
rlabel metal2 26824 30016 26824 30016 0 io_out[23]
rlabel metal3 29008 28392 29008 28392 0 io_out[24]
rlabel metal2 28504 32186 28504 32186 0 io_out[25]
rlabel metal3 30520 28504 30520 28504 0 io_out[26]
rlabel metal2 30744 30338 30744 30338 0 io_out[27]
rlabel metal2 31248 34328 31248 34328 0 io_out[28]
rlabel metal2 33152 22568 33152 22568 0 io_out[29]
rlabel metal2 30744 24864 30744 24864 0 io_out[30]
rlabel metal2 8008 31472 8008 31472 0 io_out[8]
rlabel metal2 10584 34202 10584 34202 0 io_out[9]
rlabel metal2 7896 11144 7896 11144 0 mar\[0\]
rlabel metal2 6104 8904 6104 8904 0 mar\[1\]
rlabel metal2 22344 18760 22344 18760 0 mc14500.DATA_OUT
rlabel metal3 17752 15288 17752 15288 0 mc14500.IEN_l
rlabel metal2 20384 13832 20384 13832 0 mc14500.OEN_l
rlabel metal2 12936 13384 12936 13384 0 mc14500.X1
rlabel metal2 28280 14168 28280 14168 0 mc14500.instr_l\[0\]
rlabel metal2 29624 12488 29624 12488 0 mc14500.instr_l\[1\]
rlabel metal2 30352 13720 30352 13720 0 mc14500.instr_l\[2\]
rlabel metal2 32536 15400 32536 15400 0 mc14500.instr_l\[3\]
rlabel metal2 22232 13048 22232 13048 0 mc14500.skip
rlabel metal2 31472 18760 31472 18760 0 net1
rlabel metal2 17640 17808 17640 17808 0 net10
rlabel metal2 27496 12152 27496 12152 0 net11
rlabel metal2 23688 4536 23688 4536 0 net12
rlabel metal2 24584 3416 24584 3416 0 net13
rlabel metal2 26264 3808 26264 3808 0 net14
rlabel metal2 28392 3584 28392 3584 0 net15
rlabel metal3 29064 3416 29064 3416 0 net16
rlabel metal2 31304 3808 31304 3808 0 net17
rlabel metal2 32536 4592 32536 4592 0 net18
rlabel metal2 30632 4592 30632 4592 0 net19
rlabel metal3 23688 30968 23688 30968 0 net2
rlabel metal3 9520 27496 9520 27496 0 net20
rlabel metal2 13048 26572 13048 26572 0 net21
rlabel metal2 14168 28224 14168 28224 0 net22
rlabel metal2 15288 25088 15288 25088 0 net23
rlabel metal3 10192 27944 10192 27944 0 net24
rlabel metal2 17752 28392 17752 28392 0 net25
rlabel metal2 17976 29848 17976 29848 0 net26
rlabel metal2 18648 30632 18648 30632 0 net27
rlabel metal3 25816 26768 25816 26768 0 net28
rlabel metal2 15400 25648 15400 25648 0 net29
rlabel metal2 29512 6664 29512 6664 0 net3
rlabel metal2 24360 30072 24360 30072 0 net30
rlabel metal2 24024 27776 24024 27776 0 net31
rlabel metal2 24024 25424 24024 25424 0 net32
rlabel metal2 24472 25872 24472 25872 0 net33
rlabel metal2 19880 24416 19880 24416 0 net34
rlabel metal2 26096 19208 26096 19208 0 net35
rlabel metal3 29400 24024 29400 24024 0 net36
rlabel metal2 22680 21112 22680 21112 0 net37
rlabel metal3 31584 23240 31584 23240 0 net38
rlabel metal2 16016 21784 16016 21784 0 net39
rlabel metal2 31752 12432 31752 12432 0 net4
rlabel metal2 29512 23464 29512 23464 0 net40
rlabel metal2 4816 24024 4816 24024 0 net41
rlabel metal2 8568 29456 8568 29456 0 net42
rlabel metal2 1736 8848 1736 8848 0 net43
rlabel metal2 4648 6720 4648 6720 0 net44
rlabel metal2 1736 5712 1736 5712 0 net45
rlabel metal2 2408 7000 2408 7000 0 net46
rlabel metal2 2016 3416 2016 3416 0 net47
rlabel metal2 5992 6552 5992 6552 0 net48
rlabel metal2 28112 24696 28112 24696 0 net49
rlabel metal2 32424 14168 32424 14168 0 net5
rlabel metal2 11592 8736 11592 8736 0 net50
rlabel metal3 9968 6552 9968 6552 0 net51
rlabel metal2 11928 5600 11928 5600 0 net52
rlabel metal2 9744 3640 9744 3640 0 net53
rlabel metal2 12712 5936 12712 5936 0 net54
rlabel metal3 19712 7560 19712 7560 0 net55
rlabel metal2 19768 4480 19768 4480 0 net56
rlabel metal3 20944 4200 20944 4200 0 net57
rlabel metal2 25480 27888 25480 27888 0 net58
rlabel metal2 16296 25704 16296 25704 0 net59
rlabel metal3 29176 15176 29176 15176 0 net6
rlabel metal3 5488 23240 5488 23240 0 net60
rlabel metal3 7784 26376 7784 26376 0 net61
rlabel metal2 13720 11816 13720 11816 0 net62
rlabel metal2 30184 12432 30184 12432 0 net63
rlabel metal3 29232 11144 29232 11144 0 net64
rlabel metal2 28616 14112 28616 14112 0 net65
rlabel metal2 19656 12656 19656 12656 0 net66
rlabel metal2 2296 31360 2296 31360 0 net67
rlabel metal2 1848 31556 1848 31556 0 net68
rlabel metal2 2968 31556 2968 31556 0 net69
rlabel metal2 32760 12824 32760 12824 0 net7
rlabel metal2 3920 31192 3920 31192 0 net70
rlabel metal2 4536 31976 4536 31976 0 net71
rlabel metal2 4984 31528 4984 31528 0 net72
rlabel metal3 6552 31192 6552 31192 0 net73
rlabel metal3 8624 29960 8624 29960 0 net74
rlabel metal3 26152 12712 26152 12712 0 net8
rlabel metal2 21896 18256 21896 18256 0 net9
rlabel metal2 24136 29512 24136 29512 0 rst_latency\[0\]
rlabel metal2 24584 28336 24584 28336 0 rst_latency\[1\]
rlabel metal2 26376 4368 26376 4368 0 rst_n
rlabel metal2 24304 20888 24304 20888 0 scratch\[0\]
rlabel metal2 24920 23464 24920 23464 0 scratch\[1\]
rlabel metal3 24248 21728 24248 21728 0 scratch\[2\]
rlabel metal2 28168 27496 28168 27496 0 scratch\[3\]
rlabel metal2 23128 25256 23128 25256 0 scratch\[4\]
rlabel metal2 22232 27944 22232 27944 0 scratch\[5\]
rlabel metal2 952 2142 952 2142 0 sram_addr[0]
rlabel metal2 2520 2982 2520 2982 0 sram_addr[1]
rlabel metal2 4088 2086 4088 2086 0 sram_addr[2]
rlabel metal2 5880 3640 5880 3640 0 sram_addr[3]
rlabel metal2 7224 2058 7224 2058 0 sram_addr[4]
rlabel metal2 8792 2058 8792 2058 0 sram_addr[5]
rlabel metal3 28056 25704 28056 25704 0 sram_gwe
rlabel metal2 10360 2478 10360 2478 0 sram_in[0]
rlabel metal2 11928 2058 11928 2058 0 sram_in[1]
rlabel metal2 13496 854 13496 854 0 sram_in[2]
rlabel metal2 15064 3206 15064 3206 0 sram_in[3]
rlabel metal2 16632 2058 16632 2058 0 sram_in[4]
rlabel metal2 18200 2198 18200 2198 0 sram_in[5]
rlabel metal2 19768 2058 19768 2058 0 sram_in[6]
rlabel metal2 21336 2058 21336 2058 0 sram_in[7]
rlabel metal3 24976 3416 24976 3416 0 sram_out[0]
rlabel metal2 24472 854 24472 854 0 sram_out[1]
rlabel metal2 26040 854 26040 854 0 sram_out[2]
rlabel metal2 21112 5544 21112 5544 0 sram_out[3]
rlabel metal3 28672 3528 28672 3528 0 sram_out[4]
rlabel metal2 26600 5488 26600 5488 0 sram_out[5]
rlabel metal2 22120 5320 22120 5320 0 sram_out[6]
rlabel metal2 25032 5432 25032 5432 0 sram_out[7]
<< properties >>
string FIXED_BBOX 0 0 35000 35000
<< end >>
