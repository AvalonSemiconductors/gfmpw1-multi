module hellorld (io_out,
    rst_n,
    vdd,
    vss,
    wb_clk_i,
    custom_settings);
 output io_out;
 input rst_n;
 inout vdd;
 inout vss;
 input wb_clk_i;
 input [11:0] custom_settings;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire \baud_delay[0] ;
 wire \baud_delay[10] ;
 wire \baud_delay[11] ;
 wire \baud_delay[1] ;
 wire \baud_delay[2] ;
 wire \baud_delay[3] ;
 wire \baud_delay[4] ;
 wire \baud_delay[5] ;
 wire \baud_delay[6] ;
 wire \baud_delay[7] ;
 wire \baud_delay[8] ;
 wire \baud_delay[9] ;
 wire \char_at[0] ;
 wire \char_at[1] ;
 wire \char_at[2] ;
 wire \char_at[3] ;
 wire \char_at[4] ;
 wire \char_at[5] ;
 wire \char_at[6] ;
 wire \char_pointer[0] ;
 wire \char_pointer[1] ;
 wire \char_pointer[2] ;
 wire \char_pointer[3] ;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire \frame_counter[0] ;
 wire \frame_counter[1] ;
 wire \frame_counter[2] ;
 wire \frame_counter[3] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \uart_frame[0] ;
 wire \uart_frame[1] ;
 wire \uart_frame[2] ;
 wire \uart_frame[3] ;
 wire \uart_frame[4] ;
 wire \uart_frame[5] ;
 wire \uart_frame[6] ;
 wire \uart_frame[7] ;
 wire \uart_frame[8] ;
 wire \uart_frame[9] ;

 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__204__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_120_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__217__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_120_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__251__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_120_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__401__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__415__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__416__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__417__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__418__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__421__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__423__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__430__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload1_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input10_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[7]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input11_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[8]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input12_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[9]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input13_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(rst_n));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input1_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input2_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[10]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input3_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[11]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input4_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[1]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input5_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[2]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input6_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[3]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input7_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[4]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input8_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[5]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input9_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[6]));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_11_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_14_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_1_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_20_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_35 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_24_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_24_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_24_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_24_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_24_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_24_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_4_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_7_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_7_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_7_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Left_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Left_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Left_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Left_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Left_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Left_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Left_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Left_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Left_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Left_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Left_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Left_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Left_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Left_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_22_Left_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_23_Left_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_24_Left_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Left_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Left_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Left_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Left_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Left_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Left_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Left_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Left_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _197_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_097_),
    .B(\char_at[6] ),
    .A(\uart_frame[8] ),
    .Y(_116_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _198_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_112_),
    .B(_116_),
    .A(\uart_frame[7] ),
    .Y(_117_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _199_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_117_),
    .Y(_011_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _200_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_112_),
    .B(_098_),
    .A(\uart_frame[9] ),
    .Y(_118_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _201_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_118_),
    .Y(_012_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _202_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\baud_delay[0] ),
    .Y(_119_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _203_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_100_),
    .A(_059_),
    .Y(_120_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _204_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_120_),
    .Y(_121_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _205_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_013_),
    .B(_121_),
    .A(_119_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _206_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\baud_delay[1] ),
    .Y(_122_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _207_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_122_),
    .A(_119_),
    .Y(_123_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _208_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_124_),
    .B(_122_),
    .A(_119_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _209_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_121_),
    .B(_123_),
    .C(_124_),
    .Y(_125_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _210_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_125_),
    .Y(_014_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _211_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_123_),
    .A(\baud_delay[2] ),
    .Y(_126_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _212_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_015_),
    .B(_126_),
    .A(_121_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _213_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\baud_delay[0] ),
    .B(_122_),
    .C(\baud_delay[2] ),
    .D(\baud_delay[3] ),
    .Y(_127_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _214_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\baud_delay[3] ),
    .A(_119_),
    .B(_122_),
    .C(\baud_delay[2] ),
    .Y(_128_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _215_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_129_),
    .B(_128_),
    .A(_127_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _216_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_016_),
    .B(_129_),
    .A(_121_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _217_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_120_),
    .Y(_130_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _218_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_130_),
    .Y(_131_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _219_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_132_),
    .A(\baud_delay[4] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _220_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_133_),
    .B(_127_),
    .A(_132_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _221_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_127_),
    .A(_132_),
    .Y(_134_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _222_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_131_),
    .B(_133_),
    .C(_134_),
    .Y(_135_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _223_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_135_),
    .Y(_017_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _224_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_136_),
    .A(\baud_delay[5] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _225_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_132_),
    .B(_136_),
    .C(_127_),
    .Y(_137_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _226_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_138_),
    .B(_133_),
    .A(\baud_delay[5] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _227_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_131_),
    .B(_137_),
    .C(_138_),
    .Y(_139_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _228_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_139_),
    .Y(_018_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _229_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_137_),
    .A(\baud_delay[6] ),
    .Y(_140_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _230_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_141_),
    .B(_137_),
    .A(\baud_delay[6] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _231_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_131_),
    .B(_140_),
    .C(_141_),
    .Y(_142_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _232_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_142_),
    .Y(_019_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _233_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_143_),
    .B(_140_),
    .A(\baud_delay[7] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _234_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_140_),
    .A(\baud_delay[7] ),
    .Y(_144_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _235_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_131_),
    .B(_143_),
    .C(_144_),
    .Y(_145_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _236_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_145_),
    .Y(_020_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _237_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_146_),
    .B(_144_),
    .A(\baud_delay[8] ));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _238_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\baud_delay[6] ),
    .B(\baud_delay[7] ),
    .C(_137_),
    .Y(_147_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _239_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_148_),
    .B(_147_),
    .A(\baud_delay[8] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _240_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_130_),
    .B(_146_),
    .C(_148_),
    .Y(_149_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _241_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_149_),
    .Y(_021_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _242_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_150_),
    .B(_148_),
    .A(\baud_delay[9] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _243_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_148_),
    .A(\baud_delay[9] ),
    .Y(_151_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _244_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_130_),
    .B(_150_),
    .C(_151_),
    .Y(_152_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _245_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_152_),
    .Y(_022_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _246_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_153_),
    .B(_151_),
    .A(\baud_delay[10] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _247_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_151_),
    .A(\baud_delay[10] ),
    .Y(_154_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _248_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_130_),
    .B(_153_),
    .C(_154_),
    .Y(_155_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _249_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_155_),
    .Y(_023_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _250_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_156_),
    .B(_154_),
    .A(\baud_delay[11] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _251_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_120_),
    .A(\baud_delay[10] ),
    .B(\baud_delay[11] ),
    .C(_151_),
    .Y(_157_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _252_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_024_),
    .B(_157_),
    .A(_156_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _253_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_158_),
    .B(_097_),
    .A(_100_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _254_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_158_),
    .Y(_159_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _255_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_081_),
    .Y(_160_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _256_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_161_),
    .B(net14),
    .A(_159_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _257_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_162_),
    .B(_161_),
    .A(_160_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _258_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_163_),
    .A(\uart_frame[0] ),
    .B(_159_),
    .C(_162_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _259_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_163_),
    .Y(_025_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _260_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_028_),
    .A(_085_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _261_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_158_),
    .A(_081_),
    .Y(_164_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _262_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_165_),
    .A(_101_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _263_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\uart_frame[1] ),
    .B(_164_),
    .C(_165_),
    .D(\uart_frame[0] ),
    .Y(_166_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _264_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_166_),
    .Y(_030_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _265_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\uart_frame[9] ),
    .B(_164_),
    .C(_165_),
    .D(\uart_frame[8] ),
    .Y(_167_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _266_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_167_),
    .Y(_031_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _267_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\frame_counter[0] ),
    .Y(_168_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _268_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_159_),
    .A(_168_),
    .Y(_169_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _269_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_100_),
    .Y(_170_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _270_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_171_),
    .B(_170_),
    .A(_168_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _271_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_171_),
    .A(_160_),
    .Y(_172_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _272_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_172_),
    .A(_169_),
    .Y(_173_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _273_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_173_),
    .Y(_032_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _274_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_174_),
    .B(_170_),
    .A(_098_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _275_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_175_),
    .A(\frame_counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _276_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_059_),
    .A(_175_),
    .B(_168_),
    .C(_170_),
    .Y(_176_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _277_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_176_),
    .A(\frame_counter[1] ),
    .B(_174_),
    .C(_171_),
    .Y(_177_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _278_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_177_),
    .Y(_033_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _279_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_178_),
    .B(_171_),
    .A(_175_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _280_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_178_),
    .A(\frame_counter[2] ),
    .Y(_179_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _281_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_180_),
    .B(_179_),
    .A(_160_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _282_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_034_),
    .C(_180_),
    .B(_178_),
    .A(\frame_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _283_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\frame_counter[2] ),
    .B(\frame_counter[1] ),
    .C(_168_),
    .Y(_181_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _284_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_181_),
    .A(\frame_counter[3] ),
    .Y(_182_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _285_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_183_),
    .B(\frame_counter[3] ),
    .A(_170_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _286_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_184_),
    .B(_183_),
    .A(_160_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _287_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_185_),
    .A(_159_),
    .B(_182_),
    .C(_184_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _288_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_185_),
    .Y(_035_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _289_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_036_),
    .B(_029_),
    .A(_071_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _290_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_086_),
    .A(_090_),
    .Y(_186_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _291_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_186_),
    .Y(_037_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _292_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_187_),
    .B(\frame_counter[1] ),
    .A(\frame_counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _293_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\frame_counter[2] ),
    .B(\frame_counter[0] ),
    .C(_187_),
    .Y(_188_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _294_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_188_),
    .Y(_189_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _295_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[5] ),
    .A(net8),
    .Y(_190_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _296_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[8] ),
    .A(net11),
    .Y(_191_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _297_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[7] ),
    .A(net10),
    .Y(_192_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _298_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[3] ),
    .A(net6),
    .Y(_193_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _299_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_190_),
    .B(_191_),
    .C(_192_),
    .D(_193_),
    .Y(_194_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _300_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[10] ),
    .A(net2),
    .Y(_195_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _301_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[11] ),
    .A(net3),
    .Y(_196_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _302_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[6] ),
    .A(net9),
    .Y(_038_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _303_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[9] ),
    .A(net12),
    .Y(_039_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _304_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_195_),
    .B(_196_),
    .C(_038_),
    .D(_039_),
    .Y(_040_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _305_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[2] ),
    .A(net5),
    .Y(_041_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _306_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[1] ),
    .A(net4),
    .Y(_042_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _307_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net1),
    .A(\baud_delay[0] ),
    .Y(_043_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _308_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\baud_delay[4] ),
    .A(net7),
    .Y(_044_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _309_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_041_),
    .B(_042_),
    .C(_043_),
    .D(_044_),
    .Y(_045_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _310_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_194_),
    .B(_040_),
    .C(_045_),
    .Y(_046_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _311_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_046_),
    .Y(_047_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _312_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_048_),
    .A(\char_pointer[1] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _313_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_049_),
    .A(_189_),
    .B(_047_),
    .C(_048_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _314_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_189_),
    .Y(_050_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _315_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_047_),
    .Y(_051_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _316_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_052_),
    .B(\char_pointer[2] ),
    .A(\char_pointer[3] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _317_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_053_),
    .A(\char_pointer[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _318_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_053_),
    .A(\char_pointer[1] ),
    .Y(_054_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _319_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_055_),
    .B(_054_),
    .A(_052_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _320_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\char_pointer[0] ),
    .A(_048_),
    .Y(_056_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _321_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_050_),
    .B(_051_),
    .C(_055_),
    .D(_056_),
    .Y(_057_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _322_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_058_),
    .A(net13));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _323_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_058_),
    .Y(_059_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _324_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_060_),
    .A(_049_),
    .B(_057_),
    .C(_059_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _325_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_027_),
    .A(_060_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _326_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_053_),
    .B(_188_),
    .C(_046_),
    .D(_055_),
    .Y(_061_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _327_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_062_),
    .A(_188_),
    .B(_046_),
    .C(_053_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _328_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\char_pointer[0] ),
    .A(\char_pointer[1] ),
    .Y(_063_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _329_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_063_),
    .A(\char_pointer[2] ),
    .Y(_064_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _330_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\char_pointer[3] ),
    .A(_189_),
    .B(_047_),
    .C(_064_),
    .Y(_065_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _331_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_052_),
    .B(_054_),
    .C(_064_),
    .D(\char_pointer[3] ),
    .Y(_066_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _332_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_058_),
    .A(_189_),
    .B(_047_),
    .C(_066_),
    .Y(_067_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _333_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_068_),
    .B(_067_),
    .A(_065_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _334_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_068_),
    .Y(_069_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _335_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_070_),
    .B(_063_),
    .A(\char_pointer[2] ));
 gf180mcu_as_sc_mcu7t3v3__aoi31_4 _336_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_050_),
    .B(_051_),
    .C(_064_),
    .D(_070_),
    .Y(_071_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _337_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_072_),
    .A(_050_),
    .B(_051_),
    .C(\char_pointer[2] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _338_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_073_),
    .B(_072_),
    .A(_071_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _339_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_073_),
    .A(_069_),
    .Y(_074_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _340_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_027_),
    .B(_061_),
    .C(_062_),
    .D(_074_),
    .Y(_075_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _341_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_076_),
    .A(_061_),
    .B(_062_),
    .C(_059_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _342_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_076_),
    .Y(_077_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _343_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_078_),
    .A(_060_),
    .B(_077_),
    .C(_069_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _344_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_057_),
    .A(_049_),
    .Y(_079_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _345_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_026_),
    .A(_076_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _346_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_080_),
    .A(_079_),
    .B(_026_),
    .C(_068_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _347_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net13),
    .Y(_081_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _348_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_081_),
    .B(_071_),
    .C(_072_),
    .Y(_082_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _349_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_082_),
    .B(_080_),
    .A(_078_),
    .Y(_083_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _350_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_083_),
    .A(_075_),
    .Y(_084_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _351_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_084_),
    .Y(_000_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _352_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_069_),
    .Y(_029_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _353_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_082_),
    .Y(_085_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _354_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_086_),
    .B(_085_),
    .A(_029_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _355_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_087_),
    .B(_086_),
    .A(_079_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _356_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_001_),
    .B(_087_),
    .A(_075_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _357_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_088_),
    .B(_077_),
    .A(_085_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _358_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_060_),
    .B(_085_),
    .C(_077_),
    .Y(_089_),
    .D(_069_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _359_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_026_),
    .A(_079_),
    .Y(_090_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _360_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_091_),
    .B(_090_),
    .A(_073_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _361_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_029_),
    .B(_088_),
    .C(_089_),
    .D(_091_),
    .Y(_092_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _362_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_092_),
    .Y(_002_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _363_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_080_),
    .A(_071_),
    .B(_072_),
    .C(_026_),
    .Y(_093_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _364_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_094_),
    .B(_090_),
    .A(_074_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _365_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_075_),
    .B(_093_),
    .C(_094_),
    .Y(_095_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _366_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_095_),
    .Y(_003_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _367_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_089_),
    .A(_060_),
    .B(_074_),
    .C(_077_),
    .Y(_096_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _368_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_096_),
    .Y(_004_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _369_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_050_),
    .Y(_097_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _370_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_097_),
    .Y(_098_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _371_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_098_),
    .B(\char_at[0] ),
    .A(\uart_frame[2] ),
    .Y(_099_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _372_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_051_),
    .Y(_100_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _373_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_100_),
    .A(_081_),
    .Y(_101_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _374_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_101_),
    .Y(_102_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _375_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_102_),
    .B(_099_),
    .A(\uart_frame[1] ),
    .Y(_103_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _376_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_103_),
    .Y(_005_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _377_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_098_),
    .B(\char_at[1] ),
    .A(\uart_frame[3] ),
    .Y(_104_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _378_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_102_),
    .B(_104_),
    .A(\uart_frame[2] ),
    .Y(_105_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _379_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_105_),
    .Y(_006_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _380_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_097_),
    .Y(_106_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _381_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_106_),
    .B(\char_at[2] ),
    .A(\uart_frame[4] ),
    .Y(_107_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _382_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_102_),
    .B(_107_),
    .A(\uart_frame[3] ),
    .Y(_108_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _383_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_108_),
    .Y(_007_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _384_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_106_),
    .B(\char_at[3] ),
    .A(\uart_frame[5] ),
    .Y(_109_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _385_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_102_),
    .B(_109_),
    .A(\uart_frame[4] ),
    .Y(_110_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _386_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_110_),
    .Y(_008_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _387_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_106_),
    .B(\char_at[4] ),
    .A(\uart_frame[6] ),
    .Y(_111_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _388_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_101_),
    .Y(_112_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _389_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_112_),
    .B(_111_),
    .A(\uart_frame[5] ),
    .Y(_113_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _390_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_113_),
    .Y(_009_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _391_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_106_),
    .B(\char_at[5] ),
    .A(\uart_frame[7] ),
    .Y(_114_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _392_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_112_),
    .B(_114_),
    .A(\uart_frame[6] ),
    .Y(_115_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _393_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_115_),
    .Y(_010_));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _394_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_005_),
    .Q(\uart_frame[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _395_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_006_),
    .Q(\uart_frame[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _396_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_007_),
    .Q(\uart_frame[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _397_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_008_),
    .Q(\uart_frame[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _398_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_009_),
    .Q(\uart_frame[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _399_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_010_),
    .Q(\uart_frame[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _400_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_011_),
    .Q(\uart_frame[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _401_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_012_),
    .Q(\uart_frame[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _402_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_013_),
    .Q(\baud_delay[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _403_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_014_),
    .Q(\baud_delay[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _404_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_015_),
    .Q(\baud_delay[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _405_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_016_),
    .Q(\baud_delay[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _406_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_017_),
    .Q(\baud_delay[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _407_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_018_),
    .Q(\baud_delay[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _408_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_019_),
    .Q(\baud_delay[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _409_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_020_),
    .Q(\baud_delay[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _410_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_021_),
    .Q(\baud_delay[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _411_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_022_),
    .Q(\baud_delay[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _412_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_023_),
    .Q(\baud_delay[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _413_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_024_),
    .Q(\baud_delay[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _414_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_025_),
    .Q(net14));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _415_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_026_),
    .Q(\char_pointer[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _416_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_027_),
    .Q(\char_pointer[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _417_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_028_),
    .Q(\char_pointer[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _418_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_029_),
    .Q(\char_pointer[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _419_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_030_),
    .Q(\uart_frame[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _420_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_031_),
    .Q(\uart_frame[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _421_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_032_),
    .Q(\frame_counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _422_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_033_),
    .Q(\frame_counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _423_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_034_),
    .Q(\frame_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _424_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_035_),
    .Q(\frame_counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _425_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_000_),
    .Q(\char_at[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _426_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_001_),
    .Q(\char_at[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _427_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_002_),
    .Q(\char_at[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _428_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_003_),
    .Q(\char_at[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _429_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_004_),
    .Q(\char_at[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _430_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_036_),
    .Q(\char_at[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _431_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_037_),
    .Q(\char_at[4] ));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(wb_clk_i),
    .Y(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_2_0__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_2_1__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_2_2__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_2_3__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload0 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload1 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input1 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[0]),
    .Y(net1));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[7]),
    .Y(net10));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[8]),
    .Y(net11));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[9]),
    .Y(net12));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(rst_n),
    .Y(net13));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[10]),
    .Y(net2));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input3 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[11]),
    .Y(net3));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[1]),
    .Y(net4));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[2]),
    .Y(net5));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[3]),
    .Y(net6));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[4]),
    .Y(net7));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[5]),
    .Y(net8));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[6]),
    .Y(net9));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net14),
    .Y(io_out));
endmodule
