VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ue1
  CLASS BLOCK ;
  FOREIGN ue1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    ANTENNADIFFAREA 0.877000 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 7.840 120.000 8.400 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 36.960 120.000 37.520 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 51.520 120.000 52.080 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 66.080 120.000 66.640 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 80.640 120.000 81.200 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 95.200 120.000 95.760 ;
    END
  END io_in[4]
  PIN io_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 109.760 120.000 110.320 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 8.960 116.000 9.520 120.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 116.000 20.720 120.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 116.000 31.920 120.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 116.000 43.120 120.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 116.000 54.320 120.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 116.000 65.520 120.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 116.000 76.720 120.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 116.000 87.920 120.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 116.000 99.120 120.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 116.000 110.320 120.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 22.400 120.000 22.960 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.220 15.380 20.820 102.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 45.820 15.380 47.420 102.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 72.420 15.380 74.020 102.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.020 15.380 100.620 102.220 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 32.520 15.380 34.120 102.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.120 15.380 60.720 102.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 85.720 15.380 87.320 102.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.320 15.380 113.920 102.220 ;
    END
  END vss
  OBS
      LAYER Pwell ;
        RECT 6.290 100.150 113.550 102.350 ;
      LAYER Nwell ;
        RECT 6.290 95.850 113.550 100.150 ;
      LAYER Pwell ;
        RECT 6.290 92.310 113.550 95.850 ;
      LAYER Nwell ;
        RECT 6.290 88.010 113.550 92.310 ;
      LAYER Pwell ;
        RECT 6.290 84.470 113.550 88.010 ;
      LAYER Nwell ;
        RECT 6.290 80.170 113.550 84.470 ;
      LAYER Pwell ;
        RECT 6.290 76.630 113.550 80.170 ;
      LAYER Nwell ;
        RECT 6.290 72.330 113.550 76.630 ;
      LAYER Pwell ;
        RECT 6.290 68.790 113.550 72.330 ;
      LAYER Nwell ;
        RECT 6.290 64.490 113.550 68.790 ;
      LAYER Pwell ;
        RECT 6.290 60.950 113.550 64.490 ;
      LAYER Nwell ;
        RECT 6.290 56.650 113.550 60.950 ;
      LAYER Pwell ;
        RECT 6.290 53.110 113.550 56.650 ;
      LAYER Nwell ;
        RECT 6.290 48.810 113.550 53.110 ;
      LAYER Pwell ;
        RECT 6.290 45.270 113.550 48.810 ;
      LAYER Nwell ;
        RECT 6.290 40.970 113.550 45.270 ;
      LAYER Pwell ;
        RECT 6.290 37.430 113.550 40.970 ;
      LAYER Nwell ;
        RECT 6.290 33.130 113.550 37.430 ;
      LAYER Pwell ;
        RECT 6.290 29.590 113.550 33.130 ;
      LAYER Nwell ;
        RECT 6.290 25.290 113.550 29.590 ;
      LAYER Pwell ;
        RECT 6.290 21.750 113.550 25.290 ;
      LAYER Nwell ;
        RECT 6.290 17.450 113.550 21.750 ;
      LAYER Pwell ;
        RECT 6.290 15.250 113.550 17.450 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 113.920 102.220 ;
      LAYER Metal2 ;
        RECT 9.820 115.700 19.860 116.340 ;
        RECT 21.020 115.700 31.060 116.340 ;
        RECT 32.220 115.700 42.260 116.340 ;
        RECT 43.420 115.700 53.460 116.340 ;
        RECT 54.620 115.700 64.660 116.340 ;
        RECT 65.820 115.700 75.860 116.340 ;
        RECT 77.020 115.700 87.060 116.340 ;
        RECT 88.220 115.700 98.260 116.340 ;
        RECT 99.420 115.700 109.460 116.340 ;
        RECT 110.620 115.700 113.780 116.340 ;
        RECT 9.100 7.930 113.780 115.700 ;
      LAYER Metal3 ;
        RECT 14.090 109.460 115.700 110.180 ;
        RECT 14.090 96.060 116.000 109.460 ;
        RECT 14.090 94.900 115.700 96.060 ;
        RECT 14.090 81.500 116.000 94.900 ;
        RECT 14.090 80.340 115.700 81.500 ;
        RECT 14.090 66.940 116.000 80.340 ;
        RECT 14.090 65.780 115.700 66.940 ;
        RECT 14.090 52.380 116.000 65.780 ;
        RECT 14.090 51.220 115.700 52.380 ;
        RECT 14.090 37.820 116.000 51.220 ;
        RECT 14.090 36.660 115.700 37.820 ;
        RECT 14.090 23.260 116.000 36.660 ;
        RECT 14.090 22.100 115.700 23.260 ;
        RECT 14.090 8.700 116.000 22.100 ;
        RECT 14.090 7.980 115.700 8.700 ;
      LAYER Metal4 ;
        RECT 51.660 61.130 51.940 65.430 ;
  END
END ue1
END LIBRARY

