* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuD

* Black-box entry subcircuit for wrapped_pdp11 abstract view
.subckt wrapped_pdp11 custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[12]
+ custom_settings[13] custom_settings[14] custom_settings[15] custom_settings[16]
+ custom_settings[17] custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[2]
+ custom_settings[3] custom_settings[4] custom_settings[5] custom_settings[6] custom_settings[7]
+ custom_settings[8] custom_settings[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6]
+ io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28]
+ io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for avali_logo abstract view
.subckt avali_logo vss vdd
.ends

* Black-box entry subcircuit for wrapped_sid abstract view
.subckt wrapped_sid io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[2] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_mc14500 abstract view
.subckt wrapped_mc14500 SDI clk_i custom_setting io_in[0] io_in[1] io_in[2] io_in[3]
+ io_in[4] io_in[5] io_in[6] io_in[7] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28]
+ io_out[29] io_out[2] io_out[30] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] rst_n sram_addr[0] sram_addr[1] sram_addr[2] sram_addr[3] sram_addr[4]
+ sram_addr[5] sram_gwe sram_in[0] sram_in[1] sram_in[2] sram_in[3] sram_in[4] sram_in[5]
+ sram_in[6] sram_in[7] sram_out[0] sram_out[1] sram_out[2] sram_out[3] sram_out[4]
+ sram_out[5] sram_out[6] sram_out[7] vdd vss
.ends

* Black-box entry subcircuit for blinker abstract view
.subckt blinker io_out[0] io_out[1] io_out[2] rst_n vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for multiplexer abstract view
.subckt multiplexer ay8913_do[0] ay8913_do[10] ay8913_do[11] ay8913_do[12] ay8913_do[13]
+ ay8913_do[14] ay8913_do[15] ay8913_do[16] ay8913_do[17] ay8913_do[18] ay8913_do[19]
+ ay8913_do[1] ay8913_do[20] ay8913_do[21] ay8913_do[22] ay8913_do[23] ay8913_do[24]
+ ay8913_do[25] ay8913_do[26] ay8913_do[27] ay8913_do[2] ay8913_do[3] ay8913_do[4]
+ ay8913_do[5] ay8913_do[6] ay8913_do[7] ay8913_do[8] ay8913_do[9] blinker_do[0] blinker_do[1]
+ blinker_do[2] custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[12]
+ custom_settings[13] custom_settings[14] custom_settings[15] custom_settings[16]
+ custom_settings[17] custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20]
+ custom_settings[21] custom_settings[22] custom_settings[23] custom_settings[24]
+ custom_settings[25] custom_settings[26] custom_settings[27] custom_settings[28]
+ custom_settings[29] custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3]
+ custom_settings[4] custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8]
+ custom_settings[9] diceroll_do[0] diceroll_do[1] diceroll_do[2] diceroll_do[3] diceroll_do[4]
+ diceroll_do[5] diceroll_do[6] diceroll_do[7] diceroll_do[8] hellorld_do io_in_0
+ io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16]
+ io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23]
+ io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30]
+ io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1] irq[2] mc14500_do[0] mc14500_do[10]
+ mc14500_do[11] mc14500_do[12] mc14500_do[13] mc14500_do[14] mc14500_do[15] mc14500_do[16]
+ mc14500_do[17] mc14500_do[18] mc14500_do[19] mc14500_do[1] mc14500_do[20] mc14500_do[21]
+ mc14500_do[22] mc14500_do[23] mc14500_do[24] mc14500_do[25] mc14500_do[26] mc14500_do[27]
+ mc14500_do[28] mc14500_do[29] mc14500_do[2] mc14500_do[30] mc14500_do[3] mc14500_do[4]
+ mc14500_do[5] mc14500_do[6] mc14500_do[7] mc14500_do[8] mc14500_do[9] mc14500_sram_addr[0]
+ mc14500_sram_addr[1] mc14500_sram_addr[2] mc14500_sram_addr[3] mc14500_sram_addr[4]
+ mc14500_sram_addr[5] mc14500_sram_gwe mc14500_sram_in[0] mc14500_sram_in[1] mc14500_sram_in[2]
+ mc14500_sram_in[3] mc14500_sram_in[4] mc14500_sram_in[5] mc14500_sram_in[6] mc14500_sram_in[7]
+ pdp11_do[0] pdp11_do[10] pdp11_do[11] pdp11_do[12] pdp11_do[13] pdp11_do[14] pdp11_do[15]
+ pdp11_do[16] pdp11_do[17] pdp11_do[18] pdp11_do[19] pdp11_do[1] pdp11_do[20] pdp11_do[21]
+ pdp11_do[22] pdp11_do[23] pdp11_do[24] pdp11_do[25] pdp11_do[26] pdp11_do[27] pdp11_do[28]
+ pdp11_do[29] pdp11_do[2] pdp11_do[30] pdp11_do[31] pdp11_do[32] pdp11_do[3] pdp11_do[4]
+ pdp11_do[5] pdp11_do[6] pdp11_do[7] pdp11_do[8] pdp11_do[9] pdp11_oeb[0] pdp11_oeb[10]
+ pdp11_oeb[11] pdp11_oeb[12] pdp11_oeb[13] pdp11_oeb[14] pdp11_oeb[15] pdp11_oeb[16]
+ pdp11_oeb[17] pdp11_oeb[18] pdp11_oeb[19] pdp11_oeb[1] pdp11_oeb[20] pdp11_oeb[21]
+ pdp11_oeb[22] pdp11_oeb[23] pdp11_oeb[24] pdp11_oeb[25] pdp11_oeb[26] pdp11_oeb[27]
+ pdp11_oeb[28] pdp11_oeb[29] pdp11_oeb[2] pdp11_oeb[30] pdp11_oeb[31] pdp11_oeb[32]
+ pdp11_oeb[3] pdp11_oeb[4] pdp11_oeb[5] pdp11_oeb[6] pdp11_oeb[7] pdp11_oeb[8] pdp11_oeb[9]
+ qcpu_do[0] qcpu_do[10] qcpu_do[11] qcpu_do[12] qcpu_do[13] qcpu_do[14] qcpu_do[15]
+ qcpu_do[16] qcpu_do[17] qcpu_do[18] qcpu_do[19] qcpu_do[1] qcpu_do[20] qcpu_do[21]
+ qcpu_do[22] qcpu_do[23] qcpu_do[24] qcpu_do[25] qcpu_do[26] qcpu_do[27] qcpu_do[28]
+ qcpu_do[29] qcpu_do[2] qcpu_do[30] qcpu_do[31] qcpu_do[32] qcpu_do[3] qcpu_do[4]
+ qcpu_do[5] qcpu_do[6] qcpu_do[7] qcpu_do[8] qcpu_do[9] qcpu_oeb[0] qcpu_oeb[10]
+ qcpu_oeb[11] qcpu_oeb[12] qcpu_oeb[13] qcpu_oeb[14] qcpu_oeb[15] qcpu_oeb[16] qcpu_oeb[17]
+ qcpu_oeb[18] qcpu_oeb[19] qcpu_oeb[1] qcpu_oeb[20] qcpu_oeb[21] qcpu_oeb[22] qcpu_oeb[23]
+ qcpu_oeb[24] qcpu_oeb[25] qcpu_oeb[26] qcpu_oeb[27] qcpu_oeb[28] qcpu_oeb[29] qcpu_oeb[2]
+ qcpu_oeb[30] qcpu_oeb[31] qcpu_oeb[32] qcpu_oeb[3] qcpu_oeb[4] qcpu_oeb[5] qcpu_oeb[6]
+ qcpu_oeb[7] qcpu_oeb[8] qcpu_oeb[9] qcpu_sram_addr[0] qcpu_sram_addr[1] qcpu_sram_addr[2]
+ qcpu_sram_addr[3] qcpu_sram_addr[4] qcpu_sram_addr[5] qcpu_sram_gwe qcpu_sram_in[0]
+ qcpu_sram_in[1] qcpu_sram_in[2] qcpu_sram_in[3] qcpu_sram_in[4] qcpu_sram_in[5]
+ qcpu_sram_in[6] qcpu_sram_in[7] qcpu_sram_out[0] qcpu_sram_out[1] qcpu_sram_out[2]
+ qcpu_sram_out[3] qcpu_sram_out[4] qcpu_sram_out[5] qcpu_sram_out[6] qcpu_sram_out[7]
+ rst_ay8913 rst_blinker rst_diceroll rst_hellorld rst_mc14500 rst_pdp11 rst_qcpu
+ rst_sid rst_sn76489 rst_tbb1143 rst_tholin_riscv rst_ue1 sid_do[0] sid_do[10] sid_do[11]
+ sid_do[12] sid_do[13] sid_do[14] sid_do[15] sid_do[16] sid_do[17] sid_do[18] sid_do[19]
+ sid_do[1] sid_do[20] sid_do[2] sid_do[3] sid_do[4] sid_do[5] sid_do[6] sid_do[7]
+ sid_do[8] sid_do[9] sid_oeb sn76489_do[0] sn76489_do[10] sn76489_do[11] sn76489_do[12]
+ sn76489_do[13] sn76489_do[14] sn76489_do[15] sn76489_do[16] sn76489_do[17] sn76489_do[18]
+ sn76489_do[19] sn76489_do[1] sn76489_do[20] sn76489_do[21] sn76489_do[22] sn76489_do[23]
+ sn76489_do[24] sn76489_do[25] sn76489_do[26] sn76489_do[27] sn76489_do[2] sn76489_do[3]
+ sn76489_do[4] sn76489_do[5] sn76489_do[6] sn76489_do[7] sn76489_do[8] sn76489_do[9]
+ tbb1143_do[0] tbb1143_do[1] tbb1143_do[2] tbb1143_do[3] tbb1143_do[4] tholin_riscv_do[0]
+ tholin_riscv_do[10] tholin_riscv_do[11] tholin_riscv_do[12] tholin_riscv_do[13]
+ tholin_riscv_do[14] tholin_riscv_do[15] tholin_riscv_do[16] tholin_riscv_do[17]
+ tholin_riscv_do[18] tholin_riscv_do[19] tholin_riscv_do[1] tholin_riscv_do[20] tholin_riscv_do[21]
+ tholin_riscv_do[22] tholin_riscv_do[23] tholin_riscv_do[24] tholin_riscv_do[25]
+ tholin_riscv_do[26] tholin_riscv_do[27] tholin_riscv_do[28] tholin_riscv_do[29]
+ tholin_riscv_do[2] tholin_riscv_do[30] tholin_riscv_do[31] tholin_riscv_do[32] tholin_riscv_do[3]
+ tholin_riscv_do[4] tholin_riscv_do[5] tholin_riscv_do[6] tholin_riscv_do[7] tholin_riscv_do[8]
+ tholin_riscv_do[9] tholin_riscv_oeb[0] tholin_riscv_oeb[10] tholin_riscv_oeb[11]
+ tholin_riscv_oeb[12] tholin_riscv_oeb[13] tholin_riscv_oeb[14] tholin_riscv_oeb[15]
+ tholin_riscv_oeb[16] tholin_riscv_oeb[17] tholin_riscv_oeb[18] tholin_riscv_oeb[19]
+ tholin_riscv_oeb[1] tholin_riscv_oeb[20] tholin_riscv_oeb[21] tholin_riscv_oeb[22]
+ tholin_riscv_oeb[23] tholin_riscv_oeb[24] tholin_riscv_oeb[25] tholin_riscv_oeb[26]
+ tholin_riscv_oeb[27] tholin_riscv_oeb[28] tholin_riscv_oeb[29] tholin_riscv_oeb[2]
+ tholin_riscv_oeb[30] tholin_riscv_oeb[31] tholin_riscv_oeb[32] tholin_riscv_oeb[3]
+ tholin_riscv_oeb[4] tholin_riscv_oeb[5] tholin_riscv_oeb[6] tholin_riscv_oeb[7]
+ tholin_riscv_oeb[8] tholin_riscv_oeb[9] ue1_do[0] ue1_do[1] ue1_do[2] ue1_do[3]
+ ue1_do[4] ue1_do[5] ue1_do[6] ue1_do[7] ue1_do[8] ue1_do[9] ue1_oeb vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i
+ wbs_we_i
.ends

* Black-box entry subcircuit for tholin_avalonsemi_tbb1143 abstract view
.subckt tholin_avalonsemi_tbb1143 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] rst_n vdd vss
.ends

* Black-box entry subcircuit for wrapped_tholin_riscv abstract view
.subckt wrapped_tholin_riscv custom_settings[0] custom_settings[1] io_in[0] io_in[10]
+ io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26]
+ io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[3] io_oeb[4]
+ io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11]
+ io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19]
+ io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26]
+ io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_qcpu abstract view
.subckt wrapped_qcpu custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[12]
+ custom_settings[13] custom_settings[14] custom_settings[15] custom_settings[16]
+ custom_settings[17] custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20]
+ custom_settings[21] custom_settings[22] custom_settings[23] custom_settings[24]
+ custom_settings[25] custom_settings[26] custom_settings[27] custom_settings[28]
+ custom_settings[29] custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3]
+ custom_settings[4] custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8]
+ custom_settings[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17]
+ io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24]
+ io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31]
+ io_oeb[32] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8]
+ io_out[9] rst_n sram_addr[0] sram_addr[1] sram_addr[2] sram_addr[3] sram_addr[4]
+ sram_addr[5] sram_gwe sram_in[0] sram_in[1] sram_in[2] sram_in[3] sram_in[4] sram_in[5]
+ sram_in[6] sram_in[7] sram_out[0] sram_out[1] sram_out[2] sram_out[3] sram_out[4]
+ sram_out[5] sram_out[6] sram_out[7] vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for diceroll abstract view
.subckt diceroll io_in io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] rst_n vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for ue1 abstract view
.subckt ue1 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb io_out[0] io_out[1]
+ io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ rst_n vdd vss
.ends

* Black-box entry subcircuit for hellorld abstract view
.subckt hellorld custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[1]
+ custom_settings[2] custom_settings[3] custom_settings[4] custom_settings[5] custom_settings[6]
+ custom_settings[7] custom_settings[8] custom_settings[9] io_out rst_n vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_sn76489 abstract view
.subckt wrapped_sn76489 custom_settings[0] custom_settings[1] io_in_1[0] io_in_1[1]
+ io_in_1[2] io_in_1[3] io_in_1[4] io_in_1[5] io_in_1[6] io_in_1[7] io_in_2 io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17]
+ io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24]
+ io_out[25] io_out[26] io_out[27] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_ay8913 abstract view
.subckt wrapped_ay8913 custom_settings[0] custom_settings[1] custom_settings[2] custom_settings[3]
+ io_in_1[0] io_in_1[1] io_in_1[2] io_in_1[3] io_in_1[4] io_in_1[5] io_in_1[6] io_in_1[7]
+ io_in_2[0] io_in_2[1] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[2] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xwrapped_pdp11 custom_settings\[0\] custom_settings\[10\] custom_settings\[11\] custom_settings\[12\]
+ custom_settings\[13\] custom_settings\[14\] custom_settings\[15\] custom_settings\[16\]
+ custom_settings\[17\] custom_settings\[18\] custom_settings\[19\] custom_settings\[1\]
+ custom_settings\[2\] custom_settings\[3\] custom_settings\[4\] custom_settings\[5\]
+ custom_settings\[6\] custom_settings\[7\] custom_settings\[8\] custom_settings\[9\]
+ io_in[5] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[6] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[7] io_in[35] io_in[36] io_in[37] io_in[8]
+ io_in[9] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] pdp11_oeb\[0\] pdp11_oeb\[10\]
+ pdp11_oeb\[11\] pdp11_oeb\[12\] pdp11_oeb\[13\] pdp11_oeb\[14\] pdp11_oeb\[15\]
+ pdp11_oeb\[16\] pdp11_oeb\[17\] pdp11_oeb\[18\] pdp11_oeb\[19\] pdp11_oeb\[1\] pdp11_oeb\[20\]
+ pdp11_oeb\[21\] pdp11_oeb\[22\] pdp11_oeb\[23\] pdp11_oeb\[24\] pdp11_oeb\[25\]
+ pdp11_oeb\[26\] pdp11_oeb\[27\] pdp11_oeb\[28\] pdp11_oeb\[29\] pdp11_oeb\[2\] pdp11_oeb\[30\]
+ pdp11_oeb\[31\] pdp11_oeb\[32\] pdp11_oeb\[3\] pdp11_oeb\[4\] pdp11_oeb\[5\] pdp11_oeb\[6\]
+ pdp11_oeb\[7\] pdp11_oeb\[8\] pdp11_oeb\[9\] pdp11_do\[0\] pdp11_do\[10\] pdp11_do\[11\]
+ pdp11_do\[12\] pdp11_do\[13\] pdp11_do\[14\] pdp11_do\[15\] pdp11_do\[16\] pdp11_do\[17\]
+ pdp11_do\[18\] pdp11_do\[19\] pdp11_do\[1\] pdp11_do\[20\] pdp11_do\[21\] pdp11_do\[22\]
+ pdp11_do\[23\] pdp11_do\[24\] pdp11_do\[25\] pdp11_do\[26\] pdp11_do\[27\] pdp11_do\[28\]
+ pdp11_do\[29\] pdp11_do\[2\] pdp11_do\[30\] pdp11_do\[31\] pdp11_do\[32\] pdp11_do\[3\]
+ pdp11_do\[4\] pdp11_do\[5\] pdp11_do\[6\] pdp11_do\[7\] pdp11_do\[8\] pdp11_do\[9\]
+ rst_pdp11 vdd vss wb_clk_i wrapped_pdp11
Xavali_logo vss vdd avali_logo
Xsid io_in[5] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[6] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[7] io_in[35] io_in[36] io_in[37]
+ io_in[8] io_in[9] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] sid_oeb sid_do\[0\]
+ sid_do\[10\] sid_do\[11\] sid_do\[12\] sid_do\[13\] sid_do\[14\] sid_do\[15\] sid_do\[16\]
+ sid_do\[17\] sid_do\[18\] sid_do\[19\] sid_do\[1\] sid_do\[20\] sid_do\[2\] sid_do\[3\]
+ sid_do\[4\] sid_do\[5\] sid_do\[6\] sid_do\[7\] sid_do\[8\] sid_do\[9\] rst_sid
+ vdd vss wb_clk_i wrapped_sid
Xmc14500 io_in[36] io_in[37] custom_settings\[0\] io_in[5] io_in[6] io_in[7] io_in[8]
+ io_in[9] io_in[10] io_in[11] io_in[12] mc14500_do\[0\] mc14500_do\[10\] mc14500_do\[11\]
+ mc14500_do\[12\] mc14500_do\[13\] mc14500_do\[14\] mc14500_do\[15\] mc14500_do\[16\]
+ mc14500_do\[17\] mc14500_do\[18\] mc14500_do\[19\] mc14500_do\[1\] mc14500_do\[20\]
+ mc14500_do\[21\] mc14500_do\[22\] mc14500_do\[23\] mc14500_do\[24\] mc14500_do\[25\]
+ mc14500_do\[26\] mc14500_do\[27\] mc14500_do\[28\] mc14500_do\[29\] mc14500_do\[2\]
+ mc14500_do\[30\] mc14500_do\[3\] mc14500_do\[4\] mc14500_do\[5\] mc14500_do\[6\]
+ mc14500_do\[7\] mc14500_do\[8\] mc14500_do\[9\] rst_mc14500 mc14500_sram_addr\[0\]
+ mc14500_sram_addr\[1\] mc14500_sram_addr\[2\] mc14500_sram_addr\[3\] mc14500_sram_addr\[4\]
+ mc14500_sram_addr\[5\] mc14500_sram_gwe mc14500_sram_in\[0\] mc14500_sram_in\[1\]
+ mc14500_sram_in\[2\] mc14500_sram_in\[3\] mc14500_sram_in\[4\] mc14500_sram_in\[5\]
+ mc14500_sram_in\[6\] mc14500_sram_in\[7\] qcpu_sram_out\[0\] qcpu_sram_out\[1\]
+ qcpu_sram_out\[2\] qcpu_sram_out\[3\] qcpu_sram_out\[4\] qcpu_sram_out\[5\] qcpu_sram_out\[6\]
+ qcpu_sram_out\[7\] vdd vss wrapped_mc14500
Xblinker blinker_do\[0\] blinker_do\[1\] blinker_do\[2\] rst_blinker vdd vss wb_clk_i
+ blinker
Xmultiplexer ay8913_do\[0\] ay8913_do\[10\] ay8913_do\[11\] ay8913_do\[12\] ay8913_do\[13\]
+ ay8913_do\[14\] ay8913_do\[15\] ay8913_do\[16\] ay8913_do\[17\] ay8913_do\[18\]
+ ay8913_do\[19\] ay8913_do\[1\] ay8913_do\[20\] ay8913_do\[21\] ay8913_do\[22\] ay8913_do\[23\]
+ ay8913_do\[24\] ay8913_do\[25\] ay8913_do\[26\] ay8913_do\[27\] ay8913_do\[2\] ay8913_do\[3\]
+ ay8913_do\[4\] ay8913_do\[5\] ay8913_do\[6\] ay8913_do\[7\] ay8913_do\[8\] ay8913_do\[9\]
+ blinker_do\[0\] blinker_do\[1\] blinker_do\[2\] custom_settings\[0\] custom_settings\[10\]
+ custom_settings\[11\] custom_settings\[12\] custom_settings\[13\] custom_settings\[14\]
+ custom_settings\[15\] custom_settings\[16\] custom_settings\[17\] custom_settings\[18\]
+ custom_settings\[19\] custom_settings\[1\] custom_settings\[20\] custom_settings\[21\]
+ custom_settings\[22\] custom_settings\[23\] custom_settings\[24\] custom_settings\[25\]
+ custom_settings\[26\] custom_settings\[27\] custom_settings\[28\] custom_settings\[29\]
+ custom_settings\[2\] custom_settings\[30\] custom_settings\[31\] custom_settings\[3\]
+ custom_settings\[4\] custom_settings\[5\] custom_settings\[6\] custom_settings\[7\]
+ custom_settings\[8\] custom_settings\[9\] diceroll_do\[0\] diceroll_do\[1\] diceroll_do\[2\]
+ diceroll_do\[3\] diceroll_do\[4\] diceroll_do\[5\] diceroll_do\[6\] diceroll_do\[7\]
+ diceroll_do\[8\] hellorld_do io_in[0] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ user_irq[0] user_irq[1] user_irq[2] mc14500_do\[0\] mc14500_do\[10\] mc14500_do\[11\]
+ mc14500_do\[12\] mc14500_do\[13\] mc14500_do\[14\] mc14500_do\[15\] mc14500_do\[16\]
+ mc14500_do\[17\] mc14500_do\[18\] mc14500_do\[19\] mc14500_do\[1\] mc14500_do\[20\]
+ mc14500_do\[21\] mc14500_do\[22\] mc14500_do\[23\] mc14500_do\[24\] mc14500_do\[25\]
+ mc14500_do\[26\] mc14500_do\[27\] mc14500_do\[28\] mc14500_do\[29\] mc14500_do\[2\]
+ mc14500_do\[30\] mc14500_do\[3\] mc14500_do\[4\] mc14500_do\[5\] mc14500_do\[6\]
+ mc14500_do\[7\] mc14500_do\[8\] mc14500_do\[9\] mc14500_sram_addr\[0\] mc14500_sram_addr\[1\]
+ mc14500_sram_addr\[2\] mc14500_sram_addr\[3\] mc14500_sram_addr\[4\] mc14500_sram_addr\[5\]
+ mc14500_sram_gwe mc14500_sram_in\[0\] mc14500_sram_in\[1\] mc14500_sram_in\[2\]
+ mc14500_sram_in\[3\] mc14500_sram_in\[4\] mc14500_sram_in\[5\] mc14500_sram_in\[6\]
+ mc14500_sram_in\[7\] pdp11_do\[0\] pdp11_do\[10\] pdp11_do\[11\] pdp11_do\[12\]
+ pdp11_do\[13\] pdp11_do\[14\] pdp11_do\[15\] pdp11_do\[16\] pdp11_do\[17\] pdp11_do\[18\]
+ pdp11_do\[19\] pdp11_do\[1\] pdp11_do\[20\] pdp11_do\[21\] pdp11_do\[22\] pdp11_do\[23\]
+ pdp11_do\[24\] pdp11_do\[25\] pdp11_do\[26\] pdp11_do\[27\] pdp11_do\[28\] pdp11_do\[29\]
+ pdp11_do\[2\] pdp11_do\[30\] pdp11_do\[31\] pdp11_do\[32\] pdp11_do\[3\] pdp11_do\[4\]
+ pdp11_do\[5\] pdp11_do\[6\] pdp11_do\[7\] pdp11_do\[8\] pdp11_do\[9\] pdp11_oeb\[0\]
+ pdp11_oeb\[10\] pdp11_oeb\[11\] pdp11_oeb\[12\] pdp11_oeb\[13\] pdp11_oeb\[14\]
+ pdp11_oeb\[15\] pdp11_oeb\[16\] pdp11_oeb\[17\] pdp11_oeb\[18\] pdp11_oeb\[19\]
+ pdp11_oeb\[1\] pdp11_oeb\[20\] pdp11_oeb\[21\] pdp11_oeb\[22\] pdp11_oeb\[23\] pdp11_oeb\[24\]
+ pdp11_oeb\[25\] pdp11_oeb\[26\] pdp11_oeb\[27\] pdp11_oeb\[28\] pdp11_oeb\[29\]
+ pdp11_oeb\[2\] pdp11_oeb\[30\] pdp11_oeb\[31\] pdp11_oeb\[32\] pdp11_oeb\[3\] pdp11_oeb\[4\]
+ pdp11_oeb\[5\] pdp11_oeb\[6\] pdp11_oeb\[7\] pdp11_oeb\[8\] pdp11_oeb\[9\] qcpu_do\[0\]
+ qcpu_do\[10\] qcpu_do\[11\] qcpu_do\[12\] qcpu_do\[13\] qcpu_do\[14\] qcpu_do\[15\]
+ qcpu_do\[16\] qcpu_do\[17\] qcpu_do\[18\] qcpu_do\[19\] qcpu_do\[1\] qcpu_do\[20\]
+ qcpu_do\[21\] qcpu_do\[22\] qcpu_do\[23\] qcpu_do\[24\] qcpu_do\[25\] qcpu_do\[26\]
+ qcpu_do\[27\] qcpu_do\[28\] qcpu_do\[29\] qcpu_do\[2\] qcpu_do\[30\] qcpu_do\[31\]
+ qcpu_do\[32\] qcpu_do\[3\] qcpu_do\[4\] qcpu_do\[5\] qcpu_do\[6\] qcpu_do\[7\] qcpu_do\[8\]
+ qcpu_do\[9\] qcpu_oeb\[0\] qcpu_oeb\[10\] qcpu_oeb\[11\] qcpu_oeb\[12\] qcpu_oeb\[13\]
+ qcpu_oeb\[14\] qcpu_oeb\[15\] qcpu_oeb\[16\] qcpu_oeb\[17\] qcpu_oeb\[18\] qcpu_oeb\[19\]
+ qcpu_oeb\[1\] qcpu_oeb\[20\] qcpu_oeb\[21\] qcpu_oeb\[22\] qcpu_oeb\[23\] qcpu_oeb\[24\]
+ qcpu_oeb\[25\] qcpu_oeb\[26\] qcpu_oeb\[27\] qcpu_oeb\[28\] qcpu_oeb\[29\] qcpu_oeb\[2\]
+ qcpu_oeb\[30\] qcpu_oeb\[31\] qcpu_oeb\[32\] qcpu_oeb\[3\] qcpu_oeb\[4\] qcpu_oeb\[5\]
+ qcpu_oeb\[6\] qcpu_oeb\[7\] qcpu_oeb\[8\] qcpu_oeb\[9\] qcpu_sram_addr\[0\] qcpu_sram_addr\[1\]
+ qcpu_sram_addr\[2\] qcpu_sram_addr\[3\] qcpu_sram_addr\[4\] qcpu_sram_addr\[5\]
+ qcpu_sram_gwe qcpu_sram_in\[0\] qcpu_sram_in\[1\] qcpu_sram_in\[2\] qcpu_sram_in\[3\]
+ qcpu_sram_in\[4\] qcpu_sram_in\[5\] qcpu_sram_in\[6\] qcpu_sram_in\[7\] qcpu_sram_out\[0\]
+ qcpu_sram_out\[1\] qcpu_sram_out\[2\] qcpu_sram_out\[3\] qcpu_sram_out\[4\] qcpu_sram_out\[5\]
+ qcpu_sram_out\[6\] qcpu_sram_out\[7\] rst_ay8913 rst_blinker rst_diceroll rst_hellorld
+ rst_mc14500 rst_pdp11 rst_qcpu rst_sid rst_sn76489 rst_tbb1143 rst_tholin_riscv
+ rst_ue1 sid_do\[0\] sid_do\[10\] sid_do\[11\] sid_do\[12\] sid_do\[13\] sid_do\[14\]
+ sid_do\[15\] sid_do\[16\] sid_do\[17\] sid_do\[18\] sid_do\[19\] sid_do\[1\] sid_do\[20\]
+ sid_do\[2\] sid_do\[3\] sid_do\[4\] sid_do\[5\] sid_do\[6\] sid_do\[7\] sid_do\[8\]
+ sid_do\[9\] sid_oeb sn76489_do\[0\] sn76489_do\[10\] sn76489_do\[11\] sn76489_do\[12\]
+ sn76489_do\[13\] sn76489_do\[14\] sn76489_do\[15\] sn76489_do\[16\] sn76489_do\[17\]
+ sn76489_do\[18\] sn76489_do\[19\] sn76489_do\[1\] sn76489_do\[20\] sn76489_do\[21\]
+ sn76489_do\[22\] sn76489_do\[23\] sn76489_do\[24\] sn76489_do\[25\] sn76489_do\[26\]
+ sn76489_do\[27\] sn76489_do\[2\] sn76489_do\[3\] sn76489_do\[4\] sn76489_do\[5\]
+ sn76489_do\[6\] sn76489_do\[7\] sn76489_do\[8\] sn76489_do\[9\] tbb1143_do\[0\]
+ tbb1143_do\[1\] tbb1143_do\[2\] tbb1143_do\[3\] tbb1143_do\[4\] tholin_riscv_do\[0\]
+ tholin_riscv_do\[10\] tholin_riscv_do\[11\] tholin_riscv_do\[12\] tholin_riscv_do\[13\]
+ tholin_riscv_do\[14\] tholin_riscv_do\[15\] tholin_riscv_do\[16\] tholin_riscv_do\[17\]
+ tholin_riscv_do\[18\] tholin_riscv_do\[19\] tholin_riscv_do\[1\] tholin_riscv_do\[20\]
+ tholin_riscv_do\[21\] tholin_riscv_do\[22\] tholin_riscv_do\[23\] tholin_riscv_do\[24\]
+ tholin_riscv_do\[25\] tholin_riscv_do\[26\] tholin_riscv_do\[27\] tholin_riscv_do\[28\]
+ tholin_riscv_do\[29\] tholin_riscv_do\[2\] tholin_riscv_do\[30\] tholin_riscv_do\[31\]
+ tholin_riscv_do\[32\] tholin_riscv_do\[3\] tholin_riscv_do\[4\] tholin_riscv_do\[5\]
+ tholin_riscv_do\[6\] tholin_riscv_do\[7\] tholin_riscv_do\[8\] tholin_riscv_do\[9\]
+ tholin_riscv_oeb\[0\] tholin_riscv_oeb\[10\] tholin_riscv_oeb\[11\] tholin_riscv_oeb\[12\]
+ tholin_riscv_oeb\[13\] tholin_riscv_oeb\[14\] tholin_riscv_oeb\[15\] tholin_riscv_oeb\[16\]
+ tholin_riscv_oeb\[17\] tholin_riscv_oeb\[18\] tholin_riscv_oeb\[19\] tholin_riscv_oeb\[1\]
+ tholin_riscv_oeb\[20\] tholin_riscv_oeb\[21\] tholin_riscv_oeb\[22\] tholin_riscv_oeb\[23\]
+ tholin_riscv_oeb\[24\] tholin_riscv_oeb\[25\] tholin_riscv_oeb\[26\] tholin_riscv_oeb\[27\]
+ tholin_riscv_oeb\[28\] tholin_riscv_oeb\[29\] tholin_riscv_oeb\[2\] tholin_riscv_oeb\[30\]
+ tholin_riscv_oeb\[31\] tholin_riscv_oeb\[32\] tholin_riscv_oeb\[3\] tholin_riscv_oeb\[4\]
+ tholin_riscv_oeb\[5\] tholin_riscv_oeb\[6\] tholin_riscv_oeb\[7\] tholin_riscv_oeb\[8\]
+ tholin_riscv_oeb\[9\] ue1_do\[0\] ue1_do\[1\] ue1_do\[2\] ue1_do\[3\] ue1_do\[4\]
+ ue1_do\[5\] ue1_do\[6\] ue1_do\[7\] ue1_do\[8\] ue1_do\[9\] ue1_oeb vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i
+ wbs_we_i multiplexer
Xtbb1143 io_in[11] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in[10] tbb1143_do\[0\]
+ tbb1143_do\[1\] tbb1143_do\[2\] tbb1143_do\[3\] tbb1143_do\[4\] rst_tbb1143 vdd
+ vss tholin_avalonsemi_tbb1143
Xwrapped_tholin_riscv custom_settings\[0\] custom_settings\[1\] io_in[5] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[6] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[7] io_in[35] io_in[36] io_in[37] io_in[8] io_in[9]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] tholin_riscv_oeb\[0\] tholin_riscv_oeb\[10\]
+ tholin_riscv_oeb\[11\] tholin_riscv_oeb\[12\] tholin_riscv_oeb\[13\] tholin_riscv_oeb\[14\]
+ tholin_riscv_oeb\[15\] tholin_riscv_oeb\[16\] tholin_riscv_oeb\[17\] tholin_riscv_oeb\[18\]
+ tholin_riscv_oeb\[19\] tholin_riscv_oeb\[1\] tholin_riscv_oeb\[20\] tholin_riscv_oeb\[21\]
+ tholin_riscv_oeb\[22\] tholin_riscv_oeb\[23\] tholin_riscv_oeb\[24\] tholin_riscv_oeb\[25\]
+ tholin_riscv_oeb\[26\] tholin_riscv_oeb\[27\] tholin_riscv_oeb\[28\] tholin_riscv_oeb\[29\]
+ tholin_riscv_oeb\[2\] tholin_riscv_oeb\[30\] tholin_riscv_oeb\[31\] tholin_riscv_oeb\[32\]
+ tholin_riscv_oeb\[3\] tholin_riscv_oeb\[4\] tholin_riscv_oeb\[5\] tholin_riscv_oeb\[6\]
+ tholin_riscv_oeb\[7\] tholin_riscv_oeb\[8\] tholin_riscv_oeb\[9\] tholin_riscv_do\[0\]
+ tholin_riscv_do\[10\] tholin_riscv_do\[11\] tholin_riscv_do\[12\] tholin_riscv_do\[13\]
+ tholin_riscv_do\[14\] tholin_riscv_do\[15\] tholin_riscv_do\[16\] tholin_riscv_do\[17\]
+ tholin_riscv_do\[18\] tholin_riscv_do\[19\] tholin_riscv_do\[1\] tholin_riscv_do\[20\]
+ tholin_riscv_do\[21\] tholin_riscv_do\[22\] tholin_riscv_do\[23\] tholin_riscv_do\[24\]
+ tholin_riscv_do\[25\] tholin_riscv_do\[26\] tholin_riscv_do\[27\] tholin_riscv_do\[28\]
+ tholin_riscv_do\[29\] tholin_riscv_do\[2\] tholin_riscv_do\[30\] tholin_riscv_do\[31\]
+ tholin_riscv_do\[32\] tholin_riscv_do\[3\] tholin_riscv_do\[4\] tholin_riscv_do\[5\]
+ tholin_riscv_do\[6\] tholin_riscv_do\[7\] tholin_riscv_do\[8\] tholin_riscv_do\[9\]
+ rst_tholin_riscv vdd vss wb_clk_i wrapped_tholin_riscv
Xwrapped_qcpu custom_settings\[0\] custom_settings\[10\] custom_settings\[11\] custom_settings\[12\]
+ custom_settings\[13\] custom_settings\[14\] custom_settings\[15\] custom_settings\[16\]
+ custom_settings\[17\] custom_settings\[18\] custom_settings\[19\] custom_settings\[1\]
+ custom_settings\[20\] custom_settings\[21\] custom_settings\[22\] custom_settings\[23\]
+ custom_settings\[24\] custom_settings\[25\] custom_settings\[26\] custom_settings\[27\]
+ custom_settings\[28\] custom_settings\[29\] custom_settings\[2\] custom_settings\[30\]
+ custom_settings\[31\] custom_settings\[3\] custom_settings\[4\] custom_settings\[5\]
+ custom_settings\[6\] custom_settings\[7\] custom_settings\[8\] custom_settings\[9\]
+ io_in[5] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[6] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[7] io_in[35] io_in[36] io_in[37] io_in[8]
+ io_in[9] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] qcpu_oeb\[0\] qcpu_oeb\[10\]
+ qcpu_oeb\[11\] qcpu_oeb\[12\] qcpu_oeb\[13\] qcpu_oeb\[14\] qcpu_oeb\[15\] qcpu_oeb\[16\]
+ qcpu_oeb\[17\] qcpu_oeb\[18\] qcpu_oeb\[19\] qcpu_oeb\[1\] qcpu_oeb\[20\] qcpu_oeb\[21\]
+ qcpu_oeb\[22\] qcpu_oeb\[23\] qcpu_oeb\[24\] qcpu_oeb\[25\] qcpu_oeb\[26\] qcpu_oeb\[27\]
+ qcpu_oeb\[28\] qcpu_oeb\[29\] qcpu_oeb\[2\] qcpu_oeb\[30\] qcpu_oeb\[31\] qcpu_oeb\[32\]
+ qcpu_oeb\[3\] qcpu_oeb\[4\] qcpu_oeb\[5\] qcpu_oeb\[6\] qcpu_oeb\[7\] qcpu_oeb\[8\]
+ qcpu_oeb\[9\] qcpu_do\[0\] qcpu_do\[10\] qcpu_do\[11\] qcpu_do\[12\] qcpu_do\[13\]
+ qcpu_do\[14\] qcpu_do\[15\] qcpu_do\[16\] qcpu_do\[17\] qcpu_do\[18\] qcpu_do\[19\]
+ qcpu_do\[1\] qcpu_do\[20\] qcpu_do\[21\] qcpu_do\[22\] qcpu_do\[23\] qcpu_do\[24\]
+ qcpu_do\[25\] qcpu_do\[26\] qcpu_do\[27\] qcpu_do\[28\] qcpu_do\[29\] qcpu_do\[2\]
+ qcpu_do\[30\] qcpu_do\[31\] qcpu_do\[32\] qcpu_do\[3\] qcpu_do\[4\] qcpu_do\[5\]
+ qcpu_do\[6\] qcpu_do\[7\] qcpu_do\[8\] qcpu_do\[9\] rst_qcpu qcpu_sram_addr\[0\]
+ qcpu_sram_addr\[1\] qcpu_sram_addr\[2\] qcpu_sram_addr\[3\] qcpu_sram_addr\[4\]
+ qcpu_sram_addr\[5\] qcpu_sram_gwe qcpu_sram_in\[0\] qcpu_sram_in\[1\] qcpu_sram_in\[2\]
+ qcpu_sram_in\[3\] qcpu_sram_in\[4\] qcpu_sram_in\[5\] qcpu_sram_in\[6\] qcpu_sram_in\[7\]
+ qcpu_sram_out\[0\] qcpu_sram_out\[1\] qcpu_sram_out\[2\] qcpu_sram_out\[3\] qcpu_sram_out\[4\]
+ qcpu_sram_out\[5\] qcpu_sram_out\[6\] qcpu_sram_out\[7\] vdd vss wb_clk_i wrapped_qcpu
Xdiceroll io_in[5] diceroll_do\[0\] diceroll_do\[1\] diceroll_do\[2\] diceroll_do\[3\]
+ diceroll_do\[4\] diceroll_do\[5\] diceroll_do\[6\] diceroll_do\[7\] diceroll_do\[8\]
+ rst_diceroll vdd vss wb_clk_i diceroll
Xue1 io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in[10] ue1_oeb ue1_do\[0\] ue1_do\[1\]
+ ue1_do\[2\] ue1_do\[3\] ue1_do\[4\] ue1_do\[5\] ue1_do\[6\] ue1_do\[7\] ue1_do\[8\]
+ ue1_do\[9\] rst_ue1 vdd vss ue1
Xhellorld custom_settings\[0\] custom_settings\[10\] custom_settings\[11\] custom_settings\[1\]
+ custom_settings\[2\] custom_settings\[3\] custom_settings\[4\] custom_settings\[5\]
+ custom_settings\[6\] custom_settings\[7\] custom_settings\[8\] custom_settings\[9\]
+ hellorld_do rst_hellorld vdd vss wb_clk_i hellorld
Xwrapped_sn76489 custom_settings\[0\] custom_settings\[1\] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_in[10] io_in[11] io_in[12] io_in[19] sn76489_do\[0\] sn76489_do\[10\]
+ sn76489_do\[11\] sn76489_do\[12\] sn76489_do\[13\] sn76489_do\[14\] sn76489_do\[15\]
+ sn76489_do\[16\] sn76489_do\[17\] sn76489_do\[18\] sn76489_do\[19\] sn76489_do\[1\]
+ sn76489_do\[20\] sn76489_do\[21\] sn76489_do\[22\] sn76489_do\[23\] sn76489_do\[24\]
+ sn76489_do\[25\] sn76489_do\[26\] sn76489_do\[27\] sn76489_do\[2\] sn76489_do\[3\]
+ sn76489_do\[4\] sn76489_do\[5\] sn76489_do\[6\] sn76489_do\[7\] sn76489_do\[8\]
+ sn76489_do\[9\] rst_sn76489 vdd vss wb_clk_i wrapped_sn76489
Xay8913 custom_settings\[0\] custom_settings\[1\] custom_settings\[2\] custom_settings\[3\]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in[10] io_in[11] io_in[12] io_in[19]
+ io_in[20] ay8913_do\[0\] ay8913_do\[10\] ay8913_do\[11\] ay8913_do\[12\] ay8913_do\[13\]
+ ay8913_do\[14\] ay8913_do\[15\] ay8913_do\[16\] ay8913_do\[17\] ay8913_do\[18\]
+ ay8913_do\[19\] ay8913_do\[1\] ay8913_do\[20\] ay8913_do\[21\] ay8913_do\[22\] ay8913_do\[23\]
+ ay8913_do\[24\] ay8913_do\[25\] ay8913_do\[26\] ay8913_do\[27\] ay8913_do\[2\] ay8913_do\[3\]
+ ay8913_do\[4\] ay8913_do\[5\] ay8913_do\[6\] ay8913_do\[7\] ay8913_do\[8\] ay8913_do\[9\]
+ rst_ay8913 vdd vss wb_clk_i wrapped_ay8913
.ends

