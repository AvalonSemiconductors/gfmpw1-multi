module wrapped_sn76489 (io_in_2,
    rst_n,
    vdd,
    vss,
    wb_clk_i,
    custom_settings,
    io_in_1,
    io_out);
 input io_in_2;
 input rst_n;
 inout vdd;
 inout vss;
 input wb_clk_i;
 input [1:0] custom_settings;
 input [7:0] io_in_1;
 output [27:0] io_out;

 wire net28;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \tt_um_rejunity_sn76489.DAC_clk ;
 wire \tt_um_rejunity_sn76489.DAC_dat ;
 wire \tt_um_rejunity_sn76489.DAC_le ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.in ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.in ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.in ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.in ;
 wire \tt_um_rejunity_sn76489.clk_counter[0] ;
 wire \tt_um_rejunity_sn76489.clk_counter[1] ;
 wire \tt_um_rejunity_sn76489.clk_counter[2] ;
 wire \tt_um_rejunity_sn76489.clk_counter[3] ;
 wire \tt_um_rejunity_sn76489.clk_counter[4] ;
 wire \tt_um_rejunity_sn76489.clk_counter[5] ;
 wire \tt_um_rejunity_sn76489.clk_counter[6] ;
 wire \tt_um_rejunity_sn76489.control_noise[0][0] ;
 wire \tt_um_rejunity_sn76489.control_noise[0][1] ;
 wire \tt_um_rejunity_sn76489.control_noise[0][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][0] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][1] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][3] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][4] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][5] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][6] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][7] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][8] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][9] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][0] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][1] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][3] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][4] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][5] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][6] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][7] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][8] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][9] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][0] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][1] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][3] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][4] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][5] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][6] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][7] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][8] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][9] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[0] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[10] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[1] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[2] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[3] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[4] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[5] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[6] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[7] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[8] ;
 wire \tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[9] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[0] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[10] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[1] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[2] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[3] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[4] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[5] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[6] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[7] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[8] ;
 wire \tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[9] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[0] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[10] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[1] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[2] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[3] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[4] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[5] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[6] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[7] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[8] ;
 wire \tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[9] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[0] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[10] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[1] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[2] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[3] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[4] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[5] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[6] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[7] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[8] ;
 wire \tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[9] ;
 wire \tt_um_rejunity_sn76489.latch_control_reg[0] ;
 wire \tt_um_rejunity_sn76489.latch_control_reg[1] ;
 wire \tt_um_rejunity_sn76489.latch_control_reg[2] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.restart_noise ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[0] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[10] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[11] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[12] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[1] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[2] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[3] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[4] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[5] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[6] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[7] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[8] ;
 wire \tt_um_rejunity_sn76489.pwm.accumulator[9] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.counter[0] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.counter[1] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.counter[2] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.counter[3] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.counter[4] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[0] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[10] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[11] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[1] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[2] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[3] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[4] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[5] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[6] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[7] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[8] ;
 wire \tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[9] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[7] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[8] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[9] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[7] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[8] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[9] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[7] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[8] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[9] ;

 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1465__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\tt_um_rejunity_sn76489.chan[3].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1466__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0915_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1470__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\tt_um_rejunity_sn76489.chan[3].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1474__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0915_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1477__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\tt_um_rejunity_sn76489.chan[3].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1479__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0915_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1564__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\tt_um_rejunity_sn76489.chan[3].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1603__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1050_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1618__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1059_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1618__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1067_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1619__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1050_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1689__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1133_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1689__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1136_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1690__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1133_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1690__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1136_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1714__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1159_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1715__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1159_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1740__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1184_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1758__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1201_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1758__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1202_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1759__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1184_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1771__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1201_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1772__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1202_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1780__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net11));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1781__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1222_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1782__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1223_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1787__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1224_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1789__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net11));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1805__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net8));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1806__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net9));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1807__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net10));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1810__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net7));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1811__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net6));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1815__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1817__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net11));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1820__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1252_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1820__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1256_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1824__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net3));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1834__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net4));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1839__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net5));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1844__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net6));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1848__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1252_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1848__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1256_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1862__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net8));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1865__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1866__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1294_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1866__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1256_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1881__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1305_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1884__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1306_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1891__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1314_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1899__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1321_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1900__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1322_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1907__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1322_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1913__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1322_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1919__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1222_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1920__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1339_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1922__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1340_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1927__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1321_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1928__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1346_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1932__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1349_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1938__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1351_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1945__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1351_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1952__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1346_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1956__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1223_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1961__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1314_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1965__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1340_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1972__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1351_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1978__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1346_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1986__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1346_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1994__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1401_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__1997__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1133_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2000__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1321_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2001__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1408_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2004__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1159_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2005__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1133_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2008__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1351_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2012__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1184_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2013__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1159_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2017__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1416_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2022__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1184_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2024__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1408_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2028__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1416_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2032__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1416_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2036__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1408_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2042__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1408_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2049__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0195_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2050__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0196_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2057__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0196_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2064__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1401_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2067__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1136_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2070__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0196_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2074__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1136_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2077__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1416_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2086__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0221_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2093__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0196_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2097__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0221_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2100__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1306_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2109__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0246_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2111__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0915_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2112__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0246_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2186__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net1));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2187__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net1));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2189__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0311_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2192__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0314_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2193__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0315_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2195__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0221_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2199__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0221_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2204__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0322_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2208__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0322_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2212__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0322_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2216__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1223_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2220__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1224_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2222__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1059_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2223__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1222_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2224__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1059_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2230__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0195_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2259__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1401_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2265__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0195_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2274__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0322_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2303__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0195_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2304__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0315_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2304__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0408_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2308__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0411_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2315__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0418_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2316__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0417_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2317__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0412_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2322__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0418_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2324__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0412_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2325__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0314_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2333__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0434_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2350__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1401_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2362__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1339_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2374__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0314_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2377__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0470_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2379__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0411_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2379__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0474_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2393__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0315_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2393__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0408_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2401__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0434_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2423__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1339_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2425__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0513_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2437__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0434_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2439__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0513_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2440__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0521_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2446__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0513_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2447__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0521_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2456__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0470_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2457__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0474_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2461__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0543_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2462__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0544_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2463__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0543_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2472__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0315_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2472__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0408_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2479__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0513_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2480__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0521_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2485__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1339_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2488__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0521_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2489__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0411_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2495__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0434_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2509__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0418_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2510__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0544_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2511__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0412_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2522__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1340_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2528__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0314_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2529__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1340_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2530__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0470_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2533__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0418_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2534__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0544_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2535__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0412_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2536__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0470_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2537__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0411_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2537__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0474_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2539__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1305_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2540__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1059_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2541__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1067_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2550__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0408_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2561__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1349_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2592__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1349_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2609__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0672_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2610__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net23));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2611__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net23));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2614__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0474_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2620__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0681_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2623__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net25));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2630__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net25));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2631__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1224_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2632__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0691_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2635__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1224_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2637__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\tt_um_rejunity_sn76489.DAC_dat ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2642__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1222_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2668__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1223_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2688__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net23));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2689__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0417_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2693__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0417_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2694__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0739_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2695__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net25));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2698__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1306_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2698__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0246_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2701__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net10));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2705__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net9));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2709__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1294_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2730__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net7));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2736__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net9));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2738__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net10));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2746__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0782_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2747__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1305_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2750__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1305_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2753__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1349_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2760__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0782_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2763__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0782_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2789__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net8));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2795__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1294_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2798__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net3));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2802__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net4));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2806__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net5));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2810__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net8));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2812__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net10));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2816__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0681_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2817__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1252_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2819__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0681_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2822__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0681_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2829__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net6));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2835__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1294_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2850__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net9));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2852__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1252_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2860__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1256_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2863__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1306_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2865__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0544_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2877__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1322_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2885__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0417_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2891__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1314_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2895__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1314_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2897__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net4));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2897__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_1321_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2900__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2901__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2902__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2903__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2904__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2905__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2906__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2907__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2908__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2909__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2910__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2911__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2912__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2914__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2918__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2919__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2920__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2921__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2922__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2926__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2928__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2929__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2930__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2931__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2932__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2933__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2934__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2935__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2936__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2937__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2938__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2939__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2940__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2941__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2942__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2943__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2944__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2945__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2946__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2950__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2951__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2954__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2955__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2956__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2957__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2958__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2959__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2960__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2961__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2962__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2963__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2964__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2965__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2967__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2968__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2970__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2973__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2974__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2975__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2976__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2977__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2978__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2988__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2989__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2990__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2991__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2992__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2993__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2995__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2996__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2997__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2998__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__2999__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3000__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3001__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3002__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3003__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3004__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3006__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3007__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3008__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3009__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3010__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3011__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3012__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3013__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3014__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3015__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3017__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3018__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3019__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3020__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3021__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3022__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3023__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3024__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3025__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3026__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3027__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3028__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3029__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3029__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0129_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3030__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3031__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3032__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3033__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3034__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3035__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3036__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3037__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3038__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3039__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3040__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3041__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3042__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3042__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_0142_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3043__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3044__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3046__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3049__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3050__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3052__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3053__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3054__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3055__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3056__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3057__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3058__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3059__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3060__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3061__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3062__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3063__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3064__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3065__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3066__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3067__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3069__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3071__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3079__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3083__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3084__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3085__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3086__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3087__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3088__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3089__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3109__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\tt_um_rejunity_sn76489.pwm.accumulator[12] ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__3110__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\tt_um_rejunity_sn76489.DAC_dat ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_0_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_10_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_11_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_12_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_13_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_14_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_15_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_1_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_2_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_3_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_4_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_5_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_6_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_7_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_8_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_4_9_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload11_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload12_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload13_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload14_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload1_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload2_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload3_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload4_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload5_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload7_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload9_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input10_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_2));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input11_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(rst_n));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input1_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input2_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(custom_settings[1]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input3_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[1]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input4_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[2]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input5_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[3]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input6_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[4]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input7_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[5]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input8_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[6]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input9_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in_1[7]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_output23_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net23));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_output25_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net25));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_0_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_0_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_0_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_0_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_35 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_24_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_25_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_27_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_27_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_28_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_2_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_30_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_30_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_32_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_32_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_32_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_355 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_40_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_41_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_45_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_46_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_46_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_47_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_47_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_48_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_355 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_48_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_50_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_50_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_50_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_50_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_51_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_51_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_52_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_52_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_52_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_53_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_53_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_53_9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_54_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_54_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_54_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_54_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_54_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Left_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Left_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Left_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Left_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Left_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Left_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Left_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Left_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Left_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Left_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Left_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Left_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Left_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Left_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_22_Left_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_23_Left_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_24_Left_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_25_Left_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_26_Left_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_27_Left_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_28_Left_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_29_Left_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Left_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_30_Left_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_31_Left_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_32_Left_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_33_Left_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_34_Left_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_35_Left_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_36_Left_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_37_Left_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_38_Left_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_39_Left_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Left_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_40_Left_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_41_Left_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_42_Left_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_43_Left_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_44_Left_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_45_Left_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_45_Right_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_46_Left_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_46_Right_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_47_Left_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_47_Right_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_48_Left_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_48_Right_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_49_Left_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_49_Right_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Left_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_50_Left_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_50_Right_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_51_Left_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_51_Right_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_52_Left_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_52_Right_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_53_Left_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_53_Right_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_54_Left_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_54_Right_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Left_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Left_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Left_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Left_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Left_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_50_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_51_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_52_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_53_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_54_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1446_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ),
    .Y(_0896_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1447_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0897_),
    .B(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1448_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0897_),
    .Y(_0898_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1449_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.in ),
    .Y(_0899_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1450_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0900_),
    .B(_0899_),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1451_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0901_),
    .C(_0900_),
    .B(_0898_),
    .A(_0896_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1452_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0901_),
    .Y(_0902_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1453_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ),
    .Y(_0903_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1454_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.in ),
    .Y(_0904_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1455_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0905_),
    .B(_0904_),
    .A(_0903_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1456_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0905_),
    .Y(_0906_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1457_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0907_),
    .B(_0899_),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1458_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0908_),
    .B(_0899_),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1459_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0909_),
    .B(_0908_),
    .A(_0907_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1460_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0910_),
    .B(_0909_),
    .A(_0906_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1461_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0911_),
    .B(_0908_),
    .A(_0905_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1462_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0912_),
    .B(_0911_),
    .A(_0907_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1463_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ),
    .Y(_0913_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1464_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0902_),
    .B(_0910_),
    .C(_0912_),
    .D(_0913_),
    .Y(_0914_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1465_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.in ),
    .Y(_0915_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1466_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0916_),
    .B(_0915_),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1467_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0916_),
    .Y(_0917_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1468_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0917_),
    .Y(_0918_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1469_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .Y(_0919_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1470_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0920_),
    .B(\tt_um_rejunity_sn76489.chan[3].attenuation.in ),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1471_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0920_),
    .Y(_0921_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1472_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0922_),
    .B(_0921_),
    .A(_0919_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1473_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0923_),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1474_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0924_),
    .B(_0915_),
    .A(_0923_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1475_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0924_),
    .A(_0922_),
    .Y(_0925_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1476_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0926_),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1477_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0927_),
    .B(\tt_um_rejunity_sn76489.chan[3].attenuation.in ),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1478_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0928_),
    .B(_0920_),
    .A(_0927_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1479_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0928_),
    .A(_0926_),
    .B(_0923_),
    .C(_0915_),
    .Y(_0929_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1480_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0921_),
    .A(_0919_),
    .Y(_0930_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_4 _1481_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0931_),
    .A(_0918_),
    .B(_0925_),
    .C(_0929_),
    .D(_0930_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1482_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0931_),
    .A(_0914_),
    .Y(_0932_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1483_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0933_),
    .A(_0932_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1484_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ),
    .Y(_0934_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1485_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[0].attenuation.in ),
    .Y(_0935_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1486_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0935_),
    .Y(_0936_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1487_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0937_),
    .B(_0936_),
    .A(_0934_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1488_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0937_),
    .Y(_0938_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1489_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0939_),
    .B(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ),
    .A(_0935_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1490_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0940_),
    .B(_0935_),
    .A(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _1491_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_0940_),
    .B(_0939_),
    .A(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ),
    .Y(_0941_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1492_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ),
    .Y(_0942_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1493_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0943_),
    .B(_0936_),
    .A(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1494_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ),
    .Y(_0944_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1495_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0945_),
    .B(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ),
    .A(\tt_um_rejunity_sn76489.chan[0].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1496_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0946_),
    .B(_0945_),
    .A(_0944_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _1497_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_0946_),
    .B(_0943_),
    .A(_0942_),
    .Y(_0947_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1498_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0948_),
    .A(_0938_),
    .B(_0941_),
    .C(_0947_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1499_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .Y(_0949_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1500_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0950_),
    .B(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .A(_0949_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1501_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0950_),
    .Y(_0951_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1502_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0952_),
    .B(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1503_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0952_),
    .Y(_0953_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1504_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0953_),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .Y(_0954_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_4 _1505_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0955_),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .B(_0949_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1506_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0956_),
    .B(_0954_),
    .A(_0955_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1507_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0952_),
    .Y(_0957_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1508_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .Y(_0958_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1509_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0959_),
    .B(_0949_),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _1510_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_0959_),
    .B(_0950_),
    .A(_0958_),
    .Y(_0960_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1511_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0961_),
    .B(_0960_),
    .A(_0957_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _1512_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0962_),
    .A(_0951_),
    .B(_0954_),
    .C(_0956_),
    .D(_0961_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1513_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0962_),
    .Y(_0963_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1514_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0945_),
    .Y(_0964_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _1515_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0965_),
    .A(_0942_),
    .B(_0964_),
    .C(_0939_),
    .D(_0934_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1516_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0966_),
    .B(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .A(_0935_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1517_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0967_),
    .C(_0966_),
    .B(_0940_),
    .A(_0937_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_4 _1518_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0968_),
    .C(_0943_),
    .B(_0964_),
    .A(_0942_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1519_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0969_),
    .A(_0944_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1520_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0965_),
    .B(_0967_),
    .C(_0968_),
    .D(_0969_),
    .Y(_0970_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1521_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0971_),
    .A(_0970_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1522_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0972_),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1523_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .Y(_0973_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1524_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0952_),
    .A(_0972_),
    .B(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .C(_0973_),
    .Y(_0974_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1525_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0975_),
    .B(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .A(_0973_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1526_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0976_),
    .C(_0975_),
    .B(_0953_),
    .A(_0958_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_4 _1527_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0977_),
    .C(_0955_),
    .B(_0952_),
    .A(_0958_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1528_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0972_),
    .Y(_0978_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_4 _1529_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0979_),
    .A(_0974_),
    .B(_0976_),
    .C(_0977_),
    .D(_0978_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1530_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0980_),
    .B(_0949_),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1531_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0981_),
    .A(_0980_),
    .B(_0959_),
    .C(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _1532_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0955_),
    .B(_0974_),
    .C(_0981_),
    .Y(_0982_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1533_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0983_),
    .B(_0959_),
    .A(_0953_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1534_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0984_),
    .B(_0977_),
    .A(_0983_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1535_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0985_),
    .B(_0940_),
    .A(_0937_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1536_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0939_),
    .Y(_0986_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1537_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0987_),
    .C(_0986_),
    .B(_0964_),
    .A(_0969_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _1538_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0988_),
    .A(_0985_),
    .B(_0968_),
    .C(_0987_),
    .D(_0967_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1539_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0989_),
    .A(_0982_),
    .B(_0984_),
    .C(_0988_));
 gf180mcu_as_sc_mcu7t3v3__maj3_4 _1540_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0990_),
    .A(_0971_),
    .B(_0979_),
    .C(_0989_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1541_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0991_),
    .A(_0948_),
    .B(_0963_),
    .C(_0990_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1542_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .Y(_0992_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1543_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0993_),
    .C(_0975_),
    .B(_0951_),
    .A(_0992_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1544_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .Y(_0994_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1545_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0995_),
    .C(_0994_),
    .B(_0959_),
    .A(_0980_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _1546_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_0953_),
    .B(_0992_),
    .A(_0995_),
    .Y(_0996_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1547_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0996_),
    .A(_0993_),
    .Y(_0997_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1548_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0998_),
    .A(_0986_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1549_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .Y(_0999_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1550_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1000_),
    .C(_0999_),
    .B(_0940_),
    .A(_0998_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1551_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0946_),
    .Y(_1001_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1552_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1002_),
    .A(_0944_),
    .B(_0986_),
    .C(_0966_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1553_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1003_),
    .B(_1002_),
    .A(_1001_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1554_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1004_),
    .A(_0938_),
    .B(_1000_),
    .C(_1003_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1555_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1004_),
    .A(_0997_),
    .Y(_1005_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1556_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1004_),
    .A(_0997_),
    .Y(_1006_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1557_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1007_),
    .B(_1006_),
    .A(_1005_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1558_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1007_),
    .A(_0991_),
    .Y(_1008_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1559_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1008_),
    .A(_0933_),
    .Y(_1009_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1560_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1010_),
    .B(_0924_),
    .A(_0927_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1561_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0927_),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ),
    .Y(_1011_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1562_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1011_),
    .A(_0921_),
    .Y(_1012_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1563_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ),
    .Y(_1013_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1564_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1014_),
    .B(_1013_),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1565_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1014_),
    .Y(_1015_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1566_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1016_),
    .C(_0916_),
    .B(_1014_),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _1567_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0919_),
    .B(_0923_),
    .C(_1015_),
    .Y(_1017_),
    .D(_1016_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1568_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1018_),
    .A(_1010_),
    .B(_1012_),
    .C(_1017_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1569_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1019_),
    .A(_1018_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1570_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1020_),
    .A(_0896_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1571_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1021_),
    .B(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .A(_0899_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1572_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1022_),
    .B(_1021_),
    .A(_1020_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1573_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1022_),
    .A(_0909_),
    .Y(_1023_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1574_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .Y(_1024_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1575_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1025_),
    .B(_0898_),
    .A(_0896_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1576_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1025_),
    .A(_1024_),
    .Y(_1026_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1577_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1027_),
    .A(_0901_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_4 _1578_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1028_),
    .A(_0905_),
    .B(_1023_),
    .C(_1026_),
    .D(_1027_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1579_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1029_),
    .B(_0941_),
    .A(_0938_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1580_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1030_),
    .B(_0947_),
    .A(_1029_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1581_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0962_),
    .A(_1030_),
    .Y(_1031_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1582_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1031_),
    .A(_0990_),
    .Y(_1032_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1583_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1033_),
    .A(_1019_),
    .B(_1028_),
    .C(_1032_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1584_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1028_),
    .A(_1018_),
    .Y(_1034_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1585_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1035_),
    .A(_1034_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1586_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1035_),
    .A(_1032_),
    .Y(_1036_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1587_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ),
    .Y(_1037_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1588_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1038_),
    .B(_0921_),
    .A(_0923_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _1589_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0917_),
    .B(_0928_),
    .C(_1038_),
    .Y(_1039_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1590_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0916_),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .Y(_1040_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_4 _1591_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1041_),
    .A(_1037_),
    .B(_1015_),
    .C(_1039_),
    .D(_1040_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1592_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0900_),
    .Y(_1042_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _1593_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1043_),
    .A(_1024_),
    .B(_0898_),
    .C(_1021_),
    .D(_0903_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1594_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1044_),
    .C(_0900_),
    .B(_0897_),
    .A(_1024_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1595_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1044_),
    .A(_1020_),
    .Y(_1045_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1596_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1045_),
    .A(_1042_),
    .B(_0911_),
    .C(_1043_),
    .Y(_1046_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1597_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1046_),
    .Y(_1047_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1598_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1048_),
    .B(_1047_),
    .A(_1041_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1599_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0979_),
    .A(_0970_),
    .Y(_1049_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1600_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1049_),
    .A(_0989_),
    .Y(_1050_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1601_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1037_),
    .B(_1015_),
    .C(_1039_),
    .D(_1040_),
    .Y(_1051_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1602_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1046_),
    .A(_1051_),
    .Y(_1052_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1603_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1053_),
    .B(_1052_),
    .A(_1050_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1604_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1054_),
    .B(_1053_),
    .A(_1048_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1605_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0928_),
    .A(_0917_),
    .Y(_1055_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1606_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1056_),
    .A(_0927_),
    .B(_0924_),
    .C(_1013_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1607_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1057_),
    .C(_0917_),
    .B(_1015_),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1608_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1057_),
    .A(_0928_),
    .Y(_1058_));
 gf180mcu_as_sc_mcu7t3v3__ao31_4 _1609_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1058_),
    .A(_1038_),
    .B(_1055_),
    .C(_1056_),
    .Y(_1059_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1610_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1060_),
    .B(_1044_),
    .A(_0911_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1611_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1061_),
    .B(_0897_),
    .A(_1020_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1612_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1061_),
    .A(_1042_),
    .Y(_1062_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _1613_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0907_),
    .B(_0911_),
    .C(_1062_),
    .Y(_1063_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1614_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1064_),
    .B(_1063_),
    .A(_1060_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1615_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0984_),
    .A(_0982_),
    .Y(_1065_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1616_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0985_),
    .B(_0968_),
    .C(_0987_),
    .D(_0967_),
    .Y(_1066_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1617_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1066_),
    .A(_1065_),
    .Y(_1067_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1618_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1068_),
    .A(_1059_),
    .B(_1064_),
    .C(_1067_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1619_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1052_),
    .A(_1050_),
    .Y(_1069_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1620_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1070_),
    .B(_1069_),
    .A(_1068_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1621_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1071_),
    .A(_1036_),
    .B(_1054_),
    .C(_1070_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1622_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1072_),
    .A(_1009_),
    .B(_1033_),
    .C(_1071_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1623_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1073_),
    .B(_1040_),
    .A(_1037_));
 gf180mcu_as_sc_mcu7t3v3__ao31_4 _1624_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1073_),
    .A(_1038_),
    .B(_1055_),
    .C(_1056_),
    .Y(_1074_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1625_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1022_),
    .A(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ),
    .Y(_1075_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1626_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1075_),
    .A(_1063_),
    .Y(_1076_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1627_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1076_),
    .A(_1074_),
    .Y(_1077_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1628_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0955_),
    .Y(_1078_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1629_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0994_),
    .B(_0992_),
    .C(_0980_),
    .Y(_1079_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1630_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1079_),
    .A(_1078_),
    .B(_0974_),
    .C(_0981_),
    .Y(_1080_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1631_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1081_),
    .A(_0999_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1632_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0986_),
    .A(_0969_),
    .Y(_1082_));
 gf180mcu_as_sc_mcu7t3v3__ao22_4 _1633_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1081_),
    .B(_1082_),
    .C(_0967_),
    .D(_0987_),
    .Y(_1083_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1634_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1084_),
    .A(_1083_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1635_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1084_),
    .A(_1080_),
    .Y(_1085_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1636_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0963_),
    .A(_0948_),
    .Y(_1086_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1637_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1005_),
    .A(_1086_),
    .B(_0990_),
    .C(_1006_),
    .Y(_1087_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1638_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1087_),
    .A(_1085_),
    .Y(_1088_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1639_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1088_),
    .A(_1077_),
    .Y(_1089_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1640_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1090_),
    .B(_1007_),
    .A(_0991_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1641_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1007_),
    .A(_0991_),
    .Y(_1091_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1642_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0931_),
    .A(_0914_),
    .Y(_1092_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1643_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1092_),
    .A(_0933_),
    .B(_1090_),
    .C(_1091_),
    .Y(_1093_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1644_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1093_),
    .A(_1089_),
    .Y(_1094_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1645_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1095_),
    .B(_1094_),
    .A(_1072_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1646_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1094_),
    .A(_1072_),
    .Y(_1096_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1647_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1096_),
    .A(_1095_),
    .Y(_1097_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1648_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1097_),
    .Y(net18));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1649_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1098_),
    .B(_1089_),
    .A(_1093_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1650_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1099_),
    .A(_1072_),
    .B(_1094_),
    .C(_1098_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1651_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1023_),
    .A(_1042_),
    .Y(_1100_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1652_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1100_),
    .A(_1061_),
    .Y(_1101_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1653_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1010_),
    .Y(_1102_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _1654_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0918_),
    .B(_1102_),
    .C(_1011_),
    .Y(_1103_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1655_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1103_),
    .A(_0922_),
    .Y(_1104_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1656_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1104_),
    .A(_1101_),
    .Y(_1105_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1657_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1106_),
    .B(_0957_),
    .A(_0978_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1658_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1078_),
    .A(_0960_),
    .Y(_1107_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1659_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1107_),
    .A(_1106_),
    .Y(_1108_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1660_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0964_),
    .A(_0969_),
    .Y(_1109_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1661_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1110_),
    .B(_0943_),
    .A(_0941_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1662_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1110_),
    .A(_1109_),
    .Y(_1111_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1663_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1111_),
    .A(_1108_),
    .Y(_1112_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1664_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1080_),
    .Y(_1113_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _1665_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1086_),
    .B(_0990_),
    .C(_1006_),
    .Y(_1114_),
    .D(_1005_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1666_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1115_),
    .A(_1113_),
    .B(_1083_),
    .C(_1114_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1667_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1115_),
    .A(_1112_),
    .Y(_1116_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1668_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1116_),
    .A(_1105_),
    .Y(_1117_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1669_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1118_),
    .B(_1075_),
    .A(_1063_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1670_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1119_),
    .A(_1074_),
    .B(_1118_),
    .C(_1088_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1671_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1119_),
    .A(_1117_),
    .Y(_1120_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1672_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1120_),
    .A(_1099_),
    .Y(_1121_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1673_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1121_),
    .Y(net19));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1674_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1122_),
    .A(_1099_),
    .B(_1117_),
    .C(_1119_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1675_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1123_),
    .A(_1122_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1676_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1124_),
    .A(_1012_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1677_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1057_),
    .A(_0925_),
    .Y(_1125_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1678_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1125_),
    .A(_0918_),
    .B(_0930_),
    .C(_1124_),
    .Y(_1126_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1679_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1127_),
    .B(_1022_),
    .A(_0906_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _1680_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1128_),
    .A(_0902_),
    .B(_1043_),
    .C(_1062_),
    .D(_1127_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1681_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1128_),
    .A(_1126_),
    .Y(_1129_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1682_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1130_),
    .A(_0978_),
    .B(_0951_),
    .C(_0957_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1683_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1131_),
    .A(_0977_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1684_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1132_),
    .C(_1131_),
    .B(_1106_),
    .A(_0951_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1685_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1132_),
    .A(_1130_),
    .B(_1078_),
    .C(_1106_),
    .Y(_1133_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1686_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1134_),
    .B(_1082_),
    .A(_0938_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1687_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1135_),
    .C(_0966_),
    .B(_1134_),
    .A(_1001_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1688_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1135_),
    .A(_0966_),
    .B(_1001_),
    .C(_0965_),
    .Y(_1136_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1689_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1137_),
    .B(_1136_),
    .A(_1133_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1690_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1136_),
    .A(_1133_),
    .Y(_1138_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1691_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1139_),
    .B(_1138_),
    .A(_1137_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1692_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1140_),
    .B(_1114_),
    .A(_1085_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1693_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1108_),
    .Y(_1141_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1694_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1111_),
    .Y(_1142_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _1695_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1143_),
    .A(_1113_),
    .B(_1083_),
    .C(_1141_),
    .D(_1142_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1696_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1144_),
    .B(_1142_),
    .A(_1141_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1697_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1145_),
    .C(_1144_),
    .B(_1143_),
    .A(_1140_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1698_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1145_),
    .A(_1139_),
    .Y(_1146_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1699_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1146_),
    .A(_1129_),
    .Y(_1147_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1700_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1148_),
    .A(_1101_),
    .B(_1104_),
    .C(_1116_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1701_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1148_),
    .A(_1147_),
    .Y(_1149_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1702_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1149_),
    .A(_1123_),
    .Y(_1150_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1703_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1150_),
    .Y(net20));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1704_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1151_),
    .B(_1012_),
    .A(_1102_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1705_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ),
    .B(_0922_),
    .C(_1151_),
    .D(_1057_),
    .Y(_1152_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1706_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1153_),
    .B(_1023_),
    .A(_0906_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1707_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0898_),
    .A(_1020_),
    .Y(_1154_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _1708_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1155_),
    .A(_1153_),
    .B(_1044_),
    .C(_1154_),
    .D(_0913_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1709_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1155_),
    .A(_1152_),
    .Y(_1156_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1710_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1157_),
    .A(_1156_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1711_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0957_),
    .A(_0978_),
    .Y(_1158_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_4 _1712_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1159_),
    .A(_0961_),
    .B(_0977_),
    .C(_1158_),
    .D(_0994_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_4 _1713_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1160_),
    .A(_1029_),
    .B(_0968_),
    .C(_1109_),
    .D(_0999_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1714_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1161_),
    .B(_1160_),
    .A(_1159_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1715_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1162_),
    .B(_1160_),
    .A(_1159_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _1716_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1163_),
    .B(_1162_),
    .A(_1161_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1717_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1164_),
    .A(_1137_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1718_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1165_),
    .C(_1164_),
    .B(_1145_),
    .A(_1138_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1719_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1165_),
    .A(_1163_),
    .Y(_1166_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1720_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1166_),
    .A(_1157_),
    .Y(_1167_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1721_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0902_),
    .B(_1043_),
    .C(_1062_),
    .D(_1127_),
    .Y(_1168_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1722_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1169_),
    .A(_1126_),
    .B(_1168_),
    .C(_1146_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1723_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1169_),
    .A(_1167_),
    .Y(_1170_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1724_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1171_),
    .A(_1147_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1725_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1172_),
    .A(_1122_),
    .B(_1171_),
    .C(_1148_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1726_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1173_),
    .B(_1172_),
    .A(_1170_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1727_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1172_),
    .A(_1170_),
    .Y(_1174_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1728_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1174_),
    .A(_1173_),
    .Y(_1175_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1729_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1175_),
    .Y(net21));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1730_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1176_),
    .B(_1167_),
    .A(_1169_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1731_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1177_),
    .C(_1176_),
    .B(_1172_),
    .A(_1170_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1732_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1178_),
    .B(_1016_),
    .A(_1102_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1733_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0909_),
    .A(_0902_),
    .Y(_1179_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1734_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1179_),
    .A(_1178_),
    .Y(_1180_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1735_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1143_),
    .A(_1144_),
    .Y(_1181_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1736_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1182_),
    .B(_1181_),
    .A(_1137_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1737_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1161_),
    .A(_1138_),
    .B(_1162_),
    .C(_1182_),
    .Y(_1183_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1738_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1184_),
    .B(_0954_),
    .A(_0995_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1739_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1000_),
    .A(_1001_),
    .Y(_1185_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1740_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1185_),
    .A(_1184_),
    .Y(_1186_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1741_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1186_),
    .A(_1183_),
    .Y(_1187_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1742_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1187_),
    .A(_1180_),
    .Y(_1188_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1743_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1153_),
    .B(_1044_),
    .C(_1154_),
    .D(_0913_),
    .Y(_1189_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1744_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1190_),
    .B(_1189_),
    .A(_1152_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1745_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1166_),
    .A(_1157_),
    .Y(_1191_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1746_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1192_),
    .B(_1191_),
    .A(_1190_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1747_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1192_),
    .A(_1188_),
    .Y(_1193_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1748_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1193_),
    .A(_1177_),
    .Y(_1194_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1749_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1194_),
    .Y(net22));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1750_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1191_),
    .A(_1190_),
    .Y(_1195_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1751_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1196_),
    .A(_1177_),
    .B(_1188_),
    .C(_1195_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1752_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1197_),
    .B(_0918_),
    .A(_1013_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1753_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1198_),
    .A(_1197_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1754_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1199_),
    .B(_1042_),
    .A(_0903_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1755_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1199_),
    .A(_1198_),
    .Y(_1200_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1756_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1201_),
    .B(_1078_),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1757_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1202_),
    .B(_0943_),
    .A(_0934_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1758_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1202_),
    .A(_1201_),
    .Y(_1203_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1759_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1204_),
    .A(_1183_),
    .B(_1184_),
    .C(_1185_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1760_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1204_),
    .A(_1203_),
    .Y(_1205_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1761_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1205_),
    .A(_1200_),
    .Y(_1206_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1762_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1016_),
    .A(_1102_),
    .Y(_1207_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1763_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1208_),
    .A(_1207_),
    .B(_1179_),
    .C(_1187_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1764_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1208_),
    .A(_1206_),
    .Y(_1209_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1765_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1209_),
    .A(_1196_),
    .Y(_1210_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1766_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1210_),
    .Y(net23));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1767_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1211_),
    .A(_1208_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1768_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1212_),
    .A(_1196_),
    .B(_1206_),
    .C(_1211_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1769_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1199_),
    .Y(_1213_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1770_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1214_),
    .A(_1197_),
    .B(_1213_),
    .C(_1205_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1771_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1201_),
    .Y(_1215_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1772_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1202_),
    .Y(_1216_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1773_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1217_),
    .A(_1215_),
    .B(_1216_),
    .C(_1204_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1774_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1217_),
    .A(_1214_),
    .Y(_1218_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1775_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1219_),
    .B(_1218_),
    .A(_1212_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1776_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1218_),
    .A(_1212_),
    .Y(_1220_));
 gf180mcu_as_sc_mcu7t3v3__nor2_4 _1777_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(net24),
    .A(_1219_),
    .B(_1220_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1778_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1221_),
    .A(_1214_),
    .B(_1217_),
    .C(_1219_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1779_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1221_),
    .Y(net25));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1780_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net11),
    .Y(_1222_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1781_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1222_),
    .Y(_1223_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1782_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1223_),
    .Y(_1224_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1783_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[4] ),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[3] ),
    .Y(_1225_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1784_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1226_),
    .B(_1225_),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1785_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1226_),
    .Y(_1227_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1786_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1227_),
    .Y(_1228_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1787_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1228_),
    .A(_1224_),
    .Y(_1229_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1788_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1229_),
    .Y(_0000_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1789_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net11),
    .Y(_1230_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1790_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1230_),
    .Y(_1231_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1791_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1232_),
    .B(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[4] ),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1792_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1233_),
    .B(_1232_),
    .A(_1231_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1793_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1234_),
    .B(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[1] ),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1794_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[1] ),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[0] ),
    .Y(_1235_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1795_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1233_),
    .B(_1234_),
    .C(_1235_),
    .Y(_1236_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1796_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1236_),
    .Y(_0001_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1797_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1237_),
    .B(_1235_),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1798_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1235_),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[2] ),
    .Y(_1238_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1799_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1233_),
    .B(_1237_),
    .C(_1238_),
    .Y(_1239_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1800_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1239_),
    .Y(_0002_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1801_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1238_),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[3] ),
    .Y(_1240_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1802_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0003_),
    .B(_1240_),
    .A(_1233_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1803_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1241_),
    .C(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[4] ),
    .B(_1238_),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1804_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0004_),
    .B(_1241_),
    .A(_1233_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1805_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1242_),
    .A(net8));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1806_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1243_),
    .A(net9));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1807_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1244_),
    .B(_1243_),
    .A(net10));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1808_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1244_),
    .A(_1242_),
    .Y(_1245_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1809_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1245_),
    .Y(_1246_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1810_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net7),
    .Y(_1247_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1811_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net6),
    .Y(_1248_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1812_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1249_),
    .B(_1248_),
    .A(_1247_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1813_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1249_),
    .Y(_1250_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1814_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1251_),
    .B(_1250_),
    .A(_1246_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1815_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[0]),
    .Y(_1252_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1816_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1245_),
    .Y(_1253_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1817_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1254_),
    .A(net11));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1818_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1254_),
    .Y(_1255_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1819_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1255_),
    .Y(_1256_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1820_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1256_),
    .A(_1252_),
    .B(_1253_),
    .C(_1249_),
    .Y(_1257_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1821_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1258_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][0] ),
    .B(_1251_),
    .C(_1257_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1822_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1258_),
    .Y(_0005_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1823_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1259_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1824_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1260_),
    .A(net3));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1825_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1260_),
    .Y(_1261_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1826_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1253_),
    .Y(_1262_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1827_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1249_),
    .Y(_1263_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1828_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1254_),
    .Y(_1264_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1829_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1264_),
    .Y(_1265_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1830_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1265_),
    .Y(_1266_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1831_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1266_),
    .A(_1261_),
    .B(_1262_),
    .C(_1263_),
    .Y(_1267_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1832_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0006_),
    .C(_1267_),
    .B(_1251_),
    .A(_1259_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1833_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1268_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][2] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1834_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1269_),
    .A(net4));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1835_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1269_),
    .Y(_1270_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1836_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1266_),
    .A(_1270_),
    .B(_1262_),
    .C(_1263_),
    .Y(_1271_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1837_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0007_),
    .C(_1271_),
    .B(_1251_),
    .A(_1268_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1838_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1272_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][3] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1839_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1273_),
    .A(net5));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1840_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1273_),
    .Y(_1274_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1841_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1265_),
    .Y(_1275_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1842_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1275_),
    .A(_1274_),
    .B(_1262_),
    .C(_1263_),
    .Y(_1276_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1843_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0008_),
    .C(_1276_),
    .B(_1251_),
    .A(_1272_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1844_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1277_),
    .A(net6));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1845_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1277_),
    .A(_1247_),
    .Y(_1278_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1846_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1278_),
    .Y(_1279_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1847_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1280_),
    .B(_1279_),
    .A(_1253_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1848_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1256_),
    .A(_1252_),
    .B(_1253_),
    .C(_1279_),
    .Y(_1281_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1849_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1282_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ),
    .B(_1280_),
    .C(_1281_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1850_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1282_),
    .Y(_0009_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1851_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1283_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1852_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1278_),
    .Y(_1284_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1853_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1275_),
    .A(_1261_),
    .B(_1246_),
    .C(_1284_),
    .Y(_1285_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1854_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0010_),
    .C(_1285_),
    .B(_1280_),
    .A(_1283_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1855_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1286_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1856_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1275_),
    .A(_1270_),
    .B(_1246_),
    .C(_1284_),
    .Y(_1287_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1857_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0011_),
    .C(_1287_),
    .B(_1280_),
    .A(_1286_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1858_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1288_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1859_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1275_),
    .A(_1274_),
    .B(_1246_),
    .C(_1284_),
    .Y(_1289_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1860_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0012_),
    .C(_1289_),
    .B(_1280_),
    .A(_1288_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1861_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1244_),
    .Y(_1290_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1862_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1290_),
    .A(net8),
    .Y(_1291_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1863_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1291_),
    .Y(_1292_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1864_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1293_),
    .B(_1292_),
    .A(_1250_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1865_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[0]),
    .Y(_1294_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1866_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1256_),
    .A(_1294_),
    .B(_1249_),
    .C(_1292_),
    .Y(_1295_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1867_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1296_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ),
    .B(_1293_),
    .C(_1295_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1868_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1296_),
    .Y(_0013_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1869_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1297_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1870_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1291_),
    .Y(_1298_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1871_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1265_),
    .Y(_1299_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1872_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1299_),
    .A(_1261_),
    .B(_1263_),
    .C(_1298_),
    .Y(_1300_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1873_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0014_),
    .C(_1300_),
    .B(_1293_),
    .A(_1297_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1874_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1301_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1875_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1299_),
    .A(_1270_),
    .B(_1250_),
    .C(_1298_),
    .Y(_1302_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1876_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0015_),
    .C(_1302_),
    .B(_1293_),
    .A(_1301_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1877_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1303_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1878_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1299_),
    .A(_1274_),
    .B(_1250_),
    .C(_1298_),
    .Y(_1304_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1879_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0016_),
    .C(_1304_),
    .B(_1293_),
    .A(_1303_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1880_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1265_),
    .Y(_1305_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1881_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1305_),
    .Y(_1306_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1882_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1307_),
    .B(_1064_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1883_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1064_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[0] ),
    .Y(_1308_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1884_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1306_),
    .B(_1307_),
    .C(_1308_),
    .Y(_1309_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1885_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1309_),
    .Y(_0017_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1886_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1047_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[1] ),
    .Y(_1310_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1887_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1311_),
    .B(_1047_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[1] ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1888_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1312_),
    .C(_1308_),
    .B(_1311_),
    .A(_1310_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1889_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1264_),
    .Y(_1313_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1890_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1313_),
    .Y(_1314_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1891_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1314_),
    .A(_1308_),
    .B(_1310_),
    .C(_1311_),
    .Y(_1315_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1892_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0018_),
    .B(_1315_),
    .A(_1312_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _1893_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0906_),
    .B(_1023_),
    .C(_1026_),
    .D(_1027_),
    .Y(_1316_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1894_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1316_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[2] ),
    .Y(_1317_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1895_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1318_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[1] ),
    .B(_1047_),
    .C(_1308_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1896_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1318_),
    .A(_1317_),
    .Y(_1319_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1897_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1254_),
    .Y(_1320_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1898_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1320_),
    .Y(_1321_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1899_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1321_),
    .Y(_1322_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1900_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1323_),
    .C(_1322_),
    .B(_1318_),
    .A(_1317_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1901_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1323_),
    .A(_1319_),
    .Y(_1324_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1902_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1324_),
    .Y(_0019_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1903_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1325_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1904_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0914_),
    .A(_1325_),
    .Y(_1326_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1905_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1327_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[2] ),
    .B(_1028_),
    .C(_1318_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1906_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1327_),
    .A(_1326_),
    .Y(_1328_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1907_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1329_),
    .C(_1322_),
    .B(_1327_),
    .A(_1326_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1908_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1329_),
    .A(_1328_),
    .Y(_1330_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1909_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1330_),
    .Y(_0020_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1910_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1076_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[4] ),
    .Y(_1331_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1911_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1332_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[3] ),
    .B(_0914_),
    .C(_1327_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1912_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1332_),
    .A(_1331_),
    .Y(_1333_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1913_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1334_),
    .C(_1322_),
    .B(_1332_),
    .A(_1331_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1914_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1334_),
    .A(_1333_),
    .Y(_1335_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1915_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1335_),
    .Y(_0021_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1916_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1336_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[4] ),
    .B(_1118_),
    .C(_1332_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1917_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1337_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1918_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1101_),
    .A(_1337_),
    .Y(_1338_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1919_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1222_),
    .Y(_1339_));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 _1920_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1339_),
    .Y(_1340_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1921_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1338_),
    .A(_1336_),
    .Y(_1341_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1922_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1342_),
    .B(_1341_),
    .A(_1340_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1923_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0022_),
    .C(_1342_),
    .B(_1338_),
    .A(_1336_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1924_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1128_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[6] ),
    .Y(_1343_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1925_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1344_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[5] ),
    .B(_1101_),
    .C(_1336_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1926_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1344_),
    .A(_1343_),
    .Y(_1345_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1927_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1321_),
    .Y(_1346_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1928_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1347_),
    .C(_1346_),
    .B(_1344_),
    .A(_1343_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1929_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1347_),
    .A(_1345_),
    .Y(_1348_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1930_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1348_),
    .Y(_0023_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1931_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1264_),
    .Y(_1349_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1932_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1349_),
    .Y(_1350_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1933_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1350_),
    .Y(_1351_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1934_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1155_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[7] ),
    .Y(_1352_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1935_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1353_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[6] ),
    .B(_1168_),
    .C(_1344_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1936_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1354_),
    .B(_1353_),
    .A(_1352_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1937_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1353_),
    .A(_1352_),
    .Y(_1355_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1938_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1351_),
    .B(_1354_),
    .C(_1355_),
    .Y(_1356_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1939_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1356_),
    .Y(_0024_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1940_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1357_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1941_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1179_),
    .A(_1357_),
    .Y(_1358_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1942_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1359_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[7] ),
    .B(_1189_),
    .C(_1355_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1943_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1360_),
    .B(_1359_),
    .A(_1358_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1944_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1359_),
    .A(_1358_),
    .Y(_1361_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1945_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1351_),
    .B(_1360_),
    .C(_1361_),
    .Y(_1362_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1946_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1362_),
    .Y(_0025_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1947_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1213_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[9] ),
    .Y(_1363_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1948_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1364_),
    .B(_1213_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1949_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1364_),
    .A(_1363_),
    .Y(_1365_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1950_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1366_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[8] ),
    .B(_1179_),
    .C(_1361_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1951_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1366_),
    .A(_1365_),
    .Y(_1367_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1952_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1368_),
    .C(_1346_),
    .B(_1366_),
    .A(_1365_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1953_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1368_),
    .A(_1367_),
    .Y(_1369_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1954_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1369_),
    .Y(_0026_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1955_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1370_),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[9] ),
    .B(_1213_),
    .C(_1366_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1956_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1363_),
    .A(_1223_),
    .Y(_1371_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1957_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1371_),
    .A(_1370_),
    .Y(_1372_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1958_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1372_),
    .Y(_0027_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1959_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1373_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1960_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1374_),
    .B(_1065_),
    .A(_1373_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _1961_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1314_),
    .A(_1373_),
    .B(_0982_),
    .C(_0984_),
    .Y(_1375_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1962_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0028_),
    .B(_1375_),
    .A(_1374_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1963_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0979_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[1] ),
    .Y(_1376_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1964_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1376_),
    .A(_1374_),
    .Y(_1377_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1965_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1378_),
    .B(_1377_),
    .A(_1340_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1966_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0029_),
    .C(_1378_),
    .B(_1376_),
    .A(_1374_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1967_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0963_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[2] ),
    .Y(_1379_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1968_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1380_),
    .A(_0979_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1969_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1381_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[1] ),
    .B(_1380_),
    .C(_1374_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _1970_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1382_),
    .B(_1381_),
    .A(_1379_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1971_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1381_),
    .A(_1379_),
    .Y(_1383_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _1972_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1351_),
    .B(_1382_),
    .C(_1383_),
    .Y(_1384_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1973_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1384_),
    .Y(_0030_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1974_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0997_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[3] ),
    .Y(_1385_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1975_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1386_),
    .A(_0963_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1976_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1387_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[2] ),
    .B(_1386_),
    .C(_1383_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1977_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1387_),
    .A(_1385_),
    .Y(_1388_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1978_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1389_),
    .C(_1346_),
    .B(_1387_),
    .A(_1385_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1979_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1389_),
    .A(_1388_),
    .Y(_1390_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1980_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1390_),
    .Y(_0031_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1981_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1391_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1982_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1113_),
    .A(_1391_),
    .Y(_1392_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _1983_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1393_),
    .B(_0997_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _1984_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1394_),
    .A(_1385_),
    .B(_1387_),
    .C(_1393_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1985_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1394_),
    .A(_1392_),
    .Y(_1395_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1986_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1396_),
    .C(_1346_),
    .B(_1394_),
    .A(_1392_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _1987_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1396_),
    .A(_1395_),
    .Y(_1397_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _1988_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1397_),
    .Y(_0032_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1989_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1398_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[4] ),
    .B(_1113_),
    .C(_1394_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1990_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1399_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1991_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1141_),
    .A(_1399_),
    .Y(_1400_));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 _1992_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1230_),
    .Y(_1401_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1993_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1400_),
    .A(_1398_),
    .Y(_1402_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _1994_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1403_),
    .B(_1402_),
    .A(_1401_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _1995_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0033_),
    .C(_1403_),
    .B(_1400_),
    .A(_1398_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _1996_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1404_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _1997_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1133_),
    .A(_1404_),
    .Y(_1405_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _1998_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1406_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[5] ),
    .B(_1141_),
    .C(_1398_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _1999_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1406_),
    .A(_1405_),
    .Y(_1407_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2000_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1321_),
    .Y(_1408_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2001_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1409_),
    .C(_1408_),
    .B(_1406_),
    .A(_1405_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2002_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1409_),
    .A(_1407_),
    .Y(_1410_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2003_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1410_),
    .Y(_0034_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2004_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1159_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[7] ),
    .Y(_1411_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2005_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1412_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[6] ),
    .B(_1133_),
    .C(_1406_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2006_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1413_),
    .B(_1412_),
    .A(_1411_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2007_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1412_),
    .A(_1411_),
    .Y(_1414_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2008_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1351_),
    .B(_1413_),
    .C(_1414_),
    .Y(_1415_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2009_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1415_),
    .Y(_0035_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2010_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1350_),
    .Y(_1416_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2011_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1417_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2012_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1184_),
    .A(_1417_),
    .Y(_1418_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _2013_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1419_),
    .B(_1159_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2014_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1414_),
    .A(_1419_),
    .Y(_1420_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2015_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1421_),
    .B(_1420_),
    .A(_1418_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2016_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1420_),
    .A(_1418_),
    .Y(_1422_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2017_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1416_),
    .B(_1421_),
    .C(_1422_),
    .Y(_1423_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2018_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1423_),
    .Y(_0036_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2019_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1424_),
    .B(_1215_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2020_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1215_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[9] ),
    .Y(_1425_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2021_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1426_),
    .B(_1425_),
    .A(_1424_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2022_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1427_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[8] ),
    .B(_1184_),
    .C(_1422_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2023_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1427_),
    .A(_1426_),
    .Y(_1428_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2024_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1429_),
    .C(_1408_),
    .B(_1427_),
    .A(_1426_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2025_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1429_),
    .A(_1428_),
    .Y(_1430_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2026_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1430_),
    .Y(_0037_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2027_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1431_),
    .C(_1427_),
    .B(_1215_),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2028_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1416_),
    .B(_1424_),
    .C(_1431_),
    .Y(_1432_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2029_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1432_),
    .Y(_0038_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2030_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1433_),
    .B(_1066_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2031_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1066_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[0] ),
    .Y(_1434_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2032_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1416_),
    .B(_1433_),
    .C(_1434_),
    .Y(_1435_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2033_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1435_),
    .Y(_0039_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2034_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0971_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[1] ),
    .Y(_1436_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2035_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1436_),
    .A(_1434_),
    .Y(_1437_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2036_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1438_),
    .C(_1408_),
    .B(_1436_),
    .A(_1434_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2037_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1438_),
    .A(_1437_),
    .Y(_1439_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2038_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1439_),
    .Y(_0040_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2039_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0948_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[2] ),
    .Y(_1440_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2040_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1441_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[1] ),
    .B(_0970_),
    .C(_1434_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2041_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1441_),
    .A(_1440_),
    .Y(_1442_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2042_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_1443_),
    .C(_1408_),
    .B(_1441_),
    .A(_1440_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2043_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1443_),
    .A(_1442_),
    .Y(_1444_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2044_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1444_),
    .Y(_0041_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2045_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1004_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[3] ),
    .Y(_1445_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2046_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0193_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[2] ),
    .B(_1030_),
    .C(_1441_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2047_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0193_),
    .A(_1445_),
    .Y(_0194_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2048_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1320_),
    .Y(_0195_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2049_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0195_),
    .Y(_0196_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2050_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0197_),
    .C(_0196_),
    .B(_0193_),
    .A(_1445_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2051_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0197_),
    .A(_0194_),
    .Y(_0198_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2052_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0198_),
    .Y(_0042_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2053_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1084_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[4] ),
    .Y(_0199_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2054_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0200_),
    .A(_1004_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2055_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0201_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[3] ),
    .B(_0200_),
    .C(_0193_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2056_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0201_),
    .A(_0199_),
    .Y(_0202_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2057_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0203_),
    .C(_0196_),
    .B(_0201_),
    .A(_0199_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2058_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0203_),
    .A(_0202_),
    .Y(_0204_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2059_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0204_),
    .Y(_0043_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2060_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0205_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[4] ),
    .B(_1083_),
    .C(_0201_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2061_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0206_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2062_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1142_),
    .A(_0206_),
    .Y(_0207_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2063_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0207_),
    .A(_0205_),
    .Y(_0208_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2064_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0209_),
    .B(_0208_),
    .A(_1401_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2065_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0044_),
    .C(_0209_),
    .B(_0207_),
    .A(_0205_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2066_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0210_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2067_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1136_),
    .A(_0210_),
    .Y(_0211_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2068_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0212_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[5] ),
    .B(_1142_),
    .C(_0205_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2069_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0212_),
    .A(_0211_),
    .Y(_0213_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2070_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0214_),
    .C(_0196_),
    .B(_0212_),
    .A(_0211_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2071_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0214_),
    .A(_0213_),
    .Y(_0215_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2072_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0215_),
    .Y(_0045_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2073_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1160_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[7] ),
    .Y(_0216_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2074_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0217_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[6] ),
    .B(_1136_),
    .C(_0212_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2075_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0218_),
    .B(_0217_),
    .A(_0216_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2076_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0217_),
    .A(_0216_),
    .Y(_0219_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2077_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1416_),
    .B(_0218_),
    .C(_0219_),
    .Y(_0220_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2078_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0220_),
    .Y(_0046_));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 _2079_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1350_),
    .Y(_0221_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2080_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0222_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2081_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1185_),
    .A(_0222_),
    .Y(_0223_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2082_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0224_),
    .A(_1160_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2083_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0225_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[7] ),
    .B(_0224_),
    .C(_0219_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2084_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0226_),
    .B(_0225_),
    .A(_0223_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2085_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0225_),
    .A(_0223_),
    .Y(_0227_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2086_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0221_),
    .B(_0226_),
    .C(_0227_),
    .Y(_0228_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2087_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0228_),
    .Y(_0047_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2088_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0229_),
    .B(_1216_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2089_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1216_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[9] ),
    .Y(_0230_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2090_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0231_),
    .B(_0230_),
    .A(_0229_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2091_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0232_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[8] ),
    .B(_1185_),
    .C(_0227_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2092_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0232_),
    .A(_0231_),
    .Y(_0233_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2093_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0234_),
    .C(_0196_),
    .B(_0232_),
    .A(_0231_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2094_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0234_),
    .A(_0233_),
    .Y(_0235_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2095_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0235_),
    .Y(_0048_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2096_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0236_),
    .C(_0232_),
    .B(_1216_),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2097_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0221_),
    .B(_0229_),
    .C(_0236_),
    .Y(_0237_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2098_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0237_),
    .Y(_0049_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2099_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0238_),
    .B(_1292_),
    .A(_1279_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2100_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0050_),
    .B(_0238_),
    .A(_1306_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2101_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0239_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2102_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0240_),
    .B(_0904_),
    .A(\tt_um_rejunity_sn76489.control_noise[0][0] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2103_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0241_),
    .A(\tt_um_rejunity_sn76489.control_noise[0][0] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2104_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0242_),
    .A(\tt_um_rejunity_sn76489.control_noise[0][1] ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2105_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0243_),
    .C(_0242_),
    .B(\tt_um_rejunity_sn76489.noise[0].gen.counter[6] ),
    .A(_0241_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2106_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0244_),
    .B(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .A(\tt_um_rejunity_sn76489.control_noise[0][0] ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2107_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0245_),
    .C(\tt_um_rejunity_sn76489.control_noise[0][1] ),
    .B(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ),
    .A(_0241_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2108_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0240_),
    .B(_0243_),
    .C(_0244_),
    .D(_0245_),
    .Y(_0246_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2109_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0247_),
    .B(_0246_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2110_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0247_),
    .Y(_0248_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2111_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0249_),
    .A(_0915_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2112_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0246_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ),
    .Y(_0250_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2113_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0250_),
    .Y(_0251_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2114_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_sn76489.noise[0].gen.restart_noise ),
    .A(_1264_),
    .Y(_0252_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2115_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0252_),
    .Y(_0253_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2116_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0254_),
    .A(_0249_),
    .B(_0251_),
    .C(_0253_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2117_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0051_),
    .C(_0254_),
    .B(_0248_),
    .A(_0239_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2118_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0251_),
    .Y(_0255_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2119_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0256_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2120_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0247_),
    .Y(_0257_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2121_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0258_),
    .A(_0256_),
    .B(_0257_),
    .C(_0252_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2122_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0052_),
    .C(_0258_),
    .B(_0255_),
    .A(_0239_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2123_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0253_),
    .Y(_0259_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2124_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0247_),
    .Y(_0260_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2125_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0261_),
    .B(_0260_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2126_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0262_),
    .B(_0255_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2127_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0259_),
    .B(_0261_),
    .C(_0262_),
    .Y(_0263_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2128_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0263_),
    .Y(_0053_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2129_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0264_),
    .B(_0260_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2130_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0265_),
    .B(_0255_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2131_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0259_),
    .B(_0264_),
    .C(_0265_),
    .Y(_0266_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2132_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0266_),
    .Y(_0054_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2133_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0250_),
    .Y(_0267_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2134_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0268_),
    .B(_0267_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2135_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0269_),
    .B(_0248_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2136_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0259_),
    .B(_0268_),
    .C(_0269_),
    .Y(_0270_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2137_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0270_),
    .Y(_0055_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2138_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0250_),
    .Y(_0271_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2139_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0272_),
    .B(_0271_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2140_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0273_),
    .B(_0248_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2141_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0259_),
    .B(_0272_),
    .C(_0273_),
    .Y(_0274_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2142_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0274_),
    .Y(_0056_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2143_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0253_),
    .Y(_0275_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2144_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0276_),
    .B(_0271_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2145_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0277_),
    .B(_0248_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2146_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0275_),
    .B(_0276_),
    .C(_0277_),
    .Y(_0278_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2147_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0278_),
    .Y(_0057_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2148_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0279_),
    .B(_0271_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2149_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0257_),
    .Y(_0280_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2150_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0281_),
    .B(_0280_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2151_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0275_),
    .B(_0279_),
    .C(_0281_),
    .Y(_0282_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2152_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0282_),
    .Y(_0058_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2153_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0283_),
    .B(_0260_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2154_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0284_),
    .B(_0267_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2155_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0275_),
    .B(_0283_),
    .C(_0284_),
    .Y(_0285_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2156_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0285_),
    .Y(_0059_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2157_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0286_),
    .B(_0271_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2158_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0287_),
    .B(_0280_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2159_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0275_),
    .B(_0286_),
    .C(_0287_),
    .Y(_0288_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2160_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0288_),
    .Y(_0060_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2161_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0253_),
    .Y(_0289_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2162_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0290_),
    .B(_0251_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2163_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0291_),
    .B(_0280_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2164_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0289_),
    .B(_0290_),
    .C(_0291_),
    .Y(_0292_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2165_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0292_),
    .Y(_0061_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2166_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0293_),
    .B(_0251_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2167_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0294_),
    .B(_0280_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2168_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0289_),
    .B(_0293_),
    .C(_0294_),
    .Y(_0295_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2169_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0295_),
    .Y(_0062_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2170_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0296_),
    .B(_0260_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2171_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0297_),
    .B(_0267_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2172_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0289_),
    .B(_0296_),
    .C(_0297_),
    .Y(_0298_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2173_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0298_),
    .Y(_0063_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2174_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0299_),
    .B(_0257_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2175_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0300_),
    .B(_0267_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2176_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0289_),
    .B(_0299_),
    .C(_0300_),
    .Y(_0301_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2177_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0301_),
    .Y(_0064_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2178_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ),
    .A(\tt_um_rejunity_sn76489.control_noise[0][2] ),
    .Y(_0302_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2179_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0302_),
    .A(_0249_),
    .Y(_0303_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2180_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0304_),
    .A(_0257_),
    .B(_0303_),
    .C(_0252_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2181_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0305_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ),
    .B(_0255_),
    .C(_0304_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2182_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0305_),
    .Y(_0065_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2183_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_sn76489.clk_counter[1] ),
    .A(\tt_um_rejunity_sn76489.clk_counter[0] ),
    .Y(_0306_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2184_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .B(\tt_um_rejunity_sn76489.clk_counter[2] ),
    .C(_0306_),
    .Y(_0307_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2185_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.clk_counter[5] ),
    .B(\tt_um_rejunity_sn76489.clk_counter[4] ),
    .C(\tt_um_rejunity_sn76489.clk_counter[6] ),
    .Y(_0308_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2186_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0308_),
    .A(net1),
    .Y(_0309_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2187_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0307_),
    .A(net1),
    .Y(_0310_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2188_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0311_),
    .A(net2));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2189_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0307_),
    .B(_0309_),
    .C(_0310_),
    .D(_0311_),
    .Y(_0312_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2190_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0312_),
    .Y(_0313_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2191_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0313_),
    .Y(_0314_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2192_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0314_),
    .Y(_0315_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2193_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0316_),
    .B(_0315_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2194_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0312_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ),
    .Y(_0317_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2195_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0221_),
    .B(_0316_),
    .C(_0317_),
    .Y(_0318_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2196_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0318_),
    .Y(_0066_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2197_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0319_),
    .B(_0317_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2198_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0317_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[1] ),
    .Y(_0320_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2199_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0221_),
    .B(_0319_),
    .C(_0320_),
    .Y(_0321_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2200_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0321_),
    .Y(_0067_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2201_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1350_),
    .Y(_0322_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2202_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0323_),
    .B(_0320_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2203_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0320_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[2] ),
    .Y(_0324_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2204_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0322_),
    .B(_0323_),
    .C(_0324_),
    .Y(_0325_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2205_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0325_),
    .Y(_0068_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2206_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0326_),
    .B(_0324_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2207_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0324_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[3] ),
    .Y(_0327_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2208_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0322_),
    .B(_0326_),
    .C(_0327_),
    .Y(_0328_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2209_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0328_),
    .Y(_0069_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2210_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0329_),
    .B(_0327_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2211_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0327_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ),
    .Y(_0330_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2212_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0322_),
    .B(_0329_),
    .C(_0330_),
    .Y(_0331_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2213_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0331_),
    .Y(_0070_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2214_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0332_),
    .B(_0330_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2215_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0330_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .Y(_0333_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2216_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0333_),
    .A(_1223_),
    .Y(_0334_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2217_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0334_),
    .A(_0332_),
    .Y(_0335_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2218_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0335_),
    .Y(_0071_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2219_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0332_),
    .A(\tt_um_rejunity_sn76489.noise[0].gen.counter[6] ),
    .Y(_0336_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2220_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0336_),
    .A(_1224_),
    .Y(_0337_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2221_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0337_),
    .Y(_0072_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2222_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0338_),
    .B(_1059_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2223_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1222_),
    .Y(_0339_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2224_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1059_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[0] ),
    .Y(_0340_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2225_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0340_),
    .A(_0339_),
    .Y(_0341_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2226_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0341_),
    .A(_0338_),
    .Y(_0342_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2227_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0342_),
    .Y(_0073_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2228_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1041_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[1] ),
    .Y(_0343_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2229_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0343_),
    .A(_0338_),
    .Y(_0344_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2230_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0195_),
    .Y(_0345_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2231_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0346_),
    .C(_0345_),
    .B(_0343_),
    .A(_0338_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2232_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0346_),
    .A(_0344_),
    .Y(_0347_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2233_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0347_),
    .Y(_0074_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2234_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1018_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[2] ),
    .Y(_0348_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2235_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0349_),
    .B(_1041_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2236_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0350_),
    .B(_0344_),
    .A(_0349_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2237_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0350_),
    .A(_0348_),
    .Y(_0351_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2238_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0352_),
    .C(_0345_),
    .B(_0350_),
    .A(_0348_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2239_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0352_),
    .A(_0351_),
    .Y(_0353_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2240_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0353_),
    .Y(_0075_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2241_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0354_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2242_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0931_),
    .A(_0354_),
    .Y(_0355_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2243_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0356_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[2] ),
    .B(_1019_),
    .C(_0350_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2244_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0356_),
    .A(_0355_),
    .Y(_0357_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2245_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0358_),
    .C(_0345_),
    .B(_0356_),
    .A(_0355_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2246_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0358_),
    .A(_0357_),
    .Y(_0359_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2247_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0359_),
    .Y(_0076_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2248_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0360_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2249_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1074_),
    .A(_0360_),
    .Y(_0361_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2250_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0362_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[3] ),
    .B(_0931_),
    .C(_0356_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2251_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0362_),
    .A(_0361_),
    .Y(_0363_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2252_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0364_),
    .C(_0345_),
    .B(_0362_),
    .A(_0361_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2253_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0364_),
    .A(_0363_),
    .Y(_0365_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2254_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0365_),
    .Y(_0077_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2255_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0366_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[4] ),
    .B(_1074_),
    .C(_0362_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2256_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0367_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2257_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1104_),
    .A(_0367_),
    .Y(_0368_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2258_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0368_),
    .A(_0366_),
    .Y(_0369_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2259_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0370_),
    .B(_0369_),
    .A(_1401_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2260_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0078_),
    .C(_0370_),
    .B(_0368_),
    .A(_0366_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2261_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0371_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2262_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1126_),
    .A(_0371_),
    .Y(_0372_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2263_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0373_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[5] ),
    .B(_1104_),
    .C(_0366_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2264_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0373_),
    .A(_0372_),
    .Y(_0374_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2265_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0195_),
    .Y(_0375_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2266_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0376_),
    .C(_0375_),
    .B(_0373_),
    .A(_0372_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2267_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0376_),
    .A(_0374_),
    .Y(_0377_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2268_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0377_),
    .Y(_0079_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2269_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0378_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2270_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1152_),
    .A(_0378_),
    .Y(_0379_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2271_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0380_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[6] ),
    .B(_1126_),
    .C(_0373_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2272_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0381_),
    .B(_0380_),
    .A(_0379_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2273_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0380_),
    .A(_0379_),
    .Y(_0382_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2274_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0322_),
    .B(_0381_),
    .C(_0382_),
    .Y(_0383_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2275_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0383_),
    .Y(_0080_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2276_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1178_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[8] ),
    .Y(_0384_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2277_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0385_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[7] ),
    .B(_1152_),
    .C(_0382_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2278_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0385_),
    .A(_0384_),
    .Y(_0386_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2279_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0387_),
    .C(_0375_),
    .B(_0385_),
    .A(_0384_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2280_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0387_),
    .A(_0386_),
    .Y(_0388_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2281_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0388_),
    .Y(_0081_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2282_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0389_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2283_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1197_),
    .A(_0389_),
    .Y(_0390_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2284_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0391_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[8] ),
    .B(_1207_),
    .C(_0385_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2285_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0391_),
    .A(_0390_),
    .Y(_0392_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2286_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0393_),
    .C(_0375_),
    .B(_0391_),
    .A(_0390_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2287_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0393_),
    .A(_0392_),
    .Y(_0394_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2288_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0394_),
    .Y(_0082_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2289_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0395_),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[9] ),
    .B(_1197_),
    .C(_0391_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2290_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0396_),
    .C(_0375_),
    .B(_1198_),
    .A(_0389_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2291_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0396_),
    .A(_0395_),
    .Y(_0397_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2292_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0397_),
    .Y(_0083_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2293_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0313_),
    .Y(_0398_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2294_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0398_),
    .Y(_0399_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2295_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0399_),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ),
    .Y(_0400_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2296_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0401_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2297_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0402_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2298_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0403_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2299_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0404_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2300_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0401_),
    .B(_0402_),
    .C(_0403_),
    .D(_0404_),
    .Y(_0405_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2301_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ),
    .C(_0405_),
    .Y(_0406_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2302_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0407_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ),
    .B(_0406_),
    .C(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2303_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0195_),
    .Y(_0408_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2304_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0409_),
    .C(_0408_),
    .B(_0407_),
    .A(_0315_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2305_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0409_),
    .A(_0400_),
    .Y(_0410_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2306_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0410_),
    .Y(_0084_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2307_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0398_),
    .Y(_0411_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2308_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0411_),
    .Y(_0412_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2309_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0406_),
    .Y(_0413_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2310_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0414_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ),
    .B(_0413_),
    .C(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2311_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0415_),
    .B(_0414_),
    .A(_0407_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2312_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0414_),
    .A(_0407_),
    .Y(_0416_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2313_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0339_),
    .Y(_0417_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2314_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0398_),
    .Y(_0418_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2315_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0418_),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ),
    .Y(_0419_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2316_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0420_),
    .B(_0419_),
    .A(_0417_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2317_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0412_),
    .B(_0415_),
    .C(_0416_),
    .Y(_0085_),
    .D(_0420_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2318_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0421_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ),
    .B(_0413_),
    .C(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2319_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0422_),
    .B(_0421_),
    .A(_0416_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2320_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0421_),
    .A(_0416_),
    .Y(_0423_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2321_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0339_),
    .Y(_0424_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2322_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0418_),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ),
    .Y(_0425_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2323_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0426_),
    .B(_0425_),
    .A(_0424_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2324_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0412_),
    .B(_0422_),
    .C(_0423_),
    .Y(_0086_),
    .D(_0426_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2325_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0314_),
    .Y(_0427_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2326_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0427_),
    .Y(_0428_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2327_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0429_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ),
    .B(_0413_),
    .C(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2328_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0430_),
    .B(_0429_),
    .A(_0423_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2329_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0431_),
    .B(_0429_),
    .A(_0423_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2330_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0431_),
    .Y(_0432_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2331_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0433_),
    .A(_0432_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2332_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0313_),
    .Y(_0434_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2333_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0434_),
    .Y(_0435_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2334_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0435_),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ),
    .Y(_0436_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2335_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0437_),
    .B(_0436_),
    .A(_0424_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2336_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0428_),
    .B(_0430_),
    .C(_0433_),
    .Y(_0087_),
    .D(_0437_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2337_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0413_),
    .Y(_0438_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2338_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0439_),
    .C(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ),
    .B(_0438_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][4] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2339_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0439_),
    .A(_0432_),
    .Y(_0440_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2340_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0441_),
    .B(_0439_),
    .A(_0432_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2341_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0435_),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ),
    .Y(_0442_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2342_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0443_),
    .B(_0442_),
    .A(_0424_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2343_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0428_),
    .B(_0440_),
    .C(_0441_),
    .Y(_0088_),
    .D(_0443_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2344_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0427_),
    .Y(_0444_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2345_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0445_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][5] ),
    .B(_0438_),
    .C(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2346_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0446_),
    .A(_0445_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2347_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0446_),
    .A(_0441_),
    .Y(_0447_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2348_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0398_),
    .Y(_0448_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2349_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0448_),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ),
    .Y(_0449_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2350_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0450_),
    .B(_0449_),
    .A(_1401_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2351_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0089_),
    .C(_0450_),
    .B(_0447_),
    .A(_0444_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2352_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0451_),
    .C(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ),
    .B(_0438_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][6] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2353_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0451_),
    .A(_0432_),
    .B(_0439_),
    .C(_0446_),
    .Y(_0452_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2354_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0431_),
    .B(_0439_),
    .C(_0446_),
    .D(_0451_),
    .Y(_0453_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2355_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0435_),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ),
    .Y(_0454_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2356_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0455_),
    .B(_0454_),
    .A(_0424_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2357_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0428_),
    .B(_0452_),
    .C(_0453_),
    .Y(_0090_),
    .D(_0455_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2358_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0438_),
    .Y(_0456_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2359_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0457_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][7] ),
    .B(_0456_),
    .C(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2360_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0458_),
    .B(_0457_),
    .A(_0453_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2361_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0457_),
    .A(_0453_),
    .Y(_0459_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2362_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1339_),
    .Y(_0460_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2363_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0435_),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ),
    .Y(_0461_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2364_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0462_),
    .B(_0461_),
    .A(_0460_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2365_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0428_),
    .B(_0458_),
    .C(_0459_),
    .Y(_0091_),
    .D(_0462_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2366_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0463_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][8] ),
    .B(_0456_),
    .C(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2367_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0463_),
    .A(_0459_),
    .Y(_0464_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2368_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0465_),
    .B(_0463_),
    .A(_0459_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2369_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0466_),
    .B(_0465_),
    .A(_0464_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2370_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1230_),
    .Y(_0467_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2371_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0448_),
    .A(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ),
    .Y(_0468_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2372_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0469_),
    .B(_0468_),
    .A(_0467_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2373_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0092_),
    .C(_0469_),
    .B(_0466_),
    .A(_0444_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2374_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0314_),
    .Y(_0470_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2375_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0313_),
    .Y(_0471_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2376_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\tt_um_rejunity_sn76489.tone[2].gen.counter[9] ),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][9] ),
    .B(_0471_),
    .C(_0456_),
    .Y(_0472_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2377_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0473_),
    .C(_0472_),
    .B(_0465_),
    .A(_0470_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2378_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1255_),
    .Y(_0474_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2379_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0474_),
    .A(_0411_),
    .B(_0465_),
    .C(_0472_),
    .Y(_0475_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2380_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0093_),
    .B(_0475_),
    .A(_0473_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2381_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0456_),
    .A(_0471_),
    .Y(_0476_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2382_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0476_),
    .A(_0904_),
    .Y(_0477_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2383_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0478_),
    .B(_0477_),
    .A(_0467_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2384_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0094_),
    .C(_0478_),
    .B(_0476_),
    .A(_0904_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2385_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0399_),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ),
    .Y(_0479_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2386_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0480_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2387_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0481_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2388_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0482_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2389_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0483_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2390_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0480_),
    .B(_0481_),
    .C(_0482_),
    .D(_0483_),
    .Y(_0484_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2391_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ),
    .C(_0484_),
    .Y(_0485_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2392_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0486_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ),
    .B(_0485_),
    .C(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2393_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0487_),
    .C(_0408_),
    .B(_0486_),
    .A(_0315_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2394_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0487_),
    .A(_0479_),
    .Y(_0488_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2395_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0488_),
    .Y(_0095_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2396_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0427_),
    .Y(_0489_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2397_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0485_),
    .Y(_0490_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2398_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0491_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ),
    .B(_0490_),
    .C(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2399_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0492_),
    .B(_0491_),
    .A(_0486_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2400_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0491_),
    .A(_0486_),
    .Y(_0493_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2401_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0434_),
    .Y(_0494_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2402_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0494_),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ),
    .Y(_0495_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2403_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0496_),
    .B(_0495_),
    .A(_0460_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2404_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0489_),
    .B(_0492_),
    .C(_0493_),
    .Y(_0096_),
    .D(_0496_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2405_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0497_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ),
    .B(_0490_),
    .C(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2406_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0498_),
    .B(_0497_),
    .A(_0493_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2407_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0497_),
    .A(_0493_),
    .Y(_0499_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2408_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0494_),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ),
    .Y(_0500_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2409_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0501_),
    .B(_0500_),
    .A(_0460_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2410_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0489_),
    .B(_0498_),
    .C(_0499_),
    .Y(_0097_),
    .D(_0501_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2411_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0502_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ),
    .B(_0490_),
    .C(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2412_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0503_),
    .B(_0502_),
    .A(_0499_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2413_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0504_),
    .B(_0502_),
    .A(_0499_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2414_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0504_),
    .Y(_0505_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2415_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0506_),
    .A(_0505_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2416_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0494_),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ),
    .Y(_0507_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2417_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0508_),
    .B(_0507_),
    .A(_0460_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2418_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0489_),
    .B(_0503_),
    .C(_0506_),
    .Y(_0098_),
    .D(_0508_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2419_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0490_),
    .Y(_0509_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2420_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0510_),
    .C(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ),
    .B(_0509_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][4] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2421_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0510_),
    .A(_0505_),
    .Y(_0511_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2422_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0512_),
    .B(_0510_),
    .A(_0505_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2423_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1339_),
    .Y(_0513_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2424_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0494_),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ),
    .Y(_0514_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2425_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0515_),
    .B(_0514_),
    .A(_0513_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2426_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0489_),
    .B(_0511_),
    .C(_0512_),
    .Y(_0099_),
    .D(_0515_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2427_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0516_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][5] ),
    .B(_0509_),
    .C(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2428_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0517_),
    .A(_0516_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2429_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0517_),
    .A(_0512_),
    .Y(_0518_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2430_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0448_),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ),
    .Y(_0519_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2431_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0520_),
    .B(_0519_),
    .A(_0467_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2432_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0100_),
    .C(_0520_),
    .B(_0518_),
    .A(_0444_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2433_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0427_),
    .Y(_0521_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2434_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0522_),
    .C(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ),
    .B(_0509_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][6] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2435_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0522_),
    .A(_0505_),
    .B(_0510_),
    .C(_0517_),
    .Y(_0523_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2436_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0504_),
    .B(_0510_),
    .C(_0517_),
    .D(_0522_),
    .Y(_0524_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2437_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0434_),
    .Y(_0525_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2438_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0525_),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ),
    .Y(_0526_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2439_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0527_),
    .B(_0526_),
    .A(_0513_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2440_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0521_),
    .B(_0523_),
    .C(_0524_),
    .Y(_0101_),
    .D(_0527_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2441_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0509_),
    .Y(_0528_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2442_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0529_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][7] ),
    .B(_0528_),
    .C(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2443_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0530_),
    .B(_0529_),
    .A(_0524_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2444_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0529_),
    .A(_0524_),
    .Y(_0531_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2445_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0525_),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ),
    .Y(_0532_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2446_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0533_),
    .B(_0532_),
    .A(_0513_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2447_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0521_),
    .B(_0530_),
    .C(_0531_),
    .Y(_0102_),
    .D(_0533_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2448_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0534_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][8] ),
    .B(_0528_),
    .C(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2449_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0534_),
    .A(_0531_),
    .Y(_0535_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2450_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0536_),
    .B(_0534_),
    .A(_0531_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2451_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0537_),
    .B(_0536_),
    .A(_0535_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2452_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0448_),
    .A(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ),
    .Y(_0538_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2453_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0539_),
    .B(_0538_),
    .A(_0467_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2454_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0103_),
    .C(_0539_),
    .B(_0537_),
    .A(_0444_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2455_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\tt_um_rejunity_sn76489.tone[1].gen.counter[9] ),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][9] ),
    .B(_0471_),
    .C(_0528_),
    .Y(_0540_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2456_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0541_),
    .C(_0540_),
    .B(_0536_),
    .A(_0470_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2457_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0474_),
    .A(_0399_),
    .B(_0536_),
    .C(_0540_),
    .Y(_0542_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2458_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0104_),
    .B(_0542_),
    .A(_0541_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2459_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0528_),
    .A(_0471_),
    .Y(_0543_));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 _2460_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1230_),
    .Y(_0544_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2461_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0543_),
    .A(_0973_),
    .Y(_0545_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2462_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0546_),
    .B(_0545_),
    .A(_0544_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2463_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0105_),
    .C(_0546_),
    .B(_0543_),
    .A(_0973_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2464_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0399_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ),
    .Y(_0547_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2465_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0548_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2466_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0549_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2467_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0550_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2468_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0551_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2469_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0548_),
    .B(_0549_),
    .C(_0550_),
    .D(_0551_),
    .Y(_0552_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2470_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ),
    .C(_0552_),
    .Y(_0553_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2471_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0554_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][0] ),
    .B(_0553_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2472_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0555_),
    .C(_0408_),
    .B(_0554_),
    .A(_0315_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2473_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0555_),
    .A(_0547_),
    .Y(_0556_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2474_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0556_),
    .Y(_0106_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2475_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0557_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ),
    .B(_0553_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2476_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0558_),
    .B(_0557_),
    .A(_0554_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2477_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0557_),
    .A(_0554_),
    .Y(_0559_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2478_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0525_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ),
    .Y(_0560_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2479_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0561_),
    .B(_0560_),
    .A(_0513_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2480_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0521_),
    .B(_0558_),
    .C(_0559_),
    .Y(_0107_),
    .D(_0561_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2481_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0553_),
    .Y(_0562_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2482_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0563_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][2] ),
    .B(_0562_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2483_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0564_),
    .B(_0563_),
    .A(_0559_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2484_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0563_),
    .A(_0559_),
    .Y(_0565_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2485_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1339_),
    .Y(_0566_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2486_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0525_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ),
    .Y(_0567_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2487_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0568_),
    .B(_0567_),
    .A(_0566_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2488_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0521_),
    .B(_0564_),
    .C(_0565_),
    .Y(_0108_),
    .D(_0568_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2489_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0411_),
    .Y(_0569_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2490_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0570_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][3] ),
    .B(_0562_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2491_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0571_),
    .B(_0570_),
    .A(_0565_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2492_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0572_),
    .B(_0570_),
    .A(_0565_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2493_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0572_),
    .Y(_0573_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2494_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0574_),
    .A(_0573_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2495_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0434_),
    .Y(_0575_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2496_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0575_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ),
    .Y(_0576_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2497_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0577_),
    .B(_0576_),
    .A(_0566_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2498_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0569_),
    .B(_0571_),
    .C(_0574_),
    .Y(_0109_),
    .D(_0577_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2499_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0562_),
    .Y(_0578_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2500_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0579_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ),
    .B(_0578_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][4] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2501_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0579_),
    .A(_0573_),
    .Y(_0580_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2502_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0581_),
    .B(_0579_),
    .A(_0573_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2503_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0575_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ),
    .Y(_0582_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2504_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0583_),
    .B(_0582_),
    .A(_0566_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2505_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0569_),
    .B(_0580_),
    .C(_0581_),
    .Y(_0110_),
    .D(_0583_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2506_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0584_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][5] ),
    .B(_0562_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2507_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0585_),
    .A(_0584_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2508_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0585_),
    .A(_0581_),
    .Y(_0586_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2509_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0418_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ),
    .Y(_0587_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2510_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0588_),
    .B(_0587_),
    .A(_0544_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2511_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0111_),
    .C(_0588_),
    .B(_0586_),
    .A(_0412_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2512_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0589_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ),
    .B(_0578_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][6] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2513_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0589_),
    .A(_0573_),
    .B(_0579_),
    .C(_0585_),
    .Y(_0590_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2514_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0572_),
    .B(_0579_),
    .C(_0585_),
    .D(_0589_),
    .Y(_0591_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2515_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0575_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ),
    .Y(_0592_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2516_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0593_),
    .B(_0592_),
    .A(_0566_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2517_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0569_),
    .B(_0590_),
    .C(_0591_),
    .Y(_0112_),
    .D(_0593_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2518_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0594_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][7] ),
    .B(_0578_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2519_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0595_),
    .B(_0594_),
    .A(_0591_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2520_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0594_),
    .A(_0591_),
    .Y(_0596_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2521_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0575_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ),
    .Y(_0597_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2522_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0598_),
    .B(_0597_),
    .A(_1340_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2523_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0569_),
    .B(_0595_),
    .C(_0596_),
    .Y(_0113_),
    .D(_0598_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2524_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0578_),
    .Y(_0599_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2525_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0600_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][8] ),
    .B(_0599_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2526_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0601_),
    .B(_0600_),
    .A(_0596_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2527_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0600_),
    .A(_0596_),
    .Y(_0602_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2528_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0314_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ),
    .Y(_0603_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2529_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0604_),
    .B(_0603_),
    .A(_1340_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _2530_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0470_),
    .B(_0601_),
    .C(_0602_),
    .Y(_0114_),
    .D(_0604_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2531_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0605_),
    .C(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ),
    .B(_0599_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][9] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2532_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0605_),
    .A(_0602_),
    .Y(_0606_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2533_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0418_),
    .A(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ),
    .Y(_0607_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2534_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0608_),
    .B(_0607_),
    .A(_0544_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2535_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0115_),
    .C(_0608_),
    .B(_0606_),
    .A(_0412_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2536_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0609_),
    .C(_0936_),
    .B(_0599_),
    .A(_0470_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2537_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0474_),
    .A(_0936_),
    .B(_0411_),
    .C(_0599_),
    .Y(_0610_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2538_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0116_),
    .B(_0610_),
    .A(_0609_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2539_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1305_),
    .Y(_0611_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2540_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1064_),
    .A(_1059_),
    .Y(_0612_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2541_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0612_),
    .A(_1067_),
    .Y(_0613_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2542_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0614_),
    .B(_0613_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2543_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0613_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[0] ),
    .Y(_0615_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2544_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0611_),
    .B(_0614_),
    .C(_0615_),
    .Y(_0616_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2545_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0616_),
    .Y(_0117_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2546_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0617_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[1] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2547_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1068_),
    .A(_1069_),
    .Y(_0618_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2548_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0618_),
    .A(_0617_),
    .Y(_0619_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2549_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0619_),
    .A(_0615_),
    .Y(_0620_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2550_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0621_),
    .C(_0408_),
    .B(_0619_),
    .A(_0615_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2551_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0621_),
    .A(_0620_),
    .Y(_0622_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2552_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0622_),
    .Y(_0118_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2553_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0623_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _2554_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0624_),
    .B(_1068_),
    .A(_1069_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2555_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1053_),
    .A(_1048_),
    .Y(_0625_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2556_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0625_),
    .A(_1036_),
    .Y(_0626_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2557_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0626_),
    .A(_0624_),
    .Y(_0627_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2558_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0627_),
    .A(_0623_),
    .Y(_0628_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2559_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0629_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[1] ),
    .B(_0615_),
    .C(_0618_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2560_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0629_),
    .A(_0628_),
    .Y(_0630_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2561_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1349_),
    .Y(_0631_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2562_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0632_),
    .C(_0631_),
    .B(_0629_),
    .A(_0628_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2563_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0632_),
    .A(_0630_),
    .Y(_0633_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2564_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0633_),
    .Y(_0119_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2565_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0634_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2566_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1033_),
    .A(_1009_),
    .Y(_0635_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2567_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0635_),
    .A(_1071_),
    .Y(_0636_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2568_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0636_),
    .A(_0634_),
    .Y(_0637_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2569_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0638_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[2] ),
    .B(_0627_),
    .C(_0629_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2570_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0638_),
    .A(_0637_),
    .Y(_0639_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2571_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0640_),
    .C(_0631_),
    .B(_0638_),
    .A(_0637_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2572_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0640_),
    .A(_0639_),
    .Y(_0641_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2573_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0641_),
    .Y(_0120_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2574_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0642_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2575_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net18),
    .A(_0642_),
    .Y(_0643_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2576_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0644_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[3] ),
    .B(_0636_),
    .C(_0638_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2577_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0644_),
    .A(_0643_),
    .Y(_0645_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2578_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0646_),
    .C(_0631_),
    .B(_0644_),
    .A(_0643_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2579_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0646_),
    .A(_0645_),
    .Y(_0647_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2580_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0647_),
    .Y(_0121_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2581_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0648_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2582_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net19),
    .A(_0648_),
    .Y(_0649_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2583_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0650_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[4] ),
    .B(net18),
    .C(_0644_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2584_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0650_),
    .A(_0649_),
    .Y(_0651_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2585_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0652_),
    .C(_0631_),
    .B(_0650_),
    .A(_0649_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2586_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0652_),
    .A(_0651_),
    .Y(_0653_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2587_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0653_),
    .Y(_0122_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2588_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0654_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2589_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net20),
    .A(_0654_),
    .Y(_0655_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2590_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0656_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[5] ),
    .B(net19),
    .C(_0650_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2591_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0656_),
    .A(_0655_),
    .Y(_0657_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2592_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1349_),
    .Y(_0658_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2593_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0659_),
    .C(_0658_),
    .B(_0656_),
    .A(_0655_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2594_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0659_),
    .A(_0657_),
    .Y(_0660_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2595_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0660_),
    .Y(_0123_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2596_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0661_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2597_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net21),
    .A(_0661_),
    .Y(_0662_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2598_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0663_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[6] ),
    .B(net20),
    .C(_0656_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2599_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0663_),
    .A(_0662_),
    .Y(_0664_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2600_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0665_),
    .C(_0658_),
    .B(_0663_),
    .A(_0662_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2601_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0665_),
    .A(_0664_),
    .Y(_0666_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2602_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0666_),
    .Y(_0124_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2603_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0667_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2604_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net22),
    .A(_0667_),
    .Y(_0668_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2605_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0669_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[7] ),
    .B(net21),
    .C(_0663_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2606_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0669_),
    .A(_0668_),
    .Y(_0670_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2607_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0671_),
    .C(_0658_),
    .B(_0669_),
    .A(_0668_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2608_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0671_),
    .A(_0670_),
    .Y(_0672_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2609_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0672_),
    .Y(_0125_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2610_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0673_),
    .B(net23),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2611_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net23),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[9] ),
    .Y(_0674_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2612_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0675_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[8] ),
    .B(net22),
    .C(_0669_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2613_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0676_),
    .C(_0675_),
    .B(_0674_),
    .A(_0673_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2614_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0474_),
    .A(_0675_),
    .B(_0673_),
    .C(_0674_),
    .Y(_0677_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2615_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0126_),
    .B(_0677_),
    .A(_0676_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2616_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0678_),
    .B(_0674_),
    .A(_0675_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2617_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net24),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[10] ),
    .Y(_0679_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2618_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0680_),
    .C(_0679_),
    .B(_0678_),
    .A(_0673_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2619_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1255_),
    .Y(_0681_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2620_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0681_),
    .A(_0673_),
    .B(_0678_),
    .C(_0679_),
    .Y(_0682_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2621_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0127_),
    .B(_0682_),
    .A(_0680_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2622_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0683_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[11] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2623_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net25),
    .A(_0683_),
    .Y(_0684_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2624_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0685_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[9] ),
    .B(_1210_),
    .C(_0675_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2625_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0686_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[10] ),
    .B(net24),
    .C(_0685_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2626_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0686_),
    .A(_0684_),
    .Y(_0687_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2627_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0688_),
    .C(_0658_),
    .B(_0686_),
    .A(_0684_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2628_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0688_),
    .A(_0687_),
    .Y(_0689_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2629_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0689_),
    .Y(_0128_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _2630_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0690_),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[11] ),
    .B(net25),
    .C(_0686_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2631_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0690_),
    .A(_1224_),
    .Y(_0691_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2632_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0691_),
    .Y(_0129_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2633_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1225_),
    .Y(_0692_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2634_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0692_),
    .Y(_0693_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2635_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0130_),
    .B(_0693_),
    .A(_1224_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _2636_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0694_),
    .B(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[11] ),
    .A(_1228_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2637_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0695_),
    .B(_1228_),
    .A(\tt_um_rejunity_sn76489.DAC_dat ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2638_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0611_),
    .B(_0694_),
    .C(_0695_),
    .Y(_0696_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2639_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0696_),
    .Y(_0131_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2640_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_1232_),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[0] ),
    .Y(_0697_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2641_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0697_),
    .Y(_0698_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2642_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0698_),
    .A(_1222_),
    .Y(_0699_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2643_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0699_),
    .Y(_0144_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2644_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0144_),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[0] ),
    .Y(_0700_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2645_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0700_),
    .A(_1231_),
    .B(_0693_),
    .C(_0613_),
    .Y(_0701_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2646_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0701_),
    .Y(_0132_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2647_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1231_),
    .Y(_0702_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2648_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1227_),
    .Y(_0703_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2649_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0698_),
    .Y(_0704_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2650_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[0] ),
    .B(_0703_),
    .C(_0704_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[1] ),
    .Y(_0705_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2651_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0706_),
    .A(_0693_),
    .B(_0618_),
    .C(_0705_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2652_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0706_),
    .A(_0702_),
    .Y(_0707_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2653_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0707_),
    .Y(_0133_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2654_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[1] ),
    .B(_0703_),
    .C(_0704_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[2] ),
    .Y(_0708_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2655_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0709_),
    .A(_0693_),
    .B(_0627_),
    .C(_0708_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2656_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0709_),
    .A(_0702_),
    .Y(_0710_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2657_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0710_),
    .Y(_0134_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2658_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0692_),
    .Y(_0711_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2659_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[2] ),
    .B(_0703_),
    .C(_0704_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[3] ),
    .Y(_0712_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2660_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0713_),
    .A(_0711_),
    .B(_0636_),
    .C(_0712_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2661_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0713_),
    .A(_0702_),
    .Y(_0714_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2662_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0714_),
    .Y(_0135_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2663_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0692_),
    .Y(_0715_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2664_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[3] ),
    .B(_1227_),
    .C(_0698_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[4] ),
    .Y(_0716_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2665_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0716_),
    .A(_1095_),
    .B(_1096_),
    .C(_0715_),
    .Y(_0717_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2666_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0717_),
    .A(_0702_),
    .Y(_0718_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2667_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0718_),
    .Y(_0136_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2668_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1223_),
    .Y(_0719_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2669_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[4] ),
    .B(_0703_),
    .C(_0704_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[5] ),
    .Y(_0720_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2670_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0721_),
    .A(net19),
    .B(_0711_),
    .C(_0720_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2671_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0721_),
    .A(_0719_),
    .Y(_0722_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2672_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0722_),
    .Y(_0137_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2673_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1226_),
    .Y(_0723_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2674_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0697_),
    .Y(_0724_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2675_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[5] ),
    .B(_0723_),
    .C(_0724_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[6] ),
    .Y(_0725_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2676_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0726_),
    .A(net20),
    .B(_0711_),
    .C(_0725_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2677_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0726_),
    .A(_0719_),
    .Y(_0727_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2678_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0727_),
    .Y(_0138_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2679_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[6] ),
    .B(_1227_),
    .C(_0698_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[7] ),
    .Y(_0728_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2680_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0728_),
    .A(_1173_),
    .B(_1174_),
    .C(_0715_),
    .Y(_0729_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2681_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0729_),
    .A(_0719_),
    .Y(_0730_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2682_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0730_),
    .Y(_0139_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2683_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[7] ),
    .B(_0723_),
    .C(_0724_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[8] ),
    .Y(_0731_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2684_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0732_),
    .A(net22),
    .B(_0711_),
    .C(_0731_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2685_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0732_),
    .A(_0719_),
    .Y(_0733_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2686_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0733_),
    .Y(_0140_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2687_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[8] ),
    .B(_0723_),
    .C(_0724_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[9] ),
    .Y(_0734_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2688_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0735_),
    .A(net23),
    .B(_0715_),
    .C(_0734_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2689_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0735_),
    .A(_0417_),
    .Y(_0736_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2690_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0736_),
    .Y(_0141_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2691_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[9] ),
    .B(_0723_),
    .C(_0724_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[10] ),
    .Y(_0737_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2692_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0738_),
    .A(net24),
    .B(_0715_),
    .C(_0737_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2693_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0738_),
    .A(_0417_),
    .Y(_0739_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2694_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0739_),
    .Y(_0142_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2695_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net25),
    .B(_0692_),
    .C(_1228_),
    .D(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[10] ),
    .Y(_0740_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2696_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[11] ),
    .B(_0144_),
    .C(_0740_),
    .D(_1231_),
    .Y(_0741_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2697_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0741_),
    .Y(_0143_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2698_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0145_),
    .B(_0246_),
    .A(_1306_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2699_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0742_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][4] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2700_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0743_),
    .A(\tt_um_rejunity_sn76489.latch_control_reg[2] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2701_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0744_),
    .B(net10),
    .A(_0743_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2702_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0744_),
    .Y(_0745_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2703_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.latch_control_reg[1] ),
    .Y(_0746_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2704_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.latch_control_reg[0] ),
    .Y(_0747_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2705_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0746_),
    .B(_0747_),
    .C(net9),
    .Y(_0748_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2706_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0748_),
    .Y(_0749_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2707_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0750_),
    .B(_0749_),
    .A(_0745_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2708_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0750_),
    .Y(_0751_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2709_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0752_),
    .A(_1294_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2710_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0745_),
    .Y(_0753_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2711_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0749_),
    .Y(_0754_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2712_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1299_),
    .A(_0752_),
    .B(_0753_),
    .C(_0754_),
    .Y(_0755_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2713_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0146_),
    .C(_0755_),
    .B(_0751_),
    .A(_0742_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2714_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0756_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][5] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2715_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1313_),
    .Y(_0757_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2716_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0757_),
    .A(_1260_),
    .B(_0753_),
    .C(_0754_),
    .Y(_0758_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2717_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0147_),
    .C(_0758_),
    .B(_0751_),
    .A(_0756_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2718_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0759_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][6] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2719_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0757_),
    .A(_1269_),
    .B(_0753_),
    .C(_0754_),
    .Y(_0760_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2720_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0148_),
    .C(_0760_),
    .B(_0751_),
    .A(_0759_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2721_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0761_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][7] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2722_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0757_),
    .A(_1273_),
    .B(_0753_),
    .C(_0754_),
    .Y(_0762_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2723_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0149_),
    .C(_0762_),
    .B(_0751_),
    .A(_0761_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2724_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0763_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][8] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2725_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1277_),
    .Y(_0764_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2726_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0748_),
    .Y(_0765_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2727_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0757_),
    .A(_0764_),
    .B(_0745_),
    .C(_0765_),
    .Y(_0766_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2728_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0150_),
    .C(_0766_),
    .B(_0750_),
    .A(_0763_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2729_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0767_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[2][9] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2730_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0768_),
    .A(net7));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2731_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0768_),
    .Y(_0769_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2732_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1313_),
    .Y(_0770_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2733_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0770_),
    .A(_0769_),
    .B(_0745_),
    .C(_0765_),
    .Y(_0771_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2734_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0151_),
    .C(_0771_),
    .B(_0750_),
    .A(_0767_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2735_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0772_),
    .A(\tt_um_rejunity_sn76489.latch_control_reg[1] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2736_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net9),
    .Y(_0773_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2737_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0774_),
    .A(_0747_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2738_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0775_),
    .B(net10),
    .A(\tt_um_rejunity_sn76489.latch_control_reg[2] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2739_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0775_),
    .Y(_0776_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2740_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0777_),
    .B(_0776_),
    .A(_0774_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2741_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0772_),
    .B(_0773_),
    .C(_0777_),
    .Y(_0778_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2742_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0778_),
    .Y(_0779_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2743_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0780_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][4] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2744_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1243_),
    .Y(_0781_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _2745_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0746_),
    .B(_0774_),
    .C(_0781_),
    .D(_0776_),
    .Y(_0782_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2746_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0782_),
    .Y(_0783_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2747_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0784_),
    .A(_0780_),
    .B(_0783_),
    .C(_1305_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2748_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0152_),
    .C(_0784_),
    .B(_0779_),
    .A(_0752_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2749_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0785_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][5] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2750_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0786_),
    .A(_0785_),
    .B(_0783_),
    .C(_1305_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2751_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0153_),
    .C(_0786_),
    .B(_0779_),
    .A(_1261_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2752_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0787_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][6] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2753_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1349_),
    .Y(_0788_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2754_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0789_),
    .A(_0787_),
    .B(_0783_),
    .C(_0788_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2755_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0154_),
    .C(_0789_),
    .B(_0779_),
    .A(_1270_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2756_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0790_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][7] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2757_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0791_),
    .A(_0790_),
    .B(_0783_),
    .C(_0788_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2758_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0155_),
    .C(_0791_),
    .B(_0779_),
    .A(_1274_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2759_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0792_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][8] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2760_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0793_),
    .A(_0792_),
    .B(_0782_),
    .C(_0788_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2761_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0156_),
    .C(_0793_),
    .B(_0778_),
    .A(_0764_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2762_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0794_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[1][9] ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2763_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0795_),
    .A(_0794_),
    .B(_0782_),
    .C(_0788_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2764_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0157_),
    .C(_0795_),
    .B(_0778_),
    .A(_0769_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2765_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0796_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][4] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2766_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0776_),
    .Y(_0797_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2767_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0798_),
    .B(_0797_),
    .A(_0749_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2768_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0798_),
    .Y(_0799_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2769_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0797_),
    .Y(_0800_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2770_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0770_),
    .A(_0752_),
    .B(_0765_),
    .C(_0800_),
    .Y(_0801_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2771_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0158_),
    .C(_0801_),
    .B(_0799_),
    .A(_0796_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2772_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0802_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][5] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2773_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0770_),
    .A(_1260_),
    .B(_0765_),
    .C(_0800_),
    .Y(_0803_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2774_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0159_),
    .C(_0803_),
    .B(_0799_),
    .A(_0802_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2775_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0804_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][6] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2776_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0749_),
    .Y(_0805_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2777_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0770_),
    .A(_1269_),
    .B(_0805_),
    .C(_0800_),
    .Y(_0806_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2778_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0160_),
    .C(_0806_),
    .B(_0799_),
    .A(_0804_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2779_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0807_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][7] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2780_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1313_),
    .Y(_0808_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2781_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0808_),
    .A(_1273_),
    .B(_0805_),
    .C(_0800_),
    .Y(_0809_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2782_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0161_),
    .C(_0809_),
    .B(_0799_),
    .A(_0807_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2783_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0810_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][8] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2784_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0808_),
    .A(_0764_),
    .B(_0805_),
    .C(_0797_),
    .Y(_0811_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2785_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0162_),
    .C(_0811_),
    .B(_0798_),
    .A(_0810_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _2786_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0812_),
    .A(\tt_um_rejunity_sn76489.control_tone_freq[0][9] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2787_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0808_),
    .A(_0769_),
    .B(_0805_),
    .C(_0797_),
    .Y(_0813_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2788_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0163_),
    .C(_0813_),
    .B(_0798_),
    .A(_0812_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2789_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0781_),
    .A(net8),
    .B(_1247_),
    .C(_1248_),
    .Y(_0814_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2790_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0814_),
    .Y(_0815_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2791_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1290_),
    .A(_0746_),
    .B(\tt_um_rejunity_sn76489.latch_control_reg[0] ),
    .C(_0744_),
    .Y(_0816_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2792_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0816_),
    .Y(_0817_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2793_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0818_),
    .B(_0817_),
    .A(_0815_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2794_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1320_),
    .Y(_0819_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2795_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0819_),
    .A(_1294_),
    .B(_0815_),
    .C(_0817_),
    .Y(_0820_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2796_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0821_),
    .A(_1037_),
    .B(_0818_),
    .C(_0820_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2797_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0821_),
    .Y(_0164_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2798_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net3),
    .Y(_0822_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2799_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0819_),
    .A(_0822_),
    .B(_0815_),
    .C(_0817_),
    .Y(_0823_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2800_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0824_),
    .A(_0919_),
    .B(_0818_),
    .C(_0823_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2801_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0824_),
    .Y(_0165_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2802_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net4),
    .Y(_0825_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2803_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0819_),
    .A(_0825_),
    .B(_0815_),
    .C(_0817_),
    .Y(_0826_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2804_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0827_),
    .A(_1013_),
    .B(_0818_),
    .C(_0826_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2805_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0827_),
    .Y(_0166_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2806_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net5),
    .Y(_0828_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2807_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0819_),
    .A(_0828_),
    .B(_0814_),
    .C(_0816_),
    .Y(_0829_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2808_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0830_),
    .A(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ),
    .B(_0818_),
    .C(_0829_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2809_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0830_),
    .Y(_0167_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _2810_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net8),
    .B(_0768_),
    .C(_1248_),
    .Y(_0831_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _2811_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0772_),
    .B(_0747_),
    .C(_0744_),
    .Y(_0832_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2812_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0781_),
    .A(net10),
    .Y(_0833_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2813_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0833_),
    .Y(_0834_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_4 _2814_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0835_),
    .A(_0773_),
    .B(_0831_),
    .C(_0832_),
    .D(_0834_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2815_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0773_),
    .B(_0831_),
    .C(_0832_),
    .D(_0833_),
    .Y(_0836_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2816_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0837_),
    .A(_1024_),
    .B(_0836_),
    .C(_0681_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2817_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0838_),
    .A(_1252_),
    .B(_0835_),
    .C(_0837_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2818_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0838_),
    .Y(_0168_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2819_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0839_),
    .A(_0896_),
    .B(_0836_),
    .C(_0681_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2820_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0840_),
    .A(_0822_),
    .B(_0835_),
    .C(_0839_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2821_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0840_),
    .Y(_0169_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2822_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0841_),
    .A(_0903_),
    .B(_0836_),
    .C(_0681_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2823_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0842_),
    .A(_0825_),
    .B(_0835_),
    .C(_0841_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2824_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0842_),
    .Y(_0170_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2825_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1255_),
    .Y(_0843_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2826_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0844_),
    .A(_0913_),
    .B(_0836_),
    .C(_0843_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2827_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0845_),
    .A(_0828_),
    .B(_0835_),
    .C(_0844_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2828_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0845_),
    .Y(_0171_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2829_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0781_),
    .A(_1242_),
    .B(_1247_),
    .C(net6),
    .Y(_0846_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2830_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0846_),
    .Y(_0847_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2831_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1244_),
    .A(_0746_),
    .B(\tt_um_rejunity_sn76489.latch_control_reg[0] ),
    .C(_0775_),
    .Y(_0848_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2832_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0848_),
    .Y(_0849_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2833_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0850_),
    .B(_0849_),
    .A(_0847_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2834_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1320_),
    .Y(_0851_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2835_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0851_),
    .A(_1294_),
    .B(_0847_),
    .C(_0849_),
    .Y(_0852_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2836_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0853_),
    .A(_0958_),
    .B(_0850_),
    .C(_0852_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2837_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0853_),
    .Y(_0172_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2838_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0851_),
    .A(_0822_),
    .B(_0847_),
    .C(_0849_),
    .Y(_0854_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2839_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0855_),
    .A(_0992_),
    .B(_0850_),
    .C(_0854_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2840_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0855_),
    .Y(_0173_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2841_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0851_),
    .A(_0825_),
    .B(_0847_),
    .C(_0849_),
    .Y(_0856_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2842_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0857_),
    .A(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .B(_0850_),
    .C(_0856_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2843_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0857_),
    .Y(_0174_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2844_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0851_),
    .A(_0828_),
    .B(_0846_),
    .C(_0848_),
    .Y(_0858_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2845_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0859_),
    .A(_0994_),
    .B(_0850_),
    .C(_0858_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2846_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0859_),
    .Y(_0175_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _2847_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1242_),
    .B(_0768_),
    .C(_1248_),
    .Y(_0860_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _2848_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0772_),
    .B(_0747_),
    .C(_0776_),
    .Y(_0861_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_4 _2849_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0862_),
    .A(_0773_),
    .B(_0860_),
    .C(_0861_),
    .D(_0833_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _2850_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net9),
    .B(_0860_),
    .C(_0861_),
    .D(_0833_),
    .Y(_0863_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2851_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0864_),
    .A(_0942_),
    .B(_0863_),
    .C(_0843_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2852_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0865_),
    .A(_1252_),
    .B(_0862_),
    .C(_0864_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2853_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0865_),
    .Y(_0176_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2854_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0866_),
    .A(_0944_),
    .B(_0863_),
    .C(_0843_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2855_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0867_),
    .A(_0822_),
    .B(_0862_),
    .C(_0866_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2856_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0867_),
    .Y(_0177_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2857_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0868_),
    .A(_0934_),
    .B(_0863_),
    .C(_0843_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2858_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0869_),
    .A(_0825_),
    .B(_0862_),
    .C(_0868_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2859_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0869_),
    .Y(_0178_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2860_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0870_),
    .A(_0999_),
    .B(_0863_),
    .C(_1256_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2861_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0871_),
    .A(_0828_),
    .B(_0862_),
    .C(_0870_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2862_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0871_),
    .Y(_0179_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2863_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0180_),
    .B(_1306_),
    .A(\tt_um_rejunity_sn76489.clk_counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2864_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\tt_um_rejunity_sn76489.clk_counter[1] ),
    .A(\tt_um_rejunity_sn76489.clk_counter[0] ),
    .Y(_0872_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2865_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0873_),
    .B(_0306_),
    .A(_0544_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2866_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0181_),
    .B(_0873_),
    .A(_0872_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2867_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0874_),
    .B(_0872_),
    .A(\tt_um_rejunity_sn76489.clk_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2868_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0872_),
    .A(\tt_um_rejunity_sn76489.clk_counter[2] ),
    .Y(_0875_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2869_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0611_),
    .B(_0874_),
    .C(_0875_),
    .Y(_0876_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2870_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0876_),
    .Y(_0182_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2871_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0877_),
    .B(_0875_),
    .A(\tt_um_rejunity_sn76489.clk_counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2872_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0875_),
    .A(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .Y(_0878_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2873_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0611_),
    .B(_0877_),
    .C(_0878_),
    .Y(_0879_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2874_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0879_),
    .Y(_0183_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2875_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0880_),
    .B(_0878_),
    .A(\tt_um_rejunity_sn76489.clk_counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2876_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0878_),
    .A(\tt_um_rejunity_sn76489.clk_counter[4] ),
    .Y(_0881_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _2877_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_1322_),
    .B(_0880_),
    .C(_0881_),
    .Y(_0882_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2878_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0882_),
    .Y(_0184_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _2879_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0883_),
    .B(_0881_),
    .A(\tt_um_rejunity_sn76489.clk_counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _2880_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0881_),
    .A(\tt_um_rejunity_sn76489.clk_counter[5] ),
    .Y(_0884_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2881_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0884_),
    .A(_0339_),
    .Y(_0885_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2882_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0885_),
    .A(_0883_),
    .Y(_0886_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2883_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0886_),
    .Y(_0185_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _2884_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0883_),
    .A(\tt_um_rejunity_sn76489.clk_counter[6] ),
    .Y(_0887_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _2885_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_0887_),
    .A(_0417_),
    .Y(_0888_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2886_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0888_),
    .Y(_0186_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2887_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0889_),
    .A(_0764_),
    .B(_1290_),
    .C(_1266_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2888_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0187_),
    .C(_0889_),
    .B(_0834_),
    .A(_0774_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2889_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0890_),
    .A(_0772_),
    .B(_0834_),
    .C(_1266_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2890_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0188_),
    .C(_0890_),
    .B(_1290_),
    .A(_0769_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2891_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0891_),
    .A(_0743_),
    .B(_0834_),
    .C(_1314_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _2892_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0189_),
    .B(_0891_),
    .A(_1262_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2893_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_0808_),
    .A(_0752_),
    .B(_1284_),
    .C(_1298_),
    .Y(_0892_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2894_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0190_),
    .C(_0892_),
    .B(_0238_),
    .A(_0241_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2895_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1314_),
    .A(_1260_),
    .B(_1279_),
    .C(_1292_),
    .Y(_0893_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _2896_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0191_),
    .C(_0893_),
    .B(_0238_),
    .A(_0242_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _2897_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_1321_),
    .A(net4),
    .B(_1278_),
    .C(_1291_),
    .Y(_0894_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _2898_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_0895_),
    .A(\tt_um_rejunity_sn76489.control_noise[0][2] ),
    .B(_0238_),
    .C(_0894_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _2899_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_0895_),
    .Y(_0192_));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2900_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0000_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2901_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0001_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2902_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0002_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2903_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0003_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2904_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0004_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2905_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0005_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2906_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0006_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2907_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0007_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2908_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0008_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2909_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0009_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2910_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0010_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2911_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0011_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2912_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0012_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2913_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0013_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2914_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0014_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2915_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0015_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2916_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0016_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2917_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0017_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2918_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0018_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2919_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0019_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2920_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0020_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2921_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_12_0_wb_clk_i),
    .D(_0021_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2922_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_6_0_wb_clk_i),
    .D(_0022_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2923_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0023_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2924_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0024_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2925_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0025_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2926_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_12_0_wb_clk_i),
    .D(_0026_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2927_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0027_),
    .Q(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2928_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_4_0_wb_clk_i),
    .D(_0028_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2929_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_4_0_wb_clk_i),
    .D(_0029_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2930_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_4_0_wb_clk_i),
    .D(_0030_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2931_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_4_0_wb_clk_i),
    .D(_0031_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2932_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0032_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2933_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0033_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2934_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0034_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2935_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0035_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2936_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_4_0_wb_clk_i),
    .D(_0036_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2937_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_4_0_wb_clk_i),
    .D(_0037_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2938_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0038_),
    .Q(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2939_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_4_0_wb_clk_i),
    .D(_0039_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2940_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_4_0_wb_clk_i),
    .D(_0040_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2941_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0041_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2942_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0042_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2943_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0043_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2944_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0044_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2945_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0045_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2946_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0046_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2947_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0047_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2948_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0048_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2949_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0049_),
    .Q(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2950_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_3_0_wb_clk_i),
    .D(_0050_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.restart_noise ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2951_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_3_0_wb_clk_i),
    .D(_0051_),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2952_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0052_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2953_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0053_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2954_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0054_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2955_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0055_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2956_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0056_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2957_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0057_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2958_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0058_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2959_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0059_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2960_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0060_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2961_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0061_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2962_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0062_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2963_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0063_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2964_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0064_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2965_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0065_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2966_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0066_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2967_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0067_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2968_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0068_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2969_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0069_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2970_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0070_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2971_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0071_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2972_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0072_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2973_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0073_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2974_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_6_0_wb_clk_i),
    .D(_0074_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2975_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_6_0_wb_clk_i),
    .D(_0075_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2976_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_6_0_wb_clk_i),
    .D(_0076_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2977_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_5_0_wb_clk_i),
    .D(_0077_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2978_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_6_0_wb_clk_i),
    .D(_0078_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2979_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0079_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2980_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0080_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2981_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0081_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2982_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0082_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2983_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_7_0_wb_clk_i),
    .D(_0083_),
    .Q(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2984_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0084_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2985_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0085_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2986_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0086_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2987_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0087_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2988_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0088_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2989_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0089_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2990_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0090_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2991_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0091_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2992_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0092_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2993_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0093_),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2994_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0094_),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2995_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0095_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2996_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0096_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2997_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0097_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2998_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0098_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _2999_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0099_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3000_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0100_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3001_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0101_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3002_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0102_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3003_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0103_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3004_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0104_),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3005_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0105_),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3006_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0106_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3007_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0107_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3008_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0108_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3009_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0109_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3010_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0110_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3011_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0111_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3012_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0112_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3013_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0113_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3014_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0114_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3015_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0115_),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3016_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0116_),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.in ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3017_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0117_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3018_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0118_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3019_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_12_0_wb_clk_i),
    .D(_0119_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3020_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_12_0_wb_clk_i),
    .D(_0120_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3021_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_12_0_wb_clk_i),
    .D(_0121_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3022_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_12_0_wb_clk_i),
    .D(_0122_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3023_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_12_0_wb_clk_i),
    .D(_0123_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3024_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0124_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3025_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0125_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3026_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0126_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3027_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0127_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3028_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0128_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3029_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0129_),
    .Q(\tt_um_rejunity_sn76489.pwm.accumulator[12] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3030_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_12_0_wb_clk_i),
    .D(_0130_),
    .Q(\tt_um_rejunity_sn76489.DAC_le ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3031_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0131_),
    .Q(\tt_um_rejunity_sn76489.DAC_dat ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3032_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0132_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3033_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0133_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3034_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0134_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3035_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0135_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3036_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0136_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3037_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0137_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3038_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0138_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3039_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0139_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3040_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0140_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3041_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_13_0_wb_clk_i),
    .D(_0141_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3042_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0142_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3043_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0143_),
    .Q(\tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3044_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_15_0_wb_clk_i),
    .D(_0144_),
    .Q(\tt_um_rejunity_sn76489.DAC_clk ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3045_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0145_),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3046_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_10_0_wb_clk_i),
    .D(_0146_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3047_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0147_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3048_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0148_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3049_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0149_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3050_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0150_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3051_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0151_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3052_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0152_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3053_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0153_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3054_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0154_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3055_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0155_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3056_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0156_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3057_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_8_0_wb_clk_i),
    .D(_0157_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3058_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0158_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3059_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0159_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3060_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0160_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3061_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_2_0_wb_clk_i),
    .D(_0161_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3062_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0162_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3063_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_0_0_wb_clk_i),
    .D(_0163_),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3064_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_6_0_wb_clk_i),
    .D(_0164_),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3065_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_6_0_wb_clk_i),
    .D(_0165_),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3066_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_6_0_wb_clk_i),
    .D(_0166_),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3067_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_3_0_wb_clk_i),
    .D(_0167_),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3068_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0168_),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3069_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_3_0_wb_clk_i),
    .D(_0169_),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3070_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0170_),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3071_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_6_0_wb_clk_i),
    .D(_0171_),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3072_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0172_),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3073_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0173_),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3074_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0174_),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3075_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0175_),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3076_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0176_),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3077_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0177_),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3078_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0178_),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3079_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_3_0_wb_clk_i),
    .D(_0179_),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3080_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0180_),
    .Q(\tt_um_rejunity_sn76489.clk_counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3081_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0181_),
    .Q(\tt_um_rejunity_sn76489.clk_counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3082_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_11_0_wb_clk_i),
    .D(_0182_),
    .Q(\tt_um_rejunity_sn76489.clk_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3083_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0183_),
    .Q(\tt_um_rejunity_sn76489.clk_counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3084_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0184_),
    .Q(\tt_um_rejunity_sn76489.clk_counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3085_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0185_),
    .Q(\tt_um_rejunity_sn76489.clk_counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3086_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_14_0_wb_clk_i),
    .D(_0186_),
    .Q(\tt_um_rejunity_sn76489.clk_counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3087_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_3_0_wb_clk_i),
    .D(_0187_),
    .Q(\tt_um_rejunity_sn76489.latch_control_reg[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3088_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_3_0_wb_clk_i),
    .D(_0188_),
    .Q(\tt_um_rejunity_sn76489.latch_control_reg[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3089_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_3_0_wb_clk_i),
    .D(_0189_),
    .Q(\tt_um_rejunity_sn76489.latch_control_reg[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3090_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0190_),
    .Q(\tt_um_rejunity_sn76489.control_noise[0][0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3091_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_9_0_wb_clk_i),
    .D(_0191_),
    .Q(\tt_um_rejunity_sn76489.control_noise[0][1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _3092_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_4_1_0_wb_clk_i),
    .D(_0192_),
    .Q(\tt_um_rejunity_sn76489.control_noise[0][2] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _3105_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.genblk4[0].pwm.accumulator[10] ),
    .Y(net26));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _3106_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.genblk4[1].pwm.accumulator[10] ),
    .Y(net27));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _3107_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.genblk4[2].pwm.accumulator[10] ),
    .Y(net12));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _3108_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.genblk4[3].pwm.accumulator[10] ),
    .Y(net13));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _3109_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.pwm.accumulator[12] ),
    .Y(net14));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _3110_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.DAC_dat ),
    .Y(net15));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _3111_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.DAC_le ),
    .Y(net16));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _3112_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\tt_um_rejunity_sn76489.DAC_clk ),
    .Y(net17));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(wb_clk_i),
    .Y(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_0_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_0_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_10_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_11_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_11_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_12_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_13_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_14_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_15_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_1_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_1_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_2_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_3_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_4_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_5_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_6_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_7_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_7_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_8_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_4_9_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_4_9_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload0 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_1_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload1 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_2_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_11_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_12_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_13_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_14_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_15_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_3_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload3 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_4_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_5_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_6_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_7_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkload7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_8_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_6 clkload8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_9_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_4 clkload9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_4_10_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input1 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[0]),
    .Y(net1));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_2),
    .Y(net10));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(rst_n),
    .Y(net11));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(custom_settings[1]),
    .Y(net2));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input3 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[1]),
    .Y(net3));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[2]),
    .Y(net4));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[3]),
    .Y(net5));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[4]),
    .Y(net6));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[5]),
    .Y(net7));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[6]),
    .Y(net8));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in_1[7]),
    .Y(net9));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net12),
    .Y(io_out[10]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net13),
    .Y(io_out[11]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net14),
    .Y(io_out[12]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net15),
    .Y(io_out[17]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net16),
    .Y(io_out[18]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net17),
    .Y(io_out[19]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net18),
    .Y(io_out[20]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net19),
    .Y(io_out[21]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net20),
    .Y(io_out[22]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net21),
    .Y(io_out[23]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net22),
    .Y(io_out[24]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net23),
    .Y(io_out[25]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net24),
    .Y(io_out[26]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net25),
    .Y(io_out[27]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net26),
    .Y(io_out[8]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net27),
    .Y(io_out[9]));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net28));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net29));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net30));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net31));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net32));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net33));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net34));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_35 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net35));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net36));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net37));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net38));
 gf180mcu_as_sc_mcu7t3v3__tiel_4 wrapped_sn76489_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .ZERO(net39));
 assign io_out[0] = net28;
 assign io_out[13] = net36;
 assign io_out[14] = net37;
 assign io_out[15] = net38;
 assign io_out[16] = net39;
 assign io_out[1] = net29;
 assign io_out[2] = net30;
 assign io_out[3] = net31;
 assign io_out[4] = net32;
 assign io_out[5] = net33;
 assign io_out[6] = net34;
 assign io_out[7] = net35;
endmodule
