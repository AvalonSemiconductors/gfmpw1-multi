VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_sn76489
  CLASS BLOCK ;
  FOREIGN wrapped_sn76489 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 350.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 295.680 300.000 296.240 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 330.400 300.000 330.960 ;
    END
  END custom_settings[1]
  PIN io_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 17.920 300.000 18.480 ;
    END
  END io_in_1[0]
  PIN io_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 52.640 300.000 53.200 ;
    END
  END io_in_1[1]
  PIN io_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 87.360 300.000 87.920 ;
    END
  END io_in_1[2]
  PIN io_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 122.080 300.000 122.640 ;
    END
  END io_in_1[3]
  PIN io_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 156.800 300.000 157.360 ;
    END
  END io_in_1[4]
  PIN io_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 191.520 300.000 192.080 ;
    END
  END io_in_1[5]
  PIN io_in_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 226.240 300.000 226.800 ;
    END
  END io_in_1[6]
  PIN io_in_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 260.960 300.000 261.520 ;
    END
  END io_in_1[7]
  PIN io_in_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.200 4.000 291.760 ;
    END
  END io_in_2
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 346.000 14.000 350.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 346.000 114.800 350.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 346.000 124.880 350.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 346.000 134.960 350.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 346.000 145.040 350.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 346.000 155.120 350.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 346.000 165.200 350.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 346.000 175.280 350.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 346.000 185.360 350.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 346.000 195.440 350.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 346.000 205.520 350.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 346.000 24.080 350.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 346.000 215.600 350.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 346.000 225.680 350.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 346.000 235.760 350.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 346.000 245.840 350.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 346.000 255.920 350.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 346.000 266.000 350.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 346.000 276.080 350.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 346.000 286.160 350.000 ;
    END
  END io_out[27]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 346.000 34.160 350.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 346.000 44.240 350.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 346.000 54.320 350.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 346.000 64.400 350.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 346.000 74.480 350.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 346.000 84.560 350.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 346.000 94.640 350.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 346.000 104.720 350.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 333.500 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 333.500 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 58.240 4.000 58.800 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 334.170 ;
      LAYER Metal2 ;
        RECT 8.540 345.700 13.140 346.000 ;
        RECT 14.300 345.700 23.220 346.000 ;
        RECT 24.380 345.700 33.300 346.000 ;
        RECT 34.460 345.700 43.380 346.000 ;
        RECT 44.540 345.700 53.460 346.000 ;
        RECT 54.620 345.700 63.540 346.000 ;
        RECT 64.700 345.700 73.620 346.000 ;
        RECT 74.780 345.700 83.700 346.000 ;
        RECT 84.860 345.700 93.780 346.000 ;
        RECT 94.940 345.700 103.860 346.000 ;
        RECT 105.020 345.700 113.940 346.000 ;
        RECT 115.100 345.700 124.020 346.000 ;
        RECT 125.180 345.700 134.100 346.000 ;
        RECT 135.260 345.700 144.180 346.000 ;
        RECT 145.340 345.700 154.260 346.000 ;
        RECT 155.420 345.700 164.340 346.000 ;
        RECT 165.500 345.700 174.420 346.000 ;
        RECT 175.580 345.700 184.500 346.000 ;
        RECT 185.660 345.700 194.580 346.000 ;
        RECT 195.740 345.700 204.660 346.000 ;
        RECT 205.820 345.700 214.740 346.000 ;
        RECT 215.900 345.700 224.820 346.000 ;
        RECT 225.980 345.700 234.900 346.000 ;
        RECT 236.060 345.700 244.980 346.000 ;
        RECT 246.140 345.700 255.060 346.000 ;
        RECT 256.220 345.700 265.140 346.000 ;
        RECT 266.300 345.700 275.220 346.000 ;
        RECT 276.380 345.700 285.300 346.000 ;
        RECT 286.460 345.700 292.180 346.000 ;
        RECT 8.540 15.490 292.180 345.700 ;
      LAYER Metal3 ;
        RECT 4.000 331.260 296.000 334.180 ;
        RECT 4.000 330.100 295.700 331.260 ;
        RECT 4.000 296.540 296.000 330.100 ;
        RECT 4.000 295.380 295.700 296.540 ;
        RECT 4.000 292.060 296.000 295.380 ;
        RECT 4.300 290.900 296.000 292.060 ;
        RECT 4.000 261.820 296.000 290.900 ;
        RECT 4.000 260.660 295.700 261.820 ;
        RECT 4.000 227.100 296.000 260.660 ;
        RECT 4.000 225.940 295.700 227.100 ;
        RECT 4.000 192.380 296.000 225.940 ;
        RECT 4.000 191.220 295.700 192.380 ;
        RECT 4.000 175.580 296.000 191.220 ;
        RECT 4.300 174.420 296.000 175.580 ;
        RECT 4.000 157.660 296.000 174.420 ;
        RECT 4.000 156.500 295.700 157.660 ;
        RECT 4.000 122.940 296.000 156.500 ;
        RECT 4.000 121.780 295.700 122.940 ;
        RECT 4.000 88.220 296.000 121.780 ;
        RECT 4.000 87.060 295.700 88.220 ;
        RECT 4.000 59.100 296.000 87.060 ;
        RECT 4.300 57.940 296.000 59.100 ;
        RECT 4.000 53.500 296.000 57.940 ;
        RECT 4.000 52.340 295.700 53.500 ;
        RECT 4.000 18.780 296.000 52.340 ;
        RECT 4.000 17.620 295.700 18.780 ;
        RECT 4.000 15.540 296.000 17.620 ;
      LAYER Metal4 ;
        RECT 21.420 37.050 21.940 315.750 ;
        RECT 24.140 37.050 98.740 315.750 ;
        RECT 100.940 37.050 175.540 315.750 ;
        RECT 177.740 37.050 252.340 315.750 ;
        RECT 254.540 37.050 287.700 315.750 ;
  END
END wrapped_sn76489
END LIBRARY

