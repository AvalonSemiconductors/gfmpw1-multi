VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_sid
  CLASS BLOCK ;
  FOREIGN wrapped_sid ;
  ORIGIN 0.000 0.000 ;
  SIZE 1150.000 BY 800.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 13.440 1150.000 14.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 159.040 1150.000 159.600 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 173.600 1150.000 174.160 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 188.160 1150.000 188.720 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 202.720 1150.000 203.280 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 217.280 1150.000 217.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 231.840 1150.000 232.400 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 246.400 1150.000 246.960 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 260.960 1150.000 261.520 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 275.520 1150.000 276.080 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 290.080 1150.000 290.640 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 28.000 1150.000 28.560 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 304.640 1150.000 305.200 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 319.200 1150.000 319.760 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 333.760 1150.000 334.320 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 348.320 1150.000 348.880 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 362.880 1150.000 363.440 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 377.440 1150.000 378.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 392.000 1150.000 392.560 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 406.560 1150.000 407.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 421.120 1150.000 421.680 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 435.680 1150.000 436.240 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 42.560 1150.000 43.120 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 450.240 1150.000 450.800 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 464.800 1150.000 465.360 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 479.360 1150.000 479.920 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 57.120 1150.000 57.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 71.680 1150.000 72.240 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 86.240 1150.000 86.800 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 100.800 1150.000 101.360 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 115.360 1150.000 115.920 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 129.920 1150.000 130.480 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 144.480 1150.000 145.040 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 796.000 575.120 800.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 493.920 1150.000 494.480 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 639.520 1150.000 640.080 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 654.080 1150.000 654.640 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 668.640 1150.000 669.200 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 683.200 1150.000 683.760 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 697.760 1150.000 698.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 712.320 1150.000 712.880 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 726.880 1150.000 727.440 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 741.440 1150.000 742.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 756.000 1150.000 756.560 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 770.560 1150.000 771.120 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 508.480 1150.000 509.040 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 785.120 1150.000 785.680 ;
    END
  END io_out[20]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 523.040 1150.000 523.600 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 537.600 1150.000 538.160 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 552.160 1150.000 552.720 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 566.720 1150.000 567.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 581.280 1150.000 581.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 595.840 1150.000 596.400 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 610.400 1150.000 610.960 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 624.960 1150.000 625.520 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 0.000 861.840 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 784.300 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 0.000 287.280 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Pwell ;
        RECT 6.290 782.240 1143.390 784.430 ;
      LAYER Nwell ;
        RECT 6.290 778.045 1143.390 782.240 ;
        RECT 6.290 777.920 189.990 778.045 ;
      LAYER Pwell ;
        RECT 6.290 774.400 1143.390 777.920 ;
      LAYER Nwell ;
        RECT 6.290 774.275 180.785 774.400 ;
        RECT 6.290 770.205 1143.390 774.275 ;
        RECT 6.290 770.080 111.870 770.205 ;
      LAYER Pwell ;
        RECT 6.290 766.560 1143.390 770.080 ;
      LAYER Nwell ;
        RECT 6.290 766.435 134.925 766.560 ;
        RECT 6.290 762.365 1143.390 766.435 ;
        RECT 6.290 762.240 116.350 762.365 ;
      LAYER Pwell ;
        RECT 6.290 758.720 1143.390 762.240 ;
      LAYER Nwell ;
        RECT 6.290 758.595 104.895 758.720 ;
        RECT 6.290 754.525 1143.390 758.595 ;
        RECT 6.290 754.400 74.930 754.525 ;
      LAYER Pwell ;
        RECT 6.290 750.880 1143.390 754.400 ;
      LAYER Nwell ;
        RECT 6.290 750.755 112.425 750.880 ;
        RECT 6.290 746.685 1143.390 750.755 ;
        RECT 6.290 746.560 109.105 746.685 ;
      LAYER Pwell ;
        RECT 6.290 743.040 1143.390 746.560 ;
      LAYER Nwell ;
        RECT 6.290 742.915 82.470 743.040 ;
        RECT 6.290 738.845 1143.390 742.915 ;
        RECT 6.290 738.720 82.190 738.845 ;
      LAYER Pwell ;
        RECT 6.290 735.200 1143.390 738.720 ;
      LAYER Nwell ;
        RECT 6.290 735.075 65.180 735.200 ;
        RECT 6.290 731.005 1143.390 735.075 ;
        RECT 6.290 730.880 76.635 731.005 ;
      LAYER Pwell ;
        RECT 6.290 727.360 1143.390 730.880 ;
      LAYER Nwell ;
        RECT 6.290 727.235 51.950 727.360 ;
        RECT 6.290 723.165 1143.390 727.235 ;
        RECT 6.290 723.040 79.435 723.165 ;
      LAYER Pwell ;
        RECT 6.290 719.520 1143.390 723.040 ;
      LAYER Nwell ;
        RECT 6.290 719.395 39.115 719.520 ;
        RECT 6.290 715.325 1143.390 719.395 ;
        RECT 6.290 715.200 38.510 715.325 ;
      LAYER Pwell ;
        RECT 6.290 711.680 1143.390 715.200 ;
      LAYER Nwell ;
        RECT 6.290 711.555 48.590 711.680 ;
        RECT 6.290 707.485 1143.390 711.555 ;
        RECT 6.290 707.360 12.680 707.485 ;
      LAYER Pwell ;
        RECT 6.290 703.840 1143.390 707.360 ;
      LAYER Nwell ;
        RECT 6.290 703.715 29.550 703.840 ;
        RECT 6.290 699.645 1143.390 703.715 ;
        RECT 6.290 699.520 11.070 699.645 ;
      LAYER Pwell ;
        RECT 6.290 696.000 1143.390 699.520 ;
      LAYER Nwell ;
        RECT 6.290 695.875 87.790 696.000 ;
        RECT 6.290 691.805 1143.390 695.875 ;
        RECT 6.290 691.680 31.790 691.805 ;
      LAYER Pwell ;
        RECT 6.290 688.160 1143.390 691.680 ;
      LAYER Nwell ;
        RECT 6.290 688.035 20.310 688.160 ;
        RECT 6.290 683.965 1143.390 688.035 ;
        RECT 6.290 683.840 108.510 683.965 ;
      LAYER Pwell ;
        RECT 6.290 680.320 1143.390 683.840 ;
      LAYER Nwell ;
        RECT 6.290 680.195 16.155 680.320 ;
        RECT 6.290 676.125 1143.390 680.195 ;
        RECT 6.290 676.000 14.430 676.125 ;
      LAYER Pwell ;
        RECT 6.290 672.480 1143.390 676.000 ;
      LAYER Nwell ;
        RECT 6.290 672.355 13.310 672.480 ;
        RECT 6.290 668.285 1143.390 672.355 ;
        RECT 6.290 668.160 79.390 668.285 ;
      LAYER Pwell ;
        RECT 6.290 664.640 1143.390 668.160 ;
      LAYER Nwell ;
        RECT 6.290 664.515 10.510 664.640 ;
        RECT 6.290 660.445 1143.390 664.515 ;
        RECT 6.290 660.320 18.945 660.445 ;
      LAYER Pwell ;
        RECT 6.290 656.800 1143.390 660.320 ;
      LAYER Nwell ;
        RECT 6.290 656.675 69.345 656.800 ;
        RECT 6.290 652.605 1143.390 656.675 ;
        RECT 6.290 652.480 137.115 652.605 ;
      LAYER Pwell ;
        RECT 6.290 648.960 1143.390 652.480 ;
      LAYER Nwell ;
        RECT 6.290 648.835 15.595 648.960 ;
        RECT 6.290 644.765 1143.390 648.835 ;
        RECT 6.290 644.640 42.150 644.765 ;
      LAYER Pwell ;
        RECT 6.290 641.120 1143.390 644.640 ;
      LAYER Nwell ;
        RECT 6.290 640.995 16.110 641.120 ;
        RECT 6.290 636.925 1143.390 640.995 ;
        RECT 6.290 636.800 72.670 636.925 ;
      LAYER Pwell ;
        RECT 6.290 633.280 1143.390 636.800 ;
      LAYER Nwell ;
        RECT 6.290 633.155 101.790 633.280 ;
        RECT 6.290 629.085 1143.390 633.155 ;
        RECT 6.290 628.960 10.510 629.085 ;
      LAYER Pwell ;
        RECT 6.290 625.440 1143.390 628.960 ;
      LAYER Nwell ;
        RECT 6.290 625.315 34.625 625.440 ;
        RECT 6.290 621.245 1143.390 625.315 ;
        RECT 6.290 621.120 42.150 621.245 ;
      LAYER Pwell ;
        RECT 6.290 617.600 1143.390 621.120 ;
      LAYER Nwell ;
        RECT 6.290 617.475 12.745 617.600 ;
        RECT 6.290 613.405 1143.390 617.475 ;
        RECT 6.290 613.280 84.430 613.405 ;
      LAYER Pwell ;
        RECT 6.290 609.760 1143.390 613.280 ;
      LAYER Nwell ;
        RECT 6.290 609.635 284.955 609.760 ;
        RECT 6.290 605.565 1143.390 609.635 ;
        RECT 6.290 605.440 71.550 605.565 ;
      LAYER Pwell ;
        RECT 6.290 601.920 1143.390 605.440 ;
      LAYER Nwell ;
        RECT 6.290 601.795 50.875 601.920 ;
        RECT 6.290 597.725 1143.390 601.795 ;
        RECT 6.290 597.600 31.275 597.725 ;
      LAYER Pwell ;
        RECT 6.290 594.080 1143.390 597.600 ;
      LAYER Nwell ;
        RECT 6.290 593.955 14.580 594.080 ;
        RECT 6.290 589.885 1143.390 593.955 ;
        RECT 6.290 589.760 82.190 589.885 ;
      LAYER Pwell ;
        RECT 6.290 586.240 1143.390 589.760 ;
      LAYER Nwell ;
        RECT 6.290 586.115 150.230 586.240 ;
        RECT 6.290 582.045 1143.390 586.115 ;
        RECT 6.290 581.920 16.390 582.045 ;
      LAYER Pwell ;
        RECT 6.290 578.400 1143.390 581.920 ;
      LAYER Nwell ;
        RECT 6.290 578.275 82.470 578.400 ;
        RECT 6.290 574.205 1143.390 578.275 ;
        RECT 6.290 574.080 49.710 574.205 ;
      LAYER Pwell ;
        RECT 6.290 570.560 1143.390 574.080 ;
      LAYER Nwell ;
        RECT 6.290 570.435 53.350 570.560 ;
        RECT 6.290 566.365 1143.390 570.435 ;
        RECT 6.290 566.240 36.425 566.365 ;
      LAYER Pwell ;
        RECT 6.290 562.720 1143.390 566.240 ;
      LAYER Nwell ;
        RECT 6.290 562.595 15.900 562.720 ;
        RECT 6.290 558.525 1143.390 562.595 ;
        RECT 6.290 558.400 72.950 558.525 ;
      LAYER Pwell ;
        RECT 6.290 554.880 1143.390 558.400 ;
      LAYER Nwell ;
        RECT 6.290 554.755 34.625 554.880 ;
        RECT 6.290 550.685 1143.390 554.755 ;
        RECT 6.290 550.560 119.820 550.685 ;
      LAYER Pwell ;
        RECT 6.290 547.040 1143.390 550.560 ;
      LAYER Nwell ;
        RECT 6.290 546.915 97.265 547.040 ;
        RECT 6.290 542.845 1143.390 546.915 ;
        RECT 6.290 542.720 20.940 542.845 ;
      LAYER Pwell ;
        RECT 6.290 539.200 1143.390 542.720 ;
      LAYER Nwell ;
        RECT 6.290 539.075 106.785 539.200 ;
        RECT 6.290 535.005 1143.390 539.075 ;
        RECT 6.290 534.880 39.025 535.005 ;
      LAYER Pwell ;
        RECT 6.290 531.360 1143.390 534.880 ;
      LAYER Nwell ;
        RECT 6.290 531.235 12.705 531.360 ;
        RECT 6.290 527.165 1143.390 531.235 ;
        RECT 6.290 527.040 155.505 527.165 ;
      LAYER Pwell ;
        RECT 6.290 523.520 1143.390 527.040 ;
      LAYER Nwell ;
        RECT 6.290 523.395 28.780 523.520 ;
        RECT 6.290 519.325 1143.390 523.395 ;
        RECT 6.290 519.200 12.705 519.325 ;
      LAYER Pwell ;
        RECT 6.290 515.680 1143.390 519.200 ;
      LAYER Nwell ;
        RECT 6.290 515.555 19.470 515.680 ;
        RECT 6.290 511.485 1143.390 515.555 ;
        RECT 6.290 511.360 68.190 511.485 ;
      LAYER Pwell ;
        RECT 6.290 507.840 1143.390 511.360 ;
      LAYER Nwell ;
        RECT 6.290 507.715 17.960 507.840 ;
        RECT 6.290 503.645 1143.390 507.715 ;
        RECT 6.290 503.520 90.740 503.645 ;
      LAYER Pwell ;
        RECT 6.290 500.000 1143.390 503.520 ;
      LAYER Nwell ;
        RECT 6.290 499.875 24.100 500.000 ;
        RECT 6.290 495.805 1143.390 499.875 ;
        RECT 6.290 495.680 47.960 495.805 ;
      LAYER Pwell ;
        RECT 6.290 492.160 1143.390 495.680 ;
      LAYER Nwell ;
        RECT 6.290 492.035 30.950 492.160 ;
        RECT 6.290 487.965 1143.390 492.035 ;
        RECT 6.290 487.840 93.000 487.965 ;
      LAYER Pwell ;
        RECT 6.290 484.320 1143.390 487.840 ;
      LAYER Nwell ;
        RECT 6.290 484.195 118.200 484.320 ;
        RECT 6.290 480.125 1143.390 484.195 ;
        RECT 6.290 480.000 52.300 480.125 ;
      LAYER Pwell ;
        RECT 6.290 476.480 1143.390 480.000 ;
      LAYER Nwell ;
        RECT 6.290 476.355 34.065 476.480 ;
        RECT 6.290 472.285 1143.390 476.355 ;
        RECT 6.290 472.160 34.380 472.285 ;
      LAYER Pwell ;
        RECT 6.290 468.640 1143.390 472.160 ;
      LAYER Nwell ;
        RECT 6.290 468.515 52.655 468.640 ;
        RECT 6.290 464.445 1143.390 468.515 ;
        RECT 6.290 464.320 40.540 464.445 ;
      LAYER Pwell ;
        RECT 6.290 460.800 1143.390 464.320 ;
      LAYER Nwell ;
        RECT 6.290 460.675 112.220 460.800 ;
        RECT 6.290 456.605 1143.390 460.675 ;
        RECT 6.290 456.480 15.340 456.605 ;
      LAYER Pwell ;
        RECT 6.290 452.960 1143.390 456.480 ;
      LAYER Nwell ;
        RECT 6.290 452.835 27.905 452.960 ;
        RECT 6.290 448.765 1143.390 452.835 ;
        RECT 6.290 448.640 15.270 448.765 ;
      LAYER Pwell ;
        RECT 6.290 445.120 1143.390 448.640 ;
      LAYER Nwell ;
        RECT 6.290 444.995 15.900 445.120 ;
        RECT 6.290 440.925 1143.390 444.995 ;
        RECT 6.290 440.800 18.945 440.925 ;
      LAYER Pwell ;
        RECT 6.290 437.280 1143.390 440.800 ;
      LAYER Nwell ;
        RECT 6.290 437.155 17.960 437.280 ;
        RECT 6.290 433.085 1143.390 437.155 ;
        RECT 6.290 432.960 95.155 433.085 ;
      LAYER Pwell ;
        RECT 6.290 429.440 1143.390 432.960 ;
      LAYER Nwell ;
        RECT 6.290 429.315 51.905 429.440 ;
        RECT 6.290 425.245 1143.390 429.315 ;
        RECT 6.290 425.120 33.985 425.245 ;
      LAYER Pwell ;
        RECT 6.290 421.600 1143.390 425.120 ;
      LAYER Nwell ;
        RECT 6.290 421.475 118.200 421.600 ;
        RECT 6.290 417.405 1143.390 421.475 ;
        RECT 6.290 417.280 228.305 417.405 ;
      LAYER Pwell ;
        RECT 6.290 413.760 1143.390 417.280 ;
      LAYER Nwell ;
        RECT 6.290 413.635 20.545 413.760 ;
        RECT 6.290 409.565 1143.390 413.635 ;
        RECT 6.290 409.440 89.640 409.565 ;
      LAYER Pwell ;
        RECT 6.290 405.920 1143.390 409.440 ;
      LAYER Nwell ;
        RECT 6.290 405.795 522.305 405.920 ;
        RECT 6.290 401.725 1143.390 405.795 ;
        RECT 6.290 401.600 210.945 401.725 ;
      LAYER Pwell ;
        RECT 6.290 398.080 1143.390 401.600 ;
      LAYER Nwell ;
        RECT 6.290 397.955 19.425 398.080 ;
        RECT 6.290 393.885 1143.390 397.955 ;
        RECT 6.290 393.760 162.915 393.885 ;
      LAYER Pwell ;
        RECT 6.290 390.240 1143.390 393.760 ;
      LAYER Nwell ;
        RECT 6.290 390.115 170.105 390.240 ;
        RECT 6.290 386.045 1143.390 390.115 ;
        RECT 6.290 385.920 48.200 386.045 ;
      LAYER Pwell ;
        RECT 6.290 382.400 1143.390 385.920 ;
      LAYER Nwell ;
        RECT 6.290 382.275 43.270 382.400 ;
        RECT 6.290 378.205 1143.390 382.275 ;
        RECT 6.290 378.080 45.835 378.205 ;
      LAYER Pwell ;
        RECT 6.290 374.560 1143.390 378.080 ;
      LAYER Nwell ;
        RECT 6.290 374.435 100.390 374.560 ;
        RECT 6.290 370.365 1143.390 374.435 ;
        RECT 6.290 370.240 51.390 370.365 ;
      LAYER Pwell ;
        RECT 6.290 366.720 1143.390 370.240 ;
      LAYER Nwell ;
        RECT 6.290 366.595 33.505 366.720 ;
        RECT 6.290 362.525 1143.390 366.595 ;
        RECT 6.290 362.400 129.230 362.525 ;
      LAYER Pwell ;
        RECT 6.290 358.880 1143.390 362.400 ;
      LAYER Nwell ;
        RECT 6.290 358.755 28.150 358.880 ;
        RECT 6.290 354.685 1143.390 358.755 ;
        RECT 6.290 354.560 115.275 354.685 ;
      LAYER Pwell ;
        RECT 6.290 351.040 1143.390 354.560 ;
      LAYER Nwell ;
        RECT 6.290 350.915 91.710 351.040 ;
        RECT 6.290 346.845 1143.390 350.915 ;
        RECT 6.290 346.720 56.990 346.845 ;
      LAYER Pwell ;
        RECT 6.290 343.200 1143.390 346.720 ;
      LAYER Nwell ;
        RECT 6.290 343.075 110.470 343.200 ;
        RECT 6.290 339.005 1143.390 343.075 ;
        RECT 6.290 338.880 40.470 339.005 ;
      LAYER Pwell ;
        RECT 6.290 335.360 1143.390 338.880 ;
      LAYER Nwell ;
        RECT 6.290 335.235 48.590 335.360 ;
        RECT 6.290 331.165 1143.390 335.235 ;
        RECT 6.290 331.040 194.360 331.165 ;
      LAYER Pwell ;
        RECT 6.290 327.520 1143.390 331.040 ;
      LAYER Nwell ;
        RECT 6.290 327.395 254.840 327.520 ;
        RECT 6.290 323.325 1143.390 327.395 ;
        RECT 6.290 323.200 18.395 323.325 ;
      LAYER Pwell ;
        RECT 6.290 319.680 1143.390 323.200 ;
      LAYER Nwell ;
        RECT 6.290 319.555 36.305 319.680 ;
        RECT 6.290 315.485 1143.390 319.555 ;
        RECT 6.290 315.360 78.270 315.485 ;
      LAYER Pwell ;
        RECT 6.290 311.840 1143.390 315.360 ;
      LAYER Nwell ;
        RECT 6.290 311.715 77.710 311.840 ;
        RECT 6.290 307.645 1143.390 311.715 ;
        RECT 6.290 307.520 14.710 307.645 ;
      LAYER Pwell ;
        RECT 6.290 304.000 1143.390 307.520 ;
      LAYER Nwell ;
        RECT 6.290 303.875 96.470 304.000 ;
        RECT 6.290 299.805 1143.390 303.875 ;
        RECT 6.290 299.680 131.750 299.805 ;
      LAYER Pwell ;
        RECT 6.290 296.160 1143.390 299.680 ;
      LAYER Nwell ;
        RECT 6.290 296.035 40.470 296.160 ;
        RECT 6.290 291.965 1143.390 296.035 ;
        RECT 6.290 291.840 127.270 291.965 ;
      LAYER Pwell ;
        RECT 6.290 288.320 1143.390 291.840 ;
      LAYER Nwell ;
        RECT 6.290 288.195 12.750 288.320 ;
        RECT 6.290 284.125 1143.390 288.195 ;
        RECT 6.290 284.000 38.510 284.125 ;
      LAYER Pwell ;
        RECT 6.290 280.480 1143.390 284.000 ;
      LAYER Nwell ;
        RECT 6.290 280.355 171.840 280.480 ;
        RECT 6.290 276.285 1143.390 280.355 ;
        RECT 6.290 276.160 41.355 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 1143.390 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 13.310 272.640 ;
        RECT 6.290 268.445 1143.390 272.515 ;
        RECT 6.290 268.320 127.830 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 1143.390 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 41.030 264.800 ;
        RECT 6.290 260.605 1143.390 264.675 ;
        RECT 6.290 260.480 19.750 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 1143.390 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 16.950 256.960 ;
        RECT 6.290 252.765 1143.390 256.835 ;
        RECT 6.290 252.640 111.310 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 1143.390 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 13.825 249.120 ;
        RECT 6.290 244.925 1143.390 248.995 ;
        RECT 6.290 244.800 35.710 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 1143.390 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 14.385 241.280 ;
        RECT 6.290 237.085 1143.390 241.155 ;
        RECT 6.290 236.960 110.705 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 1143.390 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 12.705 233.440 ;
        RECT 6.290 229.245 1143.390 233.315 ;
        RECT 6.290 229.120 45.745 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 1143.390 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 51.905 225.600 ;
        RECT 6.290 221.405 1143.390 225.475 ;
        RECT 6.290 221.280 13.265 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 1143.390 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 48.180 217.760 ;
        RECT 6.290 213.565 1143.390 217.635 ;
        RECT 6.290 213.440 58.280 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 1143.390 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 14.945 209.920 ;
        RECT 6.290 205.725 1143.390 209.795 ;
        RECT 6.290 205.600 79.905 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 1143.390 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 12.705 202.080 ;
        RECT 6.290 197.885 1143.390 201.955 ;
        RECT 6.290 197.760 51.560 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 1143.390 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 13.265 194.240 ;
        RECT 6.290 190.045 1143.390 194.115 ;
        RECT 6.290 189.920 39.125 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 1143.390 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 336.945 186.400 ;
        RECT 6.290 182.205 1143.390 186.275 ;
        RECT 6.290 182.080 13.825 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 1143.390 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 12.705 178.560 ;
        RECT 6.290 174.365 1143.390 178.435 ;
        RECT 6.290 174.240 39.125 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 1143.390 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 57.160 170.720 ;
        RECT 6.290 166.525 1143.390 170.595 ;
        RECT 6.290 166.400 17.960 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 1143.390 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 249.025 162.880 ;
        RECT 6.290 158.685 1143.390 162.755 ;
        RECT 6.290 158.560 71.505 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 1143.390 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 12.705 155.040 ;
        RECT 6.290 150.845 1143.390 154.915 ;
        RECT 6.290 150.720 199.960 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 1143.390 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 12.705 147.200 ;
        RECT 6.290 143.005 1143.390 147.075 ;
        RECT 6.290 142.880 42.485 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 1143.390 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 109.025 139.360 ;
        RECT 6.290 135.165 1143.390 139.235 ;
        RECT 6.290 135.040 12.705 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 1143.390 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 25.585 131.520 ;
        RECT 6.290 127.325 1143.390 131.395 ;
        RECT 6.290 127.200 14.945 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 1143.390 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 52.465 123.680 ;
        RECT 6.290 119.485 1143.390 123.555 ;
        RECT 6.290 119.360 12.705 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 1143.390 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 32.305 115.840 ;
        RECT 6.290 111.645 1143.390 115.715 ;
        RECT 6.290 111.520 34.545 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 1143.390 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 103.985 108.000 ;
        RECT 6.290 103.805 1143.390 107.875 ;
        RECT 6.290 103.680 87.960 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 1143.390 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 103.425 100.160 ;
        RECT 6.290 95.965 1143.390 100.035 ;
        RECT 6.290 95.840 160.545 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 1143.390 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 130.305 92.320 ;
        RECT 6.290 88.125 1143.390 92.195 ;
        RECT 6.290 88.000 118.545 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 1143.390 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 140.385 84.480 ;
        RECT 6.290 80.285 1143.390 84.355 ;
        RECT 6.290 80.160 124.145 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 1143.390 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 105.105 76.640 ;
        RECT 6.290 72.445 1143.390 76.515 ;
        RECT 6.290 72.320 151.765 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 1143.390 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 112.945 68.800 ;
        RECT 6.290 64.605 1143.390 68.675 ;
        RECT 6.290 64.480 156.805 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 1143.390 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 106.785 60.960 ;
        RECT 6.290 56.765 1143.390 60.835 ;
        RECT 6.290 56.640 362.680 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 1143.390 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 139.825 53.120 ;
        RECT 6.290 48.925 1143.390 52.995 ;
        RECT 6.290 48.800 123.025 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 1143.390 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 146.200 45.280 ;
        RECT 6.290 41.085 1143.390 45.155 ;
        RECT 6.290 40.960 250.145 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 1143.390 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 209.265 37.440 ;
        RECT 6.290 33.245 1143.390 37.315 ;
        RECT 6.290 33.120 149.905 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 1143.390 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 171.745 29.600 ;
        RECT 6.290 25.405 1143.390 29.475 ;
        RECT 6.290 25.280 250.920 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 1143.390 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 188.545 21.760 ;
        RECT 6.290 17.565 1143.390 21.635 ;
        RECT 6.290 17.440 514.680 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 1143.390 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 1142.960 784.300 ;
      LAYER Metal2 ;
        RECT 7.980 795.700 574.260 796.000 ;
        RECT 575.420 795.700 1141.700 796.000 ;
        RECT 7.980 4.300 1141.700 795.700 ;
        RECT 7.980 3.450 286.420 4.300 ;
        RECT 287.580 3.450 860.980 4.300 ;
        RECT 862.140 3.450 1141.700 4.300 ;
      LAYER Metal3 ;
        RECT 7.930 785.980 1146.000 792.820 ;
        RECT 7.930 784.820 1145.700 785.980 ;
        RECT 7.930 771.420 1146.000 784.820 ;
        RECT 7.930 770.260 1145.700 771.420 ;
        RECT 7.930 756.860 1146.000 770.260 ;
        RECT 7.930 755.700 1145.700 756.860 ;
        RECT 7.930 742.300 1146.000 755.700 ;
        RECT 7.930 741.140 1145.700 742.300 ;
        RECT 7.930 727.740 1146.000 741.140 ;
        RECT 7.930 726.580 1145.700 727.740 ;
        RECT 7.930 713.180 1146.000 726.580 ;
        RECT 7.930 712.020 1145.700 713.180 ;
        RECT 7.930 698.620 1146.000 712.020 ;
        RECT 7.930 697.460 1145.700 698.620 ;
        RECT 7.930 684.060 1146.000 697.460 ;
        RECT 7.930 682.900 1145.700 684.060 ;
        RECT 7.930 669.500 1146.000 682.900 ;
        RECT 7.930 668.340 1145.700 669.500 ;
        RECT 7.930 654.940 1146.000 668.340 ;
        RECT 7.930 653.780 1145.700 654.940 ;
        RECT 7.930 640.380 1146.000 653.780 ;
        RECT 7.930 639.220 1145.700 640.380 ;
        RECT 7.930 625.820 1146.000 639.220 ;
        RECT 7.930 624.660 1145.700 625.820 ;
        RECT 7.930 611.260 1146.000 624.660 ;
        RECT 7.930 610.100 1145.700 611.260 ;
        RECT 7.930 596.700 1146.000 610.100 ;
        RECT 7.930 595.540 1145.700 596.700 ;
        RECT 7.930 582.140 1146.000 595.540 ;
        RECT 7.930 580.980 1145.700 582.140 ;
        RECT 7.930 567.580 1146.000 580.980 ;
        RECT 7.930 566.420 1145.700 567.580 ;
        RECT 7.930 553.020 1146.000 566.420 ;
        RECT 7.930 551.860 1145.700 553.020 ;
        RECT 7.930 538.460 1146.000 551.860 ;
        RECT 7.930 537.300 1145.700 538.460 ;
        RECT 7.930 523.900 1146.000 537.300 ;
        RECT 7.930 522.740 1145.700 523.900 ;
        RECT 7.930 509.340 1146.000 522.740 ;
        RECT 7.930 508.180 1145.700 509.340 ;
        RECT 7.930 494.780 1146.000 508.180 ;
        RECT 7.930 493.620 1145.700 494.780 ;
        RECT 7.930 480.220 1146.000 493.620 ;
        RECT 7.930 479.060 1145.700 480.220 ;
        RECT 7.930 465.660 1146.000 479.060 ;
        RECT 7.930 464.500 1145.700 465.660 ;
        RECT 7.930 451.100 1146.000 464.500 ;
        RECT 7.930 449.940 1145.700 451.100 ;
        RECT 7.930 436.540 1146.000 449.940 ;
        RECT 7.930 435.380 1145.700 436.540 ;
        RECT 7.930 421.980 1146.000 435.380 ;
        RECT 7.930 420.820 1145.700 421.980 ;
        RECT 7.930 407.420 1146.000 420.820 ;
        RECT 7.930 406.260 1145.700 407.420 ;
        RECT 7.930 392.860 1146.000 406.260 ;
        RECT 7.930 391.700 1145.700 392.860 ;
        RECT 7.930 378.300 1146.000 391.700 ;
        RECT 7.930 377.140 1145.700 378.300 ;
        RECT 7.930 363.740 1146.000 377.140 ;
        RECT 7.930 362.580 1145.700 363.740 ;
        RECT 7.930 349.180 1146.000 362.580 ;
        RECT 7.930 348.020 1145.700 349.180 ;
        RECT 7.930 334.620 1146.000 348.020 ;
        RECT 7.930 333.460 1145.700 334.620 ;
        RECT 7.930 320.060 1146.000 333.460 ;
        RECT 7.930 318.900 1145.700 320.060 ;
        RECT 7.930 305.500 1146.000 318.900 ;
        RECT 7.930 304.340 1145.700 305.500 ;
        RECT 7.930 290.940 1146.000 304.340 ;
        RECT 7.930 289.780 1145.700 290.940 ;
        RECT 7.930 276.380 1146.000 289.780 ;
        RECT 7.930 275.220 1145.700 276.380 ;
        RECT 7.930 261.820 1146.000 275.220 ;
        RECT 7.930 260.660 1145.700 261.820 ;
        RECT 7.930 247.260 1146.000 260.660 ;
        RECT 7.930 246.100 1145.700 247.260 ;
        RECT 7.930 232.700 1146.000 246.100 ;
        RECT 7.930 231.540 1145.700 232.700 ;
        RECT 7.930 218.140 1146.000 231.540 ;
        RECT 7.930 216.980 1145.700 218.140 ;
        RECT 7.930 203.580 1146.000 216.980 ;
        RECT 7.930 202.420 1145.700 203.580 ;
        RECT 7.930 189.020 1146.000 202.420 ;
        RECT 7.930 187.860 1145.700 189.020 ;
        RECT 7.930 174.460 1146.000 187.860 ;
        RECT 7.930 173.300 1145.700 174.460 ;
        RECT 7.930 159.900 1146.000 173.300 ;
        RECT 7.930 158.740 1145.700 159.900 ;
        RECT 7.930 145.340 1146.000 158.740 ;
        RECT 7.930 144.180 1145.700 145.340 ;
        RECT 7.930 130.780 1146.000 144.180 ;
        RECT 7.930 129.620 1145.700 130.780 ;
        RECT 7.930 116.220 1146.000 129.620 ;
        RECT 7.930 115.060 1145.700 116.220 ;
        RECT 7.930 101.660 1146.000 115.060 ;
        RECT 7.930 100.500 1145.700 101.660 ;
        RECT 7.930 87.100 1146.000 100.500 ;
        RECT 7.930 85.940 1145.700 87.100 ;
        RECT 7.930 72.540 1146.000 85.940 ;
        RECT 7.930 71.380 1145.700 72.540 ;
        RECT 7.930 57.980 1146.000 71.380 ;
        RECT 7.930 56.820 1145.700 57.980 ;
        RECT 7.930 43.420 1146.000 56.820 ;
        RECT 7.930 42.260 1145.700 43.420 ;
        RECT 7.930 28.860 1146.000 42.260 ;
        RECT 7.930 27.700 1145.700 28.860 ;
        RECT 7.930 14.300 1146.000 27.700 ;
        RECT 7.930 13.140 1145.700 14.300 ;
        RECT 7.930 3.500 1146.000 13.140 ;
      LAYER Metal4 ;
        RECT 63.420 784.600 1133.300 791.750 ;
        RECT 63.420 15.080 98.740 784.600 ;
        RECT 100.940 15.080 175.540 784.600 ;
        RECT 177.740 15.080 252.340 784.600 ;
        RECT 254.540 15.080 329.140 784.600 ;
        RECT 331.340 15.080 405.940 784.600 ;
        RECT 408.140 15.080 482.740 784.600 ;
        RECT 484.940 15.080 559.540 784.600 ;
        RECT 561.740 15.080 636.340 784.600 ;
        RECT 638.540 15.080 713.140 784.600 ;
        RECT 715.340 15.080 789.940 784.600 ;
        RECT 792.140 15.080 866.740 784.600 ;
        RECT 868.940 15.080 943.540 784.600 ;
        RECT 945.740 15.080 1020.340 784.600 ;
        RECT 1022.540 15.080 1097.140 784.600 ;
        RECT 1099.340 15.080 1133.300 784.600 ;
        RECT 63.420 4.570 1133.300 15.080 ;
  END
END wrapped_sid
END LIBRARY

