magic
tech gf180mcuD
magscale 1 10
timestamp 1702458816
<< metal1 >>
rect 1344 42362 44576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 44576 42362
rect 1344 42276 44576 42310
rect 18286 42194 18338 42206
rect 18286 42130 18338 42142
rect 33518 42194 33570 42206
rect 33518 42130 33570 42142
rect 6190 42082 6242 42094
rect 9986 42030 9998 42082
rect 10050 42030 10062 42082
rect 6190 42018 6242 42030
rect 5070 41970 5122 41982
rect 5070 41906 5122 41918
rect 5854 41970 5906 41982
rect 5854 41906 5906 41918
rect 8878 41970 8930 41982
rect 8878 41906 8930 41918
rect 9662 41970 9714 41982
rect 13458 41918 13470 41970
rect 13522 41918 13534 41970
rect 17266 41918 17278 41970
rect 17330 41918 17342 41970
rect 21074 41918 21086 41970
rect 21138 41918 21150 41970
rect 24882 41918 24894 41970
rect 24946 41918 24958 41970
rect 28690 41918 28702 41970
rect 28754 41918 28766 41970
rect 32498 41918 32510 41970
rect 32562 41918 32574 41970
rect 36306 41918 36318 41970
rect 36370 41918 36382 41970
rect 40114 41918 40126 41970
rect 40178 41918 40190 41970
rect 9662 41906 9714 41918
rect 14478 41858 14530 41870
rect 14478 41794 14530 41806
rect 22094 41858 22146 41870
rect 22094 41794 22146 41806
rect 25902 41858 25954 41870
rect 25902 41794 25954 41806
rect 29710 41858 29762 41870
rect 29710 41794 29762 41806
rect 37326 41858 37378 41870
rect 37326 41794 37378 41806
rect 41134 41858 41186 41870
rect 41134 41794 41186 41806
rect 1344 41578 44576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 44576 41578
rect 1344 41492 44576 41526
rect 43586 41246 43598 41298
rect 43650 41246 43662 41298
rect 41570 41134 41582 41186
rect 41634 41134 41646 41186
rect 13918 40962 13970 40974
rect 13918 40898 13970 40910
rect 28478 40962 28530 40974
rect 28478 40898 28530 40910
rect 39790 40962 39842 40974
rect 39790 40898 39842 40910
rect 1344 40794 44576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 44576 40794
rect 1344 40708 44576 40742
rect 6302 40626 6354 40638
rect 6302 40562 6354 40574
rect 10446 40626 10498 40638
rect 10446 40562 10498 40574
rect 32622 40626 32674 40638
rect 32622 40562 32674 40574
rect 10222 40514 10274 40526
rect 34178 40462 34190 40514
rect 34242 40462 34254 40514
rect 10222 40450 10274 40462
rect 10110 40402 10162 40414
rect 17614 40402 17666 40414
rect 3042 40350 3054 40402
rect 3106 40350 3118 40402
rect 10770 40350 10782 40402
rect 10834 40350 10846 40402
rect 14018 40350 14030 40402
rect 14082 40350 14094 40402
rect 10110 40338 10162 40350
rect 17614 40338 17666 40350
rect 20078 40402 20130 40414
rect 31838 40402 31890 40414
rect 36878 40402 36930 40414
rect 20290 40350 20302 40402
rect 20354 40350 20366 40402
rect 25330 40350 25342 40402
rect 25394 40350 25406 40402
rect 28466 40350 28478 40402
rect 28530 40350 28542 40402
rect 29250 40350 29262 40402
rect 29314 40350 29326 40402
rect 33394 40350 33406 40402
rect 33458 40350 33470 40402
rect 20078 40338 20130 40350
rect 31838 40338 31890 40350
rect 36878 40338 36930 40350
rect 3714 40238 3726 40290
rect 3778 40238 3790 40290
rect 5842 40238 5854 40290
rect 5906 40238 5918 40290
rect 11442 40238 11454 40290
rect 11506 40238 11518 40290
rect 13570 40238 13582 40290
rect 13634 40238 13646 40290
rect 14690 40238 14702 40290
rect 14754 40238 14766 40290
rect 16818 40238 16830 40290
rect 16882 40238 16894 40290
rect 21074 40238 21086 40290
rect 21138 40238 21150 40290
rect 23202 40238 23214 40290
rect 23266 40238 23278 40290
rect 26002 40238 26014 40290
rect 26066 40238 26078 40290
rect 28130 40238 28142 40290
rect 28194 40238 28206 40290
rect 31378 40238 31390 40290
rect 31442 40238 31454 40290
rect 36306 40238 36318 40290
rect 36370 40238 36382 40290
rect 1344 40010 44576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 44576 40010
rect 1344 39924 44576 39958
rect 9102 39842 9154 39854
rect 9102 39778 9154 39790
rect 6414 39730 6466 39742
rect 6414 39666 6466 39678
rect 11342 39730 11394 39742
rect 11342 39666 11394 39678
rect 17054 39730 17106 39742
rect 34974 39730 35026 39742
rect 20290 39678 20302 39730
rect 20354 39678 20366 39730
rect 34402 39678 34414 39730
rect 34466 39678 34478 39730
rect 17054 39666 17106 39678
rect 34974 39666 35026 39678
rect 37998 39730 38050 39742
rect 38322 39678 38334 39730
rect 38386 39678 38398 39730
rect 37998 39666 38050 39678
rect 6974 39618 7026 39630
rect 6974 39554 7026 39566
rect 7758 39618 7810 39630
rect 7758 39554 7810 39566
rect 7982 39618 8034 39630
rect 7982 39554 8034 39566
rect 9214 39618 9266 39630
rect 9214 39554 9266 39566
rect 9662 39618 9714 39630
rect 9662 39554 9714 39566
rect 10222 39618 10274 39630
rect 10222 39554 10274 39566
rect 10782 39618 10834 39630
rect 10782 39554 10834 39566
rect 11230 39618 11282 39630
rect 11230 39554 11282 39566
rect 11790 39618 11842 39630
rect 41470 39618 41522 39630
rect 17490 39566 17502 39618
rect 17554 39566 17566 39618
rect 31490 39566 31502 39618
rect 31554 39566 31566 39618
rect 41122 39566 41134 39618
rect 41186 39566 41198 39618
rect 11790 39554 11842 39566
rect 41470 39554 41522 39566
rect 41806 39618 41858 39630
rect 41806 39554 41858 39566
rect 7646 39506 7698 39518
rect 7646 39442 7698 39454
rect 9774 39506 9826 39518
rect 9774 39442 9826 39454
rect 11902 39506 11954 39518
rect 11902 39442 11954 39454
rect 13918 39506 13970 39518
rect 13918 39442 13970 39454
rect 14254 39506 14306 39518
rect 41694 39506 41746 39518
rect 18162 39454 18174 39506
rect 18226 39454 18238 39506
rect 32162 39454 32174 39506
rect 32226 39454 32238 39506
rect 40450 39454 40462 39506
rect 40514 39454 40526 39506
rect 14254 39442 14306 39454
rect 41694 39442 41746 39454
rect 42142 39506 42194 39518
rect 42142 39442 42194 39454
rect 6302 39394 6354 39406
rect 6302 39330 6354 39342
rect 6526 39394 6578 39406
rect 6526 39330 6578 39342
rect 7310 39394 7362 39406
rect 7310 39330 7362 39342
rect 7534 39394 7586 39406
rect 7534 39330 7586 39342
rect 8318 39394 8370 39406
rect 8318 39330 8370 39342
rect 8542 39394 8594 39406
rect 8542 39330 8594 39342
rect 8654 39394 8706 39406
rect 8654 39330 8706 39342
rect 9102 39394 9154 39406
rect 9102 39330 9154 39342
rect 9886 39394 9938 39406
rect 9886 39330 9938 39342
rect 11454 39394 11506 39406
rect 11454 39330 11506 39342
rect 12126 39394 12178 39406
rect 12126 39330 12178 39342
rect 28254 39394 28306 39406
rect 28254 39330 28306 39342
rect 1344 39226 44576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 44576 39226
rect 1344 39140 44576 39174
rect 5182 39058 5234 39070
rect 5182 38994 5234 39006
rect 7982 39058 8034 39070
rect 7982 38994 8034 39006
rect 9550 39058 9602 39070
rect 39230 39058 39282 39070
rect 12114 39006 12126 39058
rect 12178 39006 12190 39058
rect 9550 38994 9602 39006
rect 39230 38994 39282 39006
rect 40350 39058 40402 39070
rect 40350 38994 40402 39006
rect 7646 38946 7698 38958
rect 2594 38894 2606 38946
rect 2658 38894 2670 38946
rect 7646 38882 7698 38894
rect 7758 38946 7810 38958
rect 7758 38882 7810 38894
rect 8878 38946 8930 38958
rect 11566 38946 11618 38958
rect 10770 38894 10782 38946
rect 10834 38894 10846 38946
rect 8878 38882 8930 38894
rect 11566 38882 11618 38894
rect 40126 38946 40178 38958
rect 40126 38882 40178 38894
rect 8990 38834 9042 38846
rect 1922 38782 1934 38834
rect 1986 38782 1998 38834
rect 8990 38770 9042 38782
rect 9886 38834 9938 38846
rect 9886 38770 9938 38782
rect 10222 38834 10274 38846
rect 10222 38770 10274 38782
rect 11790 38834 11842 38846
rect 11790 38770 11842 38782
rect 40014 38834 40066 38846
rect 41122 38782 41134 38834
rect 41186 38782 41198 38834
rect 40014 38770 40066 38782
rect 39678 38722 39730 38734
rect 4722 38670 4734 38722
rect 4786 38670 4798 38722
rect 41906 38670 41918 38722
rect 41970 38670 41982 38722
rect 44034 38670 44046 38722
rect 44098 38670 44110 38722
rect 39678 38658 39730 38670
rect 10446 38610 10498 38622
rect 10446 38546 10498 38558
rect 1344 38442 44576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 44576 38442
rect 1344 38356 44576 38390
rect 37874 38222 37886 38274
rect 37938 38222 37950 38274
rect 10110 38162 10162 38174
rect 42030 38162 42082 38174
rect 38322 38110 38334 38162
rect 38386 38110 38398 38162
rect 10110 38098 10162 38110
rect 42030 38098 42082 38110
rect 9662 38050 9714 38062
rect 9662 37986 9714 37998
rect 10222 38050 10274 38062
rect 25790 38050 25842 38062
rect 40798 38050 40850 38062
rect 10546 37998 10558 38050
rect 10610 37998 10622 38050
rect 25554 37998 25566 38050
rect 25618 37998 25630 38050
rect 38098 37998 38110 38050
rect 38162 37998 38174 38050
rect 10222 37986 10274 37998
rect 25790 37986 25842 37998
rect 40798 37986 40850 37998
rect 41022 38050 41074 38062
rect 41022 37986 41074 37998
rect 41358 38050 41410 38062
rect 41358 37986 41410 37998
rect 41806 38050 41858 38062
rect 41806 37986 41858 37998
rect 24894 37938 24946 37950
rect 11442 37886 11454 37938
rect 11506 37886 11518 37938
rect 24894 37874 24946 37886
rect 40462 37938 40514 37950
rect 40462 37874 40514 37886
rect 41582 37938 41634 37950
rect 41582 37874 41634 37886
rect 42142 37938 42194 37950
rect 42142 37874 42194 37886
rect 42366 37938 42418 37950
rect 42366 37874 42418 37886
rect 42702 37938 42754 37950
rect 42702 37874 42754 37886
rect 43150 37938 43202 37950
rect 43150 37874 43202 37886
rect 12126 37826 12178 37838
rect 12126 37762 12178 37774
rect 26350 37826 26402 37838
rect 26350 37762 26402 37774
rect 39790 37826 39842 37838
rect 39790 37762 39842 37774
rect 40238 37826 40290 37838
rect 40238 37762 40290 37774
rect 40574 37826 40626 37838
rect 40574 37762 40626 37774
rect 41134 37826 41186 37838
rect 41134 37762 41186 37774
rect 42590 37826 42642 37838
rect 42590 37762 42642 37774
rect 1344 37658 44576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 44576 37658
rect 1344 37572 44576 37606
rect 19742 37490 19794 37502
rect 6850 37438 6862 37490
rect 6914 37438 6926 37490
rect 19742 37426 19794 37438
rect 30830 37378 30882 37390
rect 25554 37326 25566 37378
rect 25618 37326 25630 37378
rect 30830 37314 30882 37326
rect 25230 37266 25282 37278
rect 37774 37266 37826 37278
rect 7074 37214 7086 37266
rect 7138 37214 7150 37266
rect 20066 37214 20078 37266
rect 20130 37214 20142 37266
rect 24322 37214 24334 37266
rect 24386 37214 24398 37266
rect 27570 37214 27582 37266
rect 27634 37214 27646 37266
rect 34626 37214 34638 37266
rect 34690 37214 34702 37266
rect 25230 37202 25282 37214
rect 37774 37202 37826 37214
rect 23662 37154 23714 37166
rect 20850 37102 20862 37154
rect 20914 37102 20926 37154
rect 22978 37102 22990 37154
rect 23042 37102 23054 37154
rect 24546 37102 24558 37154
rect 24610 37102 24622 37154
rect 28242 37102 28254 37154
rect 28306 37102 28318 37154
rect 30370 37102 30382 37154
rect 30434 37102 30446 37154
rect 35298 37102 35310 37154
rect 35362 37102 35374 37154
rect 37426 37102 37438 37154
rect 37490 37102 37502 37154
rect 38210 37102 38222 37154
rect 38274 37102 38286 37154
rect 23662 37090 23714 37102
rect 1344 36874 44576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 44576 36874
rect 1344 36788 44576 36822
rect 21534 36706 21586 36718
rect 21534 36642 21586 36654
rect 21870 36706 21922 36718
rect 21870 36642 21922 36654
rect 24222 36706 24274 36718
rect 24222 36642 24274 36654
rect 27918 36706 27970 36718
rect 27918 36642 27970 36654
rect 27134 36594 27186 36606
rect 27134 36530 27186 36542
rect 37662 36594 37714 36606
rect 37662 36530 37714 36542
rect 17278 36482 17330 36494
rect 17278 36418 17330 36430
rect 17502 36482 17554 36494
rect 17502 36418 17554 36430
rect 24334 36482 24386 36494
rect 24334 36418 24386 36430
rect 26798 36482 26850 36494
rect 26798 36418 26850 36430
rect 29486 36482 29538 36494
rect 31278 36482 31330 36494
rect 30818 36430 30830 36482
rect 30882 36430 30894 36482
rect 29486 36418 29538 36430
rect 31278 36418 31330 36430
rect 7086 36370 7138 36382
rect 7086 36306 7138 36318
rect 15598 36370 15650 36382
rect 18062 36370 18114 36382
rect 16930 36318 16942 36370
rect 16994 36318 17006 36370
rect 15598 36306 15650 36318
rect 18062 36306 18114 36318
rect 26910 36370 26962 36382
rect 26910 36306 26962 36318
rect 27246 36370 27298 36382
rect 27246 36306 27298 36318
rect 27582 36370 27634 36382
rect 27582 36306 27634 36318
rect 27806 36370 27858 36382
rect 30382 36370 30434 36382
rect 29138 36318 29150 36370
rect 29202 36318 29214 36370
rect 27806 36306 27858 36318
rect 30382 36306 30434 36318
rect 7198 36258 7250 36270
rect 7198 36194 7250 36206
rect 10446 36258 10498 36270
rect 10446 36194 10498 36206
rect 15486 36258 15538 36270
rect 15486 36194 15538 36206
rect 17726 36258 17778 36270
rect 17726 36194 17778 36206
rect 17950 36258 18002 36270
rect 17950 36194 18002 36206
rect 20862 36258 20914 36270
rect 20862 36194 20914 36206
rect 21646 36258 21698 36270
rect 21646 36194 21698 36206
rect 24222 36258 24274 36270
rect 24222 36194 24274 36206
rect 28366 36258 28418 36270
rect 28366 36194 28418 36206
rect 1344 36090 44576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 44576 36090
rect 1344 36004 44576 36038
rect 19070 35922 19122 35934
rect 10658 35870 10670 35922
rect 10722 35870 10734 35922
rect 19070 35858 19122 35870
rect 41358 35922 41410 35934
rect 41358 35858 41410 35870
rect 7646 35810 7698 35822
rect 2594 35758 2606 35810
rect 2658 35758 2670 35810
rect 7646 35746 7698 35758
rect 11118 35810 11170 35822
rect 11118 35746 11170 35758
rect 11230 35810 11282 35822
rect 11230 35746 11282 35758
rect 14702 35810 14754 35822
rect 14702 35746 14754 35758
rect 17950 35810 18002 35822
rect 17950 35746 18002 35758
rect 18622 35810 18674 35822
rect 18622 35746 18674 35758
rect 19630 35810 19682 35822
rect 19630 35746 19682 35758
rect 41806 35810 41858 35822
rect 41806 35746 41858 35758
rect 41918 35810 41970 35822
rect 41918 35746 41970 35758
rect 7982 35698 8034 35710
rect 1922 35646 1934 35698
rect 1986 35646 1998 35698
rect 7982 35634 8034 35646
rect 11342 35698 11394 35710
rect 15262 35698 15314 35710
rect 14914 35646 14926 35698
rect 14978 35646 14990 35698
rect 11342 35634 11394 35646
rect 15262 35634 15314 35646
rect 15710 35698 15762 35710
rect 15710 35634 15762 35646
rect 16382 35698 16434 35710
rect 17838 35698 17890 35710
rect 18734 35698 18786 35710
rect 17378 35646 17390 35698
rect 17442 35646 17454 35698
rect 18162 35646 18174 35698
rect 18226 35646 18238 35698
rect 16382 35634 16434 35646
rect 17838 35634 17890 35646
rect 18734 35634 18786 35646
rect 19182 35698 19234 35710
rect 20526 35698 20578 35710
rect 20066 35646 20078 35698
rect 20130 35646 20142 35698
rect 19182 35634 19234 35646
rect 20526 35634 20578 35646
rect 41582 35698 41634 35710
rect 41582 35634 41634 35646
rect 5182 35586 5234 35598
rect 4722 35534 4734 35586
rect 4786 35534 4798 35586
rect 5182 35522 5234 35534
rect 10334 35586 10386 35598
rect 16258 35534 16270 35586
rect 16322 35534 16334 35586
rect 10334 35522 10386 35534
rect 10110 35474 10162 35486
rect 9762 35422 9774 35474
rect 9826 35422 9838 35474
rect 10110 35410 10162 35422
rect 14590 35474 14642 35486
rect 14590 35410 14642 35422
rect 15934 35474 15986 35486
rect 15934 35410 15986 35422
rect 16494 35474 16546 35486
rect 16494 35410 16546 35422
rect 18622 35474 18674 35486
rect 18622 35410 18674 35422
rect 1344 35306 44576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 44576 35306
rect 1344 35220 44576 35254
rect 17166 35138 17218 35150
rect 17166 35074 17218 35086
rect 17726 35138 17778 35150
rect 17726 35074 17778 35086
rect 18062 35138 18114 35150
rect 18062 35074 18114 35086
rect 9886 35026 9938 35038
rect 9886 34962 9938 34974
rect 10782 35026 10834 35038
rect 10782 34962 10834 34974
rect 11342 35026 11394 35038
rect 11342 34962 11394 34974
rect 15598 35026 15650 35038
rect 15598 34962 15650 34974
rect 16830 35026 16882 35038
rect 40574 35026 40626 35038
rect 33058 34974 33070 35026
rect 33122 34974 33134 35026
rect 43810 34974 43822 35026
rect 43874 34974 43886 35026
rect 16830 34962 16882 34974
rect 40574 34962 40626 34974
rect 8766 34914 8818 34926
rect 8766 34850 8818 34862
rect 9326 34914 9378 34926
rect 9326 34850 9378 34862
rect 10222 34914 10274 34926
rect 10222 34850 10274 34862
rect 11118 34914 11170 34926
rect 11118 34850 11170 34862
rect 11566 34914 11618 34926
rect 11566 34850 11618 34862
rect 11678 34914 11730 34926
rect 15374 34914 15426 34926
rect 14690 34862 14702 34914
rect 14754 34862 14766 34914
rect 11678 34850 11730 34862
rect 15374 34850 15426 34862
rect 25566 34914 25618 34926
rect 33518 34914 33570 34926
rect 30258 34862 30270 34914
rect 30322 34862 30334 34914
rect 41010 34862 41022 34914
rect 41074 34862 41086 34914
rect 25566 34850 25618 34862
rect 33518 34850 33570 34862
rect 14366 34802 14418 34814
rect 14366 34738 14418 34750
rect 14926 34802 14978 34814
rect 14926 34738 14978 34750
rect 15934 34802 15986 34814
rect 15934 34738 15986 34750
rect 17390 34802 17442 34814
rect 17390 34738 17442 34750
rect 25790 34802 25842 34814
rect 30930 34750 30942 34802
rect 30994 34750 31006 34802
rect 41682 34750 41694 34802
rect 41746 34750 41758 34802
rect 25790 34738 25842 34750
rect 9774 34690 9826 34702
rect 9090 34638 9102 34690
rect 9154 34638 9166 34690
rect 9774 34626 9826 34638
rect 9998 34690 10050 34702
rect 9998 34626 10050 34638
rect 10670 34690 10722 34702
rect 10670 34626 10722 34638
rect 10894 34690 10946 34702
rect 10894 34626 10946 34638
rect 12350 34690 12402 34702
rect 12350 34626 12402 34638
rect 14142 34690 14194 34702
rect 14142 34626 14194 34638
rect 14478 34690 14530 34702
rect 14478 34626 14530 34638
rect 15710 34690 15762 34702
rect 15710 34626 15762 34638
rect 17838 34690 17890 34702
rect 17838 34626 17890 34638
rect 25678 34690 25730 34702
rect 25678 34626 25730 34638
rect 26014 34690 26066 34702
rect 26014 34626 26066 34638
rect 27134 34690 27186 34702
rect 27134 34626 27186 34638
rect 1344 34522 44576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 44576 34522
rect 1344 34436 44576 34470
rect 10110 34354 10162 34366
rect 26574 34354 26626 34366
rect 14690 34302 14702 34354
rect 14754 34302 14766 34354
rect 10110 34290 10162 34302
rect 26574 34290 26626 34302
rect 26798 34354 26850 34366
rect 26798 34290 26850 34302
rect 27358 34354 27410 34366
rect 27358 34290 27410 34302
rect 27694 34354 27746 34366
rect 27694 34290 27746 34302
rect 38894 34354 38946 34366
rect 38894 34290 38946 34302
rect 9662 34242 9714 34254
rect 4946 34190 4958 34242
rect 5010 34190 5022 34242
rect 9662 34178 9714 34190
rect 27918 34242 27970 34254
rect 31826 34190 31838 34242
rect 31890 34190 31902 34242
rect 27918 34178 27970 34190
rect 9550 34130 9602 34142
rect 14142 34130 14194 34142
rect 27470 34130 27522 34142
rect 4274 34078 4286 34130
rect 4338 34078 4350 34130
rect 10546 34078 10558 34130
rect 10610 34078 10622 34130
rect 26338 34078 26350 34130
rect 26402 34078 26414 34130
rect 27122 34078 27134 34130
rect 27186 34078 27198 34130
rect 9550 34066 9602 34078
rect 14142 34066 14194 34078
rect 27470 34066 27522 34078
rect 28030 34130 28082 34142
rect 32050 34078 32062 34130
rect 32114 34078 32126 34130
rect 38322 34078 38334 34130
rect 38386 34078 38398 34130
rect 42242 34078 42254 34130
rect 42306 34078 42318 34130
rect 28030 34066 28082 34078
rect 7534 34018 7586 34030
rect 11454 34018 11506 34030
rect 7074 33966 7086 34018
rect 7138 33966 7150 34018
rect 10882 33966 10894 34018
rect 10946 33966 10958 34018
rect 26674 33966 26686 34018
rect 26738 33966 26750 34018
rect 35522 33966 35534 34018
rect 35586 33966 35598 34018
rect 37650 33966 37662 34018
rect 37714 33966 37726 34018
rect 41906 33966 41918 34018
rect 41970 33966 41982 34018
rect 7534 33954 7586 33966
rect 11454 33954 11506 33966
rect 14366 33906 14418 33918
rect 41458 33854 41470 33906
rect 41522 33854 41534 33906
rect 14366 33842 14418 33854
rect 1344 33738 44576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 44576 33738
rect 1344 33652 44576 33686
rect 30830 33570 30882 33582
rect 30830 33506 30882 33518
rect 10222 33458 10274 33470
rect 10222 33394 10274 33406
rect 23102 33458 23154 33470
rect 23102 33394 23154 33406
rect 25118 33458 25170 33470
rect 25118 33394 25170 33406
rect 35870 33458 35922 33470
rect 35870 33394 35922 33406
rect 37102 33458 37154 33470
rect 37102 33394 37154 33406
rect 41806 33458 41858 33470
rect 41806 33394 41858 33406
rect 11342 33346 11394 33358
rect 27022 33346 27074 33358
rect 31390 33346 31442 33358
rect 23762 33294 23774 33346
rect 23826 33294 23838 33346
rect 30930 33294 30942 33346
rect 30994 33294 31006 33346
rect 11342 33282 11394 33294
rect 27022 33282 27074 33294
rect 31390 33282 31442 33294
rect 32958 33346 33010 33358
rect 32958 33282 33010 33294
rect 36094 33346 36146 33358
rect 36094 33282 36146 33294
rect 37326 33346 37378 33358
rect 37326 33282 37378 33294
rect 37774 33346 37826 33358
rect 37774 33282 37826 33294
rect 41694 33346 41746 33358
rect 41694 33282 41746 33294
rect 42254 33346 42306 33358
rect 42254 33282 42306 33294
rect 26686 33234 26738 33246
rect 24658 33182 24670 33234
rect 24722 33182 24734 33234
rect 26686 33170 26738 33182
rect 30718 33234 30770 33246
rect 30718 33170 30770 33182
rect 31614 33234 31666 33246
rect 31614 33170 31666 33182
rect 31726 33234 31778 33246
rect 31726 33170 31778 33182
rect 32622 33234 32674 33246
rect 32622 33170 32674 33182
rect 32734 33234 32786 33246
rect 32734 33170 32786 33182
rect 35758 33234 35810 33246
rect 35758 33170 35810 33182
rect 36318 33234 36370 33246
rect 36318 33170 36370 33182
rect 36990 33234 37042 33246
rect 36990 33170 37042 33182
rect 37550 33234 37602 33246
rect 37550 33170 37602 33182
rect 38110 33234 38162 33246
rect 38110 33170 38162 33182
rect 42030 33234 42082 33246
rect 42030 33170 42082 33182
rect 26798 33122 26850 33134
rect 11666 33070 11678 33122
rect 11730 33070 11742 33122
rect 26798 33058 26850 33070
rect 27470 33122 27522 33134
rect 27470 33058 27522 33070
rect 31166 33122 31218 33134
rect 31166 33058 31218 33070
rect 34750 33122 34802 33134
rect 34750 33058 34802 33070
rect 35086 33122 35138 33134
rect 37998 33122 38050 33134
rect 35410 33070 35422 33122
rect 35474 33070 35486 33122
rect 35086 33058 35138 33070
rect 37998 33058 38050 33070
rect 1344 32954 44576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 44576 32954
rect 1344 32868 44576 32902
rect 19630 32786 19682 32798
rect 19630 32722 19682 32734
rect 30830 32786 30882 32798
rect 30830 32722 30882 32734
rect 31054 32786 31106 32798
rect 31054 32722 31106 32734
rect 31502 32786 31554 32798
rect 31502 32722 31554 32734
rect 32398 32786 32450 32798
rect 32398 32722 32450 32734
rect 36878 32786 36930 32798
rect 36878 32722 36930 32734
rect 37102 32786 37154 32798
rect 37102 32722 37154 32734
rect 37214 32786 37266 32798
rect 37214 32722 37266 32734
rect 42142 32786 42194 32798
rect 42142 32722 42194 32734
rect 37438 32674 37490 32686
rect 15474 32622 15486 32674
rect 15538 32622 15550 32674
rect 37438 32610 37490 32622
rect 41918 32674 41970 32686
rect 41918 32610 41970 32622
rect 24110 32562 24162 32574
rect 15250 32510 15262 32562
rect 15314 32510 15326 32562
rect 19954 32510 19966 32562
rect 20018 32510 20030 32562
rect 23874 32510 23886 32562
rect 23938 32510 23950 32562
rect 24110 32498 24162 32510
rect 26574 32562 26626 32574
rect 26574 32498 26626 32510
rect 31166 32562 31218 32574
rect 32062 32562 32114 32574
rect 31714 32510 31726 32562
rect 31778 32510 31790 32562
rect 31166 32498 31218 32510
rect 32062 32498 32114 32510
rect 32286 32562 32338 32574
rect 32286 32498 32338 32510
rect 36766 32562 36818 32574
rect 36766 32498 36818 32510
rect 37550 32562 37602 32574
rect 37550 32498 37602 32510
rect 41806 32562 41858 32574
rect 41806 32498 41858 32510
rect 23214 32450 23266 32462
rect 27022 32450 27074 32462
rect 20738 32398 20750 32450
rect 20802 32398 20814 32450
rect 22866 32398 22878 32450
rect 22930 32398 22942 32450
rect 26114 32398 26126 32450
rect 26178 32398 26190 32450
rect 23214 32386 23266 32398
rect 27022 32386 27074 32398
rect 31838 32450 31890 32462
rect 31838 32386 31890 32398
rect 32398 32338 32450 32350
rect 32398 32274 32450 32286
rect 1344 32170 44576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 44576 32170
rect 1344 32084 44576 32118
rect 21534 32002 21586 32014
rect 21534 31938 21586 31950
rect 21870 32002 21922 32014
rect 21870 31938 21922 31950
rect 25678 31890 25730 31902
rect 5058 31838 5070 31890
rect 5122 31838 5134 31890
rect 25678 31826 25730 31838
rect 26238 31890 26290 31902
rect 26238 31826 26290 31838
rect 27134 31890 27186 31902
rect 27134 31826 27186 31838
rect 27582 31890 27634 31902
rect 27582 31826 27634 31838
rect 12910 31778 12962 31790
rect 14030 31778 14082 31790
rect 25790 31778 25842 31790
rect 2146 31726 2158 31778
rect 2210 31726 2222 31778
rect 13570 31726 13582 31778
rect 13634 31726 13646 31778
rect 19954 31726 19966 31778
rect 20018 31726 20030 31778
rect 12910 31714 12962 31726
rect 14030 31714 14082 31726
rect 25790 31714 25842 31726
rect 26686 31778 26738 31790
rect 30034 31726 30046 31778
rect 30098 31726 30110 31778
rect 26686 31714 26738 31726
rect 25342 31666 25394 31678
rect 2930 31614 2942 31666
rect 2994 31614 3006 31666
rect 15138 31614 15150 31666
rect 15202 31614 15214 31666
rect 25342 31602 25394 31614
rect 26126 31666 26178 31678
rect 26126 31602 26178 31614
rect 26462 31666 26514 31678
rect 40338 31614 40350 31666
rect 40402 31614 40414 31666
rect 26462 31602 26514 31614
rect 5742 31554 5794 31566
rect 5742 31490 5794 31502
rect 20750 31554 20802 31566
rect 20750 31490 20802 31502
rect 21646 31554 21698 31566
rect 21646 31490 21698 31502
rect 25566 31554 25618 31566
rect 30718 31554 30770 31566
rect 30258 31502 30270 31554
rect 30322 31502 30334 31554
rect 25566 31490 25618 31502
rect 30718 31490 30770 31502
rect 36430 31554 36482 31566
rect 36430 31490 36482 31502
rect 36990 31554 37042 31566
rect 39678 31554 39730 31566
rect 37314 31502 37326 31554
rect 37378 31502 37390 31554
rect 36990 31490 37042 31502
rect 39678 31490 39730 31502
rect 40014 31554 40066 31566
rect 40014 31490 40066 31502
rect 1344 31386 44576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 44576 31386
rect 1344 31300 44576 31334
rect 4174 31218 4226 31230
rect 4174 31154 4226 31166
rect 16270 31218 16322 31230
rect 16270 31154 16322 31166
rect 31726 31218 31778 31230
rect 31726 31154 31778 31166
rect 41470 31218 41522 31230
rect 41470 31154 41522 31166
rect 30718 31106 30770 31118
rect 30718 31042 30770 31054
rect 31502 31106 31554 31118
rect 40014 31106 40066 31118
rect 36642 31054 36654 31106
rect 36706 31054 36718 31106
rect 31502 31042 31554 31054
rect 40014 31042 40066 31054
rect 40126 31106 40178 31118
rect 40126 31042 40178 31054
rect 41806 31106 41858 31118
rect 41806 31042 41858 31054
rect 16494 30994 16546 31006
rect 17950 30994 18002 31006
rect 6066 30942 6078 30994
rect 6130 30942 6142 30994
rect 15922 30942 15934 30994
rect 15986 30942 15998 30994
rect 16818 30942 16830 30994
rect 16882 30942 16894 30994
rect 16494 30930 16546 30942
rect 17950 30930 18002 30942
rect 30606 30994 30658 31006
rect 30606 30930 30658 30942
rect 30942 30994 30994 31006
rect 30942 30930 30994 30942
rect 31390 30994 31442 31006
rect 31390 30930 31442 30942
rect 32510 30994 32562 31006
rect 40350 30994 40402 31006
rect 33394 30942 33406 30994
rect 33458 30942 33470 30994
rect 32510 30930 32562 30942
rect 40350 30930 40402 30942
rect 41134 30994 41186 31006
rect 41134 30930 41186 30942
rect 41582 30994 41634 31006
rect 41582 30930 41634 30942
rect 4286 30882 4338 30894
rect 9662 30882 9714 30894
rect 16382 30882 16434 30894
rect 6850 30830 6862 30882
rect 6914 30830 6926 30882
rect 8978 30830 8990 30882
rect 9042 30830 9054 30882
rect 10882 30830 10894 30882
rect 10946 30830 10958 30882
rect 4286 30818 4338 30830
rect 9662 30818 9714 30830
rect 16382 30818 16434 30830
rect 17502 30882 17554 30894
rect 17502 30818 17554 30830
rect 20190 30882 20242 30894
rect 20190 30818 20242 30830
rect 1344 30602 44576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 44576 30602
rect 1344 30516 44576 30550
rect 15822 30434 15874 30446
rect 15822 30370 15874 30382
rect 9538 30270 9550 30322
rect 9602 30270 9614 30322
rect 16146 30270 16158 30322
rect 16210 30270 16222 30322
rect 41458 30270 41470 30322
rect 41522 30270 41534 30322
rect 43586 30270 43598 30322
rect 43650 30270 43662 30322
rect 13022 30210 13074 30222
rect 19630 30210 19682 30222
rect 12450 30158 12462 30210
rect 12514 30158 12526 30210
rect 14914 30158 14926 30210
rect 14978 30158 14990 30210
rect 18946 30158 18958 30210
rect 19010 30158 19022 30210
rect 13022 30146 13074 30158
rect 19630 30146 19682 30158
rect 28590 30210 28642 30222
rect 35310 30210 35362 30222
rect 30146 30158 30158 30210
rect 30210 30158 30222 30210
rect 28590 30146 28642 30158
rect 35310 30146 35362 30158
rect 37438 30210 37490 30222
rect 40674 30158 40686 30210
rect 40738 30158 40750 30210
rect 37438 30146 37490 30158
rect 15710 30098 15762 30110
rect 34974 30098 35026 30110
rect 36990 30098 37042 30110
rect 11666 30046 11678 30098
rect 11730 30046 11742 30098
rect 18274 30046 18286 30098
rect 18338 30046 18350 30098
rect 33506 30046 33518 30098
rect 33570 30046 33582 30098
rect 35970 30046 35982 30098
rect 36034 30046 36046 30098
rect 15710 30034 15762 30046
rect 34974 30034 35026 30046
rect 36990 30034 37042 30046
rect 37326 30098 37378 30110
rect 37326 30034 37378 30046
rect 39118 30098 39170 30110
rect 39118 30034 39170 30046
rect 39342 30098 39394 30110
rect 39342 30034 39394 30046
rect 39454 30098 39506 30110
rect 39454 30034 39506 30046
rect 15150 29986 15202 29998
rect 15150 29922 15202 29934
rect 15598 29986 15650 29998
rect 15598 29922 15650 29934
rect 35198 29986 35250 29998
rect 35198 29922 35250 29934
rect 35646 29986 35698 29998
rect 35646 29922 35698 29934
rect 36430 29986 36482 29998
rect 36430 29922 36482 29934
rect 37102 29986 37154 29998
rect 37102 29922 37154 29934
rect 40350 29986 40402 29998
rect 40350 29922 40402 29934
rect 1344 29818 44576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 44576 29818
rect 1344 29732 44576 29766
rect 5854 29650 5906 29662
rect 5854 29586 5906 29598
rect 11230 29650 11282 29662
rect 11230 29586 11282 29598
rect 11902 29650 11954 29662
rect 11902 29586 11954 29598
rect 22990 29650 23042 29662
rect 22990 29586 23042 29598
rect 24110 29650 24162 29662
rect 24110 29586 24162 29598
rect 32062 29650 32114 29662
rect 32062 29586 32114 29598
rect 38222 29650 38274 29662
rect 38222 29586 38274 29598
rect 41470 29650 41522 29662
rect 41470 29586 41522 29598
rect 41694 29538 41746 29550
rect 23202 29486 23214 29538
rect 23266 29486 23278 29538
rect 36978 29486 36990 29538
rect 37042 29486 37054 29538
rect 41694 29474 41746 29486
rect 41806 29538 41858 29550
rect 41806 29474 41858 29486
rect 1922 29374 1934 29426
rect 1986 29374 1998 29426
rect 11442 29374 11454 29426
rect 11506 29374 11518 29426
rect 14354 29374 14366 29426
rect 14418 29374 14430 29426
rect 23426 29374 23438 29426
rect 23490 29374 23502 29426
rect 28802 29374 28814 29426
rect 28866 29374 28878 29426
rect 37762 29374 37774 29426
rect 37826 29374 37838 29426
rect 5518 29314 5570 29326
rect 2594 29262 2606 29314
rect 2658 29262 2670 29314
rect 4834 29262 4846 29314
rect 4898 29262 4910 29314
rect 5518 29250 5570 29262
rect 23998 29314 24050 29326
rect 29474 29262 29486 29314
rect 29538 29262 29550 29314
rect 31602 29262 31614 29314
rect 31666 29262 31678 29314
rect 34850 29262 34862 29314
rect 34914 29262 34926 29314
rect 23998 29250 24050 29262
rect 11118 29202 11170 29214
rect 13906 29150 13918 29202
rect 13970 29150 13982 29202
rect 11118 29138 11170 29150
rect 1344 29034 44576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 44576 29034
rect 1344 28948 44576 28982
rect 4510 28866 4562 28878
rect 29262 28866 29314 28878
rect 15922 28814 15934 28866
rect 15986 28814 15998 28866
rect 4510 28802 4562 28814
rect 29262 28802 29314 28814
rect 29822 28866 29874 28878
rect 29822 28802 29874 28814
rect 30382 28866 30434 28878
rect 30382 28802 30434 28814
rect 5742 28754 5794 28766
rect 5742 28690 5794 28702
rect 6974 28754 7026 28766
rect 27022 28754 27074 28766
rect 15138 28702 15150 28754
rect 15202 28702 15214 28754
rect 6974 28690 7026 28702
rect 27022 28690 27074 28702
rect 11902 28642 11954 28654
rect 6402 28590 6414 28642
rect 6466 28590 6478 28642
rect 11554 28590 11566 28642
rect 11618 28590 11630 28642
rect 11902 28578 11954 28590
rect 12350 28642 12402 28654
rect 12350 28578 12402 28590
rect 12462 28642 12514 28654
rect 12462 28578 12514 28590
rect 12686 28642 12738 28654
rect 12686 28578 12738 28590
rect 12910 28642 12962 28654
rect 12910 28578 12962 28590
rect 15710 28642 15762 28654
rect 15710 28578 15762 28590
rect 16270 28642 16322 28654
rect 16270 28578 16322 28590
rect 16494 28642 16546 28654
rect 16494 28578 16546 28590
rect 16718 28642 16770 28654
rect 16718 28578 16770 28590
rect 17278 28642 17330 28654
rect 17278 28578 17330 28590
rect 21310 28642 21362 28654
rect 21310 28578 21362 28590
rect 21534 28642 21586 28654
rect 21534 28578 21586 28590
rect 21982 28642 22034 28654
rect 21982 28578 22034 28590
rect 22318 28642 22370 28654
rect 22318 28578 22370 28590
rect 26574 28642 26626 28654
rect 26574 28578 26626 28590
rect 29598 28642 29650 28654
rect 31950 28642 32002 28654
rect 30930 28590 30942 28642
rect 30994 28590 31006 28642
rect 29598 28578 29650 28590
rect 31950 28578 32002 28590
rect 32510 28642 32562 28654
rect 32510 28578 32562 28590
rect 32846 28642 32898 28654
rect 32846 28578 32898 28590
rect 34638 28642 34690 28654
rect 34638 28578 34690 28590
rect 35982 28642 36034 28654
rect 35982 28578 36034 28590
rect 5070 28530 5122 28542
rect 5070 28466 5122 28478
rect 5854 28530 5906 28542
rect 5854 28466 5906 28478
rect 5966 28530 6018 28542
rect 5966 28466 6018 28478
rect 17390 28530 17442 28542
rect 17390 28466 17442 28478
rect 26238 28530 26290 28542
rect 26238 28466 26290 28478
rect 29374 28530 29426 28542
rect 29374 28466 29426 28478
rect 29934 28530 29986 28542
rect 32734 28530 32786 28542
rect 32274 28478 32286 28530
rect 32338 28478 32350 28530
rect 36306 28478 36318 28530
rect 36370 28478 36382 28530
rect 29934 28466 29986 28478
rect 32734 28466 32786 28478
rect 4622 28418 4674 28430
rect 4622 28354 4674 28366
rect 4846 28418 4898 28430
rect 4846 28354 4898 28366
rect 5630 28418 5682 28430
rect 5630 28354 5682 28366
rect 15150 28418 15202 28430
rect 15150 28354 15202 28366
rect 15374 28418 15426 28430
rect 15374 28354 15426 28366
rect 17166 28418 17218 28430
rect 17166 28354 17218 28366
rect 21758 28418 21810 28430
rect 21758 28354 21810 28366
rect 28590 28418 28642 28430
rect 28590 28354 28642 28366
rect 29262 28418 29314 28430
rect 29262 28354 29314 28366
rect 30158 28418 30210 28430
rect 30158 28354 30210 28366
rect 30494 28418 30546 28430
rect 30494 28354 30546 28366
rect 30718 28418 30770 28430
rect 34962 28366 34974 28418
rect 35026 28366 35038 28418
rect 30718 28354 30770 28366
rect 1344 28250 44576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 44576 28250
rect 1344 28164 44576 28198
rect 5406 28082 5458 28094
rect 5406 28018 5458 28030
rect 5630 28082 5682 28094
rect 5630 28018 5682 28030
rect 11454 28082 11506 28094
rect 11454 28018 11506 28030
rect 12350 28082 12402 28094
rect 12350 28018 12402 28030
rect 12574 28082 12626 28094
rect 12574 28018 12626 28030
rect 22878 28082 22930 28094
rect 22878 28018 22930 28030
rect 23662 28082 23714 28094
rect 23662 28018 23714 28030
rect 28590 28082 28642 28094
rect 28590 28018 28642 28030
rect 5742 27970 5794 27982
rect 5742 27906 5794 27918
rect 11902 27970 11954 27982
rect 23102 27970 23154 27982
rect 21858 27918 21870 27970
rect 21922 27918 21934 27970
rect 11902 27906 11954 27918
rect 23102 27906 23154 27918
rect 23214 27970 23266 27982
rect 41694 27970 41746 27982
rect 26002 27918 26014 27970
rect 26066 27918 26078 27970
rect 23214 27906 23266 27918
rect 41694 27906 41746 27918
rect 12686 27858 12738 27870
rect 30158 27858 30210 27870
rect 11666 27806 11678 27858
rect 11730 27806 11742 27858
rect 22642 27806 22654 27858
rect 22706 27806 22718 27858
rect 25330 27806 25342 27858
rect 25394 27806 25406 27858
rect 12686 27794 12738 27806
rect 30158 27794 30210 27806
rect 41582 27858 41634 27870
rect 41582 27794 41634 27806
rect 13134 27746 13186 27758
rect 42254 27746 42306 27758
rect 11442 27694 11454 27746
rect 11506 27694 11518 27746
rect 19730 27694 19742 27746
rect 19794 27694 19806 27746
rect 28130 27694 28142 27746
rect 28194 27694 28206 27746
rect 13134 27682 13186 27694
rect 42254 27682 42306 27694
rect 41694 27634 41746 27646
rect 41694 27570 41746 27582
rect 42142 27634 42194 27646
rect 42142 27570 42194 27582
rect 1344 27466 44576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 44576 27466
rect 1344 27380 44576 27414
rect 5966 27186 6018 27198
rect 12126 27186 12178 27198
rect 11330 27134 11342 27186
rect 11394 27134 11406 27186
rect 5966 27122 6018 27134
rect 12126 27122 12178 27134
rect 16606 27186 16658 27198
rect 41794 27134 41806 27186
rect 41858 27134 41870 27186
rect 43922 27134 43934 27186
rect 43986 27134 43998 27186
rect 16606 27122 16658 27134
rect 9886 27074 9938 27086
rect 9886 27010 9938 27022
rect 10446 27074 10498 27086
rect 17166 27074 17218 27086
rect 10882 27022 10894 27074
rect 10946 27022 10958 27074
rect 11554 27022 11566 27074
rect 11618 27022 11630 27074
rect 10446 27010 10498 27022
rect 17166 27010 17218 27022
rect 30830 27074 30882 27086
rect 30830 27010 30882 27022
rect 31614 27074 31666 27086
rect 31614 27010 31666 27022
rect 31950 27074 32002 27086
rect 31950 27010 32002 27022
rect 37886 27074 37938 27086
rect 41010 27022 41022 27074
rect 41074 27022 41086 27074
rect 37886 27010 37938 27022
rect 30718 26962 30770 26974
rect 30718 26898 30770 26910
rect 37550 26962 37602 26974
rect 37550 26898 37602 26910
rect 40686 26962 40738 26974
rect 40686 26898 40738 26910
rect 5854 26850 5906 26862
rect 5854 26786 5906 26798
rect 6078 26850 6130 26862
rect 6078 26786 6130 26798
rect 6302 26850 6354 26862
rect 6302 26786 6354 26798
rect 11118 26850 11170 26862
rect 11118 26786 11170 26798
rect 11342 26850 11394 26862
rect 11342 26786 11394 26798
rect 30494 26850 30546 26862
rect 30494 26786 30546 26798
rect 31838 26850 31890 26862
rect 31838 26786 31890 26798
rect 37774 26850 37826 26862
rect 37774 26786 37826 26798
rect 1344 26682 44576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 44576 26682
rect 1344 26596 44576 26630
rect 12238 26514 12290 26526
rect 4050 26462 4062 26514
rect 4114 26462 4126 26514
rect 12238 26450 12290 26462
rect 13022 26514 13074 26526
rect 13022 26450 13074 26462
rect 13134 26514 13186 26526
rect 33070 26514 33122 26526
rect 18722 26462 18734 26514
rect 18786 26462 18798 26514
rect 13134 26450 13186 26462
rect 33070 26450 33122 26462
rect 33294 26514 33346 26526
rect 33294 26450 33346 26462
rect 36990 26514 37042 26526
rect 36990 26450 37042 26462
rect 41694 26514 41746 26526
rect 41694 26450 41746 26462
rect 5294 26402 5346 26414
rect 5294 26338 5346 26350
rect 9886 26402 9938 26414
rect 9886 26338 9938 26350
rect 11118 26402 11170 26414
rect 15374 26402 15426 26414
rect 11890 26350 11902 26402
rect 11954 26350 11966 26402
rect 11118 26338 11170 26350
rect 15374 26338 15426 26350
rect 16606 26402 16658 26414
rect 33518 26402 33570 26414
rect 17714 26350 17726 26402
rect 17778 26350 17790 26402
rect 16606 26338 16658 26350
rect 33518 26338 33570 26350
rect 36654 26402 36706 26414
rect 36654 26338 36706 26350
rect 36766 26402 36818 26414
rect 36766 26338 36818 26350
rect 41806 26402 41858 26414
rect 42018 26350 42030 26402
rect 42082 26350 42094 26402
rect 41806 26338 41858 26350
rect 4510 26290 4562 26302
rect 4510 26226 4562 26238
rect 4622 26290 4674 26302
rect 5406 26290 5458 26302
rect 4834 26238 4846 26290
rect 4898 26238 4910 26290
rect 4622 26226 4674 26238
rect 5406 26226 5458 26238
rect 5518 26290 5570 26302
rect 10782 26290 10834 26302
rect 10546 26238 10558 26290
rect 10610 26238 10622 26290
rect 5518 26226 5570 26238
rect 10782 26226 10834 26238
rect 12910 26290 12962 26302
rect 12910 26226 12962 26238
rect 13582 26290 13634 26302
rect 13582 26226 13634 26238
rect 16270 26290 16322 26302
rect 16270 26226 16322 26238
rect 17390 26290 17442 26302
rect 17390 26226 17442 26238
rect 18398 26290 18450 26302
rect 41470 26290 41522 26302
rect 36194 26238 36206 26290
rect 36258 26238 36270 26290
rect 18398 26226 18450 26238
rect 41470 26226 41522 26238
rect 32510 26178 32562 26190
rect 9538 26126 9550 26178
rect 9602 26126 9614 26178
rect 15138 26126 15150 26178
rect 15202 26126 15214 26178
rect 32510 26114 32562 26126
rect 33182 26178 33234 26190
rect 33182 26114 33234 26126
rect 35870 26178 35922 26190
rect 41134 26178 41186 26190
rect 36642 26126 36654 26178
rect 36706 26126 36718 26178
rect 42242 26126 42254 26178
rect 42306 26126 42318 26178
rect 35870 26114 35922 26126
rect 41134 26114 41186 26126
rect 11006 26066 11058 26078
rect 5954 26014 5966 26066
rect 6018 26014 6030 26066
rect 11006 26002 11058 26014
rect 1344 25898 44576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 44576 25898
rect 1344 25812 44576 25846
rect 13570 25678 13582 25730
rect 13634 25678 13646 25730
rect 3614 25618 3666 25630
rect 3614 25554 3666 25566
rect 4734 25618 4786 25630
rect 22654 25618 22706 25630
rect 8306 25566 8318 25618
rect 8370 25566 8382 25618
rect 4734 25554 4786 25566
rect 22654 25554 22706 25566
rect 23102 25618 23154 25630
rect 35982 25618 36034 25630
rect 25218 25566 25230 25618
rect 25282 25566 25294 25618
rect 30482 25566 30494 25618
rect 30546 25566 30558 25618
rect 23102 25554 23154 25566
rect 35982 25554 36034 25566
rect 36430 25618 36482 25630
rect 39218 25566 39230 25618
rect 39282 25566 39294 25618
rect 36430 25554 36482 25566
rect 4398 25506 4450 25518
rect 5966 25506 6018 25518
rect 4834 25454 4846 25506
rect 4898 25454 4910 25506
rect 4398 25442 4450 25454
rect 5966 25442 6018 25454
rect 6190 25506 6242 25518
rect 6190 25442 6242 25454
rect 7198 25506 7250 25518
rect 11342 25506 11394 25518
rect 16046 25506 16098 25518
rect 23774 25506 23826 25518
rect 36990 25506 37042 25518
rect 7970 25454 7982 25506
rect 8034 25454 8046 25506
rect 8194 25454 8206 25506
rect 8258 25454 8270 25506
rect 14130 25454 14142 25506
rect 14194 25454 14206 25506
rect 14354 25454 14366 25506
rect 14418 25454 14430 25506
rect 14578 25454 14590 25506
rect 14642 25454 14654 25506
rect 21634 25454 21646 25506
rect 21698 25454 21710 25506
rect 24210 25454 24222 25506
rect 24274 25454 24286 25506
rect 24882 25454 24894 25506
rect 24946 25454 24958 25506
rect 30594 25454 30606 25506
rect 30658 25454 30670 25506
rect 30818 25454 30830 25506
rect 30882 25454 30894 25506
rect 38994 25454 39006 25506
rect 39058 25454 39070 25506
rect 40898 25454 40910 25506
rect 40962 25454 40974 25506
rect 7198 25442 7250 25454
rect 11342 25442 11394 25454
rect 16046 25442 16098 25454
rect 23774 25442 23826 25454
rect 36990 25442 37042 25454
rect 3838 25394 3890 25406
rect 3838 25330 3890 25342
rect 4622 25394 4674 25406
rect 4622 25330 4674 25342
rect 5742 25394 5794 25406
rect 5742 25330 5794 25342
rect 10782 25394 10834 25406
rect 10782 25330 10834 25342
rect 11006 25394 11058 25406
rect 21310 25394 21362 25406
rect 15698 25342 15710 25394
rect 15762 25342 15774 25394
rect 11006 25330 11058 25342
rect 21310 25330 21362 25342
rect 21422 25394 21474 25406
rect 39902 25394 39954 25406
rect 26002 25342 26014 25394
rect 26066 25342 26078 25394
rect 37314 25342 37326 25394
rect 37378 25342 37390 25394
rect 21422 25330 21474 25342
rect 39902 25330 39954 25342
rect 3726 25282 3778 25294
rect 3726 25218 3778 25230
rect 4062 25282 4114 25294
rect 4062 25218 4114 25230
rect 5070 25282 5122 25294
rect 5070 25218 5122 25230
rect 6078 25282 6130 25294
rect 6078 25218 6130 25230
rect 10670 25282 10722 25294
rect 10670 25218 10722 25230
rect 18062 25282 18114 25294
rect 24446 25282 24498 25294
rect 23426 25230 23438 25282
rect 23490 25230 23502 25282
rect 18062 25218 18114 25230
rect 24446 25218 24498 25230
rect 25678 25282 25730 25294
rect 25678 25218 25730 25230
rect 31054 25282 31106 25294
rect 31054 25218 31106 25230
rect 31278 25282 31330 25294
rect 31278 25218 31330 25230
rect 36318 25282 36370 25294
rect 41122 25230 41134 25282
rect 41186 25230 41198 25282
rect 36318 25218 36370 25230
rect 1344 25114 44576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 44576 25114
rect 1344 25028 44576 25062
rect 4734 24946 4786 24958
rect 4734 24882 4786 24894
rect 5070 24946 5122 24958
rect 5070 24882 5122 24894
rect 5854 24946 5906 24958
rect 5854 24882 5906 24894
rect 7870 24946 7922 24958
rect 7870 24882 7922 24894
rect 8766 24946 8818 24958
rect 8766 24882 8818 24894
rect 11118 24946 11170 24958
rect 11118 24882 11170 24894
rect 15934 24946 15986 24958
rect 15934 24882 15986 24894
rect 16382 24946 16434 24958
rect 16382 24882 16434 24894
rect 25342 24946 25394 24958
rect 25342 24882 25394 24894
rect 26238 24946 26290 24958
rect 26238 24882 26290 24894
rect 27134 24946 27186 24958
rect 27134 24882 27186 24894
rect 41022 24946 41074 24958
rect 41022 24882 41074 24894
rect 4622 24834 4674 24846
rect 4622 24770 4674 24782
rect 5294 24834 5346 24846
rect 5294 24770 5346 24782
rect 7646 24834 7698 24846
rect 7646 24770 7698 24782
rect 10110 24834 10162 24846
rect 10110 24770 10162 24782
rect 10558 24834 10610 24846
rect 10558 24770 10610 24782
rect 23886 24834 23938 24846
rect 23886 24770 23938 24782
rect 31950 24834 32002 24846
rect 40910 24834 40962 24846
rect 36194 24782 36206 24834
rect 36258 24782 36270 24834
rect 31950 24770 32002 24782
rect 40910 24770 40962 24782
rect 5406 24722 5458 24734
rect 5406 24658 5458 24670
rect 8094 24722 8146 24734
rect 8094 24658 8146 24670
rect 8318 24722 8370 24734
rect 8318 24658 8370 24670
rect 16158 24722 16210 24734
rect 16158 24658 16210 24670
rect 16606 24722 16658 24734
rect 16606 24658 16658 24670
rect 16830 24722 16882 24734
rect 25902 24722 25954 24734
rect 17378 24670 17390 24722
rect 17442 24670 17454 24722
rect 24210 24670 24222 24722
rect 24274 24670 24286 24722
rect 16830 24658 16882 24670
rect 25902 24658 25954 24670
rect 31278 24722 31330 24734
rect 31278 24658 31330 24670
rect 31614 24722 31666 24734
rect 38782 24722 38834 24734
rect 35522 24670 35534 24722
rect 35586 24670 35598 24722
rect 31614 24658 31666 24670
rect 38782 24658 38834 24670
rect 41246 24722 41298 24734
rect 41246 24658 41298 24670
rect 17950 24610 18002 24622
rect 17950 24546 18002 24558
rect 23998 24610 24050 24622
rect 23998 24546 24050 24558
rect 24670 24610 24722 24622
rect 31502 24610 31554 24622
rect 26674 24558 26686 24610
rect 26738 24558 26750 24610
rect 27570 24558 27582 24610
rect 27634 24558 27646 24610
rect 38322 24558 38334 24610
rect 38386 24558 38398 24610
rect 24670 24546 24722 24558
rect 31502 24546 31554 24558
rect 4846 24498 4898 24510
rect 4846 24434 4898 24446
rect 7758 24498 7810 24510
rect 7758 24434 7810 24446
rect 10222 24498 10274 24510
rect 10222 24434 10274 24446
rect 10670 24498 10722 24510
rect 10670 24434 10722 24446
rect 17726 24498 17778 24510
rect 17726 24434 17778 24446
rect 1344 24330 44576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 44576 24330
rect 1344 24244 44576 24278
rect 7198 24162 7250 24174
rect 21522 24110 21534 24162
rect 21586 24110 21598 24162
rect 7198 24098 7250 24110
rect 7758 24050 7810 24062
rect 7758 23986 7810 23998
rect 17950 24050 18002 24062
rect 17950 23986 18002 23998
rect 20862 24050 20914 24062
rect 40910 24050 40962 24062
rect 29922 23998 29934 24050
rect 29986 23998 29998 24050
rect 32050 23998 32062 24050
rect 32114 23998 32126 24050
rect 32386 23998 32398 24050
rect 32450 23998 32462 24050
rect 34514 23998 34526 24050
rect 34578 23998 34590 24050
rect 20862 23986 20914 23998
rect 40910 23986 40962 23998
rect 6190 23938 6242 23950
rect 6190 23874 6242 23886
rect 6750 23938 6802 23950
rect 22094 23938 22146 23950
rect 18274 23886 18286 23938
rect 18338 23886 18350 23938
rect 18498 23886 18510 23938
rect 18562 23886 18574 23938
rect 19618 23886 19630 23938
rect 19682 23886 19694 23938
rect 21522 23886 21534 23938
rect 21586 23886 21598 23938
rect 6750 23874 6802 23886
rect 22094 23874 22146 23886
rect 22430 23938 22482 23950
rect 22430 23874 22482 23886
rect 22542 23938 22594 23950
rect 22542 23874 22594 23886
rect 23102 23938 23154 23950
rect 23102 23874 23154 23886
rect 25454 23938 25506 23950
rect 25454 23874 25506 23886
rect 26014 23938 26066 23950
rect 35870 23938 35922 23950
rect 29250 23886 29262 23938
rect 29314 23886 29326 23938
rect 35298 23886 35310 23938
rect 35362 23886 35374 23938
rect 26014 23874 26066 23886
rect 35870 23874 35922 23886
rect 41246 23938 41298 23950
rect 41246 23874 41298 23886
rect 6526 23826 6578 23838
rect 6526 23762 6578 23774
rect 7086 23826 7138 23838
rect 7086 23762 7138 23774
rect 7198 23826 7250 23838
rect 22654 23826 22706 23838
rect 18722 23774 18734 23826
rect 18786 23774 18798 23826
rect 21858 23774 21870 23826
rect 21922 23774 21934 23826
rect 7198 23762 7250 23774
rect 22654 23762 22706 23774
rect 41470 23826 41522 23838
rect 41470 23762 41522 23774
rect 41582 23826 41634 23838
rect 41682 23774 41694 23826
rect 41746 23774 41758 23826
rect 41582 23762 41634 23774
rect 6302 23714 6354 23726
rect 6302 23650 6354 23662
rect 19966 23714 20018 23726
rect 19966 23650 20018 23662
rect 21982 23714 22034 23726
rect 21982 23650 22034 23662
rect 41358 23714 41410 23726
rect 41358 23650 41410 23662
rect 1344 23546 44576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 44576 23546
rect 1344 23460 44576 23494
rect 4958 23378 5010 23390
rect 4958 23314 5010 23326
rect 31166 23378 31218 23390
rect 31166 23314 31218 23326
rect 32398 23378 32450 23390
rect 34626 23326 34638 23378
rect 34690 23326 34702 23378
rect 32398 23314 32450 23326
rect 31278 23266 31330 23278
rect 14354 23214 14366 23266
rect 14418 23214 14430 23266
rect 15250 23214 15262 23266
rect 15314 23214 15326 23266
rect 20178 23214 20190 23266
rect 20242 23214 20254 23266
rect 31278 23202 31330 23214
rect 41806 23266 41858 23278
rect 41806 23202 41858 23214
rect 5294 23154 5346 23166
rect 14466 23102 14478 23154
rect 14530 23102 14542 23154
rect 14914 23102 14926 23154
rect 14978 23102 14990 23154
rect 18610 23102 18622 23154
rect 18674 23102 18686 23154
rect 19506 23102 19518 23154
rect 19570 23102 19582 23154
rect 34850 23102 34862 23154
rect 34914 23102 34926 23154
rect 5294 23090 5346 23102
rect 21198 23042 21250 23054
rect 18498 22990 18510 23042
rect 18562 22990 18574 23042
rect 21198 22978 21250 22990
rect 35422 23042 35474 23054
rect 35422 22978 35474 22990
rect 16046 22930 16098 22942
rect 41694 22930 41746 22942
rect 17826 22878 17838 22930
rect 17890 22878 17902 22930
rect 16046 22866 16098 22878
rect 41694 22866 41746 22878
rect 1344 22762 44576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 44576 22762
rect 1344 22676 44576 22710
rect 16830 22594 16882 22606
rect 16830 22530 16882 22542
rect 16270 22482 16322 22494
rect 2594 22430 2606 22482
rect 2658 22430 2670 22482
rect 4722 22430 4734 22482
rect 4786 22430 4798 22482
rect 9986 22430 9998 22482
rect 10050 22430 10062 22482
rect 16270 22418 16322 22430
rect 16494 22482 16546 22494
rect 16494 22418 16546 22430
rect 17166 22482 17218 22494
rect 41570 22430 41582 22482
rect 41634 22430 41646 22482
rect 43698 22430 43710 22482
rect 43762 22430 43774 22482
rect 17166 22418 17218 22430
rect 17726 22370 17778 22382
rect 1922 22318 1934 22370
rect 1986 22318 1998 22370
rect 7074 22318 7086 22370
rect 7138 22318 7150 22370
rect 8642 22318 8654 22370
rect 8706 22318 8718 22370
rect 17726 22306 17778 22318
rect 21534 22370 21586 22382
rect 21746 22318 21758 22370
rect 21810 22318 21822 22370
rect 40898 22318 40910 22370
rect 40962 22318 40974 22370
rect 21534 22306 21586 22318
rect 5742 22258 5794 22270
rect 7858 22206 7870 22258
rect 7922 22206 7934 22258
rect 8754 22206 8766 22258
rect 8818 22206 8830 22258
rect 26786 22206 26798 22258
rect 26850 22206 26862 22258
rect 5742 22194 5794 22206
rect 40462 22146 40514 22158
rect 40462 22082 40514 22094
rect 1344 21978 44576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 44576 21978
rect 1344 21892 44576 21926
rect 7534 21810 7586 21822
rect 15822 21810 15874 21822
rect 11442 21758 11454 21810
rect 11506 21758 11518 21810
rect 7534 21746 7586 21758
rect 15822 21746 15874 21758
rect 11566 21698 11618 21710
rect 10434 21646 10446 21698
rect 10498 21646 10510 21698
rect 12674 21646 12686 21698
rect 12738 21646 12750 21698
rect 13682 21646 13694 21698
rect 13746 21646 13758 21698
rect 22194 21646 22206 21698
rect 22258 21646 22270 21698
rect 11566 21634 11618 21646
rect 7422 21586 7474 21598
rect 16494 21586 16546 21598
rect 6402 21534 6414 21586
rect 6466 21534 6478 21586
rect 10770 21534 10782 21586
rect 10834 21534 10846 21586
rect 11778 21534 11790 21586
rect 11842 21534 11854 21586
rect 12114 21534 12126 21586
rect 12178 21534 12190 21586
rect 13794 21534 13806 21586
rect 13858 21534 13870 21586
rect 22978 21534 22990 21586
rect 23042 21534 23054 21586
rect 36082 21534 36094 21586
rect 36146 21534 36158 21586
rect 7422 21522 7474 21534
rect 16494 21522 16546 21534
rect 23550 21474 23602 21486
rect 39454 21474 39506 21486
rect 6514 21422 6526 21474
rect 6578 21422 6590 21474
rect 15362 21422 15374 21474
rect 15426 21422 15438 21474
rect 20066 21422 20078 21474
rect 20130 21422 20142 21474
rect 36866 21422 36878 21474
rect 36930 21422 36942 21474
rect 38994 21422 39006 21474
rect 39058 21422 39070 21474
rect 23550 21410 23602 21422
rect 39454 21410 39506 21422
rect 16270 21362 16322 21374
rect 16270 21298 16322 21310
rect 16606 21362 16658 21374
rect 16606 21298 16658 21310
rect 1344 21194 44576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 44576 21194
rect 1344 21108 44576 21142
rect 34626 20974 34638 21026
rect 34690 20974 34702 21026
rect 37326 20914 37378 20926
rect 8306 20862 8318 20914
rect 8370 20862 8382 20914
rect 13794 20862 13806 20914
rect 13858 20862 13870 20914
rect 37326 20850 37378 20862
rect 8194 20750 8206 20802
rect 8258 20750 8270 20802
rect 9090 20750 9102 20802
rect 9154 20750 9166 20802
rect 9986 20750 9998 20802
rect 10050 20750 10062 20802
rect 10546 20750 10558 20802
rect 10610 20750 10622 20802
rect 11442 20750 11454 20802
rect 11506 20750 11518 20802
rect 12674 20750 12686 20802
rect 12738 20750 12750 20802
rect 13458 20750 13470 20802
rect 13522 20750 13534 20802
rect 14914 20750 14926 20802
rect 14978 20750 14990 20802
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 17378 20750 17390 20802
rect 17442 20750 17454 20802
rect 37538 20750 37550 20802
rect 37602 20750 37614 20802
rect 17950 20690 18002 20702
rect 7746 20638 7758 20690
rect 7810 20638 7822 20690
rect 9874 20638 9886 20690
rect 9938 20638 9950 20690
rect 11330 20638 11342 20690
rect 11394 20638 11406 20690
rect 13906 20638 13918 20690
rect 13970 20638 13982 20690
rect 15362 20638 15374 20690
rect 15426 20638 15438 20690
rect 17950 20626 18002 20638
rect 34974 20690 35026 20702
rect 34974 20626 35026 20638
rect 35198 20690 35250 20702
rect 35198 20626 35250 20638
rect 35422 20690 35474 20702
rect 35422 20626 35474 20638
rect 37214 20690 37266 20702
rect 37214 20626 37266 20638
rect 10670 20578 10722 20590
rect 14702 20578 14754 20590
rect 8978 20526 8990 20578
rect 9042 20526 9054 20578
rect 10546 20526 10558 20578
rect 10610 20526 10622 20578
rect 12338 20526 12350 20578
rect 12402 20526 12414 20578
rect 12562 20526 12574 20578
rect 12626 20526 12638 20578
rect 16930 20526 16942 20578
rect 16994 20526 17006 20578
rect 10670 20514 10722 20526
rect 14702 20514 14754 20526
rect 1344 20410 44576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 44576 20410
rect 1344 20324 44576 20358
rect 5394 20190 5406 20242
rect 5458 20190 5470 20242
rect 34962 20190 34974 20242
rect 35026 20190 35038 20242
rect 5966 20130 6018 20142
rect 3154 20078 3166 20130
rect 3218 20078 3230 20130
rect 5966 20066 6018 20078
rect 7758 20130 7810 20142
rect 7758 20066 7810 20078
rect 16718 20130 16770 20142
rect 16718 20066 16770 20078
rect 22654 20130 22706 20142
rect 35410 20078 35422 20130
rect 35474 20078 35486 20130
rect 35634 20078 35646 20130
rect 35698 20078 35710 20130
rect 22654 20066 22706 20078
rect 2370 19966 2382 20018
rect 2434 19966 2446 20018
rect 7074 19966 7086 20018
rect 7138 19966 7150 20018
rect 7522 19966 7534 20018
rect 7586 19966 7598 20018
rect 12114 19966 12126 20018
rect 12178 19966 12190 20018
rect 12898 19966 12910 20018
rect 12962 19966 12974 20018
rect 13794 19966 13806 20018
rect 13858 19966 13870 20018
rect 14242 19966 14254 20018
rect 14306 19966 14318 20018
rect 22866 19966 22878 20018
rect 22930 19966 22942 20018
rect 25778 19966 25790 20018
rect 25842 19966 25854 20018
rect 29922 19966 29934 20018
rect 29986 19966 29998 20018
rect 31378 19966 31390 20018
rect 31442 19966 31454 20018
rect 35970 19966 35982 20018
rect 36034 19966 36046 20018
rect 9998 19906 10050 19918
rect 16158 19906 16210 19918
rect 31950 19906 32002 19918
rect 11778 19854 11790 19906
rect 11842 19854 11854 19906
rect 15250 19854 15262 19906
rect 15314 19854 15326 19906
rect 26562 19854 26574 19906
rect 26626 19854 26638 19906
rect 28690 19854 28702 19906
rect 28754 19854 28766 19906
rect 30034 19854 30046 19906
rect 30098 19854 30110 19906
rect 9998 19842 10050 19854
rect 16158 19842 16210 19854
rect 31950 19842 32002 19854
rect 10110 19794 10162 19806
rect 10110 19730 10162 19742
rect 22878 19794 22930 19806
rect 22878 19730 22930 19742
rect 23214 19794 23266 19806
rect 31726 19794 31778 19806
rect 29250 19742 29262 19794
rect 29314 19742 29326 19794
rect 23214 19730 23266 19742
rect 31726 19730 31778 19742
rect 1344 19626 44576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 44576 19626
rect 1344 19540 44576 19574
rect 26686 19458 26738 19470
rect 26686 19394 26738 19406
rect 38894 19458 38946 19470
rect 38894 19394 38946 19406
rect 26574 19346 26626 19358
rect 23650 19294 23662 19346
rect 23714 19294 23726 19346
rect 25778 19294 25790 19346
rect 25842 19294 25854 19346
rect 26574 19282 26626 19294
rect 27134 19346 27186 19358
rect 27134 19282 27186 19294
rect 29262 19346 29314 19358
rect 29262 19282 29314 19294
rect 30046 19346 30098 19358
rect 37550 19346 37602 19358
rect 35410 19294 35422 19346
rect 35474 19294 35486 19346
rect 30046 19282 30098 19294
rect 37550 19282 37602 19294
rect 9102 19234 9154 19246
rect 16270 19234 16322 19246
rect 30718 19234 30770 19246
rect 8306 19182 8318 19234
rect 8370 19182 8382 19234
rect 9426 19182 9438 19234
rect 9490 19182 9502 19234
rect 11666 19182 11678 19234
rect 11730 19182 11742 19234
rect 22978 19182 22990 19234
rect 23042 19182 23054 19234
rect 26338 19182 26350 19234
rect 26402 19182 26414 19234
rect 30370 19182 30382 19234
rect 30434 19182 30446 19234
rect 9102 19170 9154 19182
rect 16270 19170 16322 19182
rect 30718 19170 30770 19182
rect 31502 19234 31554 19246
rect 38334 19234 38386 19246
rect 32050 19182 32062 19234
rect 32114 19182 32126 19234
rect 34066 19182 34078 19234
rect 34130 19182 34142 19234
rect 37986 19182 37998 19234
rect 38050 19182 38062 19234
rect 31502 19170 31554 19182
rect 38334 19170 38386 19182
rect 38670 19234 38722 19246
rect 38670 19170 38722 19182
rect 34638 19122 34690 19134
rect 10882 19070 10894 19122
rect 10946 19070 10958 19122
rect 16482 19070 16494 19122
rect 16546 19070 16558 19122
rect 17266 19070 17278 19122
rect 17330 19070 17342 19122
rect 32162 19070 32174 19122
rect 32226 19070 32238 19122
rect 34638 19058 34690 19070
rect 11902 19010 11954 19022
rect 30606 19010 30658 19022
rect 16594 18958 16606 19010
rect 16658 18958 16670 19010
rect 11902 18946 11954 18958
rect 30606 18946 30658 18958
rect 31166 19010 31218 19022
rect 31166 18946 31218 18958
rect 31390 19010 31442 19022
rect 31390 18946 31442 18958
rect 31614 19010 31666 19022
rect 39218 18958 39230 19010
rect 39282 18958 39294 19010
rect 31614 18946 31666 18958
rect 1344 18842 44576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 44576 18842
rect 1344 18756 44576 18790
rect 16158 18562 16210 18574
rect 16482 18510 16494 18562
rect 16546 18510 16558 18562
rect 31602 18510 31614 18562
rect 31666 18510 31678 18562
rect 16158 18498 16210 18510
rect 15374 18450 15426 18462
rect 22094 18450 22146 18462
rect 39118 18450 39170 18462
rect 14914 18398 14926 18450
rect 14978 18398 14990 18450
rect 21634 18398 21646 18450
rect 21698 18398 21710 18450
rect 32386 18398 32398 18450
rect 32450 18398 32462 18450
rect 35746 18398 35758 18450
rect 35810 18398 35822 18450
rect 41794 18398 41806 18450
rect 41858 18398 41870 18450
rect 15374 18386 15426 18398
rect 22094 18386 22146 18398
rect 39118 18386 39170 18398
rect 26014 18338 26066 18350
rect 33182 18338 33234 18350
rect 10098 18286 10110 18338
rect 10162 18286 10174 18338
rect 18722 18286 18734 18338
rect 18786 18286 18798 18338
rect 20850 18286 20862 18338
rect 20914 18286 20926 18338
rect 29474 18286 29486 18338
rect 29538 18286 29550 18338
rect 36530 18286 36542 18338
rect 36594 18286 36606 18338
rect 38658 18286 38670 18338
rect 38722 18286 38734 18338
rect 41682 18286 41694 18338
rect 41746 18286 41758 18338
rect 26014 18274 26066 18286
rect 33182 18274 33234 18286
rect 41470 18226 41522 18238
rect 41470 18162 41522 18174
rect 1344 18058 44576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 44576 18058
rect 1344 17972 44576 18006
rect 8878 17890 8930 17902
rect 8878 17826 8930 17838
rect 12350 17890 12402 17902
rect 12350 17826 12402 17838
rect 36990 17890 37042 17902
rect 36990 17826 37042 17838
rect 37326 17890 37378 17902
rect 37326 17826 37378 17838
rect 10558 17778 10610 17790
rect 10558 17714 10610 17726
rect 12238 17778 12290 17790
rect 12238 17714 12290 17726
rect 19518 17778 19570 17790
rect 19518 17714 19570 17726
rect 20190 17778 20242 17790
rect 20190 17714 20242 17726
rect 39566 17778 39618 17790
rect 39566 17714 39618 17726
rect 40014 17778 40066 17790
rect 41682 17726 41694 17778
rect 41746 17726 41758 17778
rect 43810 17726 43822 17778
rect 43874 17726 43886 17778
rect 40014 17714 40066 17726
rect 9886 17666 9938 17678
rect 9650 17614 9662 17666
rect 9714 17614 9726 17666
rect 9886 17602 9938 17614
rect 10110 17666 10162 17678
rect 10110 17602 10162 17614
rect 16158 17666 16210 17678
rect 37102 17666 37154 17678
rect 40686 17666 40738 17678
rect 19730 17614 19742 17666
rect 19794 17614 19806 17666
rect 37538 17614 37550 17666
rect 37602 17614 37614 17666
rect 40898 17614 40910 17666
rect 40962 17614 40974 17666
rect 16158 17602 16210 17614
rect 37102 17602 37154 17614
rect 40686 17602 40738 17614
rect 8990 17554 9042 17566
rect 8990 17490 9042 17502
rect 9998 17554 10050 17566
rect 9998 17490 10050 17502
rect 10670 17554 10722 17566
rect 10670 17490 10722 17502
rect 19406 17554 19458 17566
rect 19406 17490 19458 17502
rect 40350 17554 40402 17566
rect 40350 17490 40402 17502
rect 40462 17554 40514 17566
rect 40462 17490 40514 17502
rect 9214 17442 9266 17454
rect 17054 17442 17106 17454
rect 15810 17390 15822 17442
rect 15874 17390 15886 17442
rect 9214 17378 9266 17390
rect 17054 17378 17106 17390
rect 36430 17442 36482 17454
rect 36430 17378 36482 17390
rect 1344 17274 44576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 44576 17274
rect 1344 17188 44576 17222
rect 6974 17106 7026 17118
rect 10334 17106 10386 17118
rect 9874 17054 9886 17106
rect 9938 17054 9950 17106
rect 6974 17042 7026 17054
rect 10334 17042 10386 17054
rect 11118 17106 11170 17118
rect 11118 17042 11170 17054
rect 13134 17106 13186 17118
rect 13134 17042 13186 17054
rect 40238 17106 40290 17118
rect 40238 17042 40290 17054
rect 41470 17106 41522 17118
rect 41470 17042 41522 17054
rect 11902 16994 11954 17006
rect 4386 16942 4398 16994
rect 4450 16942 4462 16994
rect 11902 16930 11954 16942
rect 13806 16994 13858 17006
rect 13806 16930 13858 16942
rect 14030 16994 14082 17006
rect 14030 16930 14082 16942
rect 14142 16994 14194 17006
rect 14142 16930 14194 16942
rect 17390 16994 17442 17006
rect 17390 16930 17442 16942
rect 40126 16994 40178 17006
rect 40126 16930 40178 16942
rect 41246 16994 41298 17006
rect 41246 16930 41298 16942
rect 9550 16882 9602 16894
rect 3602 16830 3614 16882
rect 3666 16830 3678 16882
rect 9550 16818 9602 16830
rect 10222 16882 10274 16894
rect 11566 16882 11618 16894
rect 13694 16882 13746 16894
rect 11106 16830 11118 16882
rect 11170 16830 11182 16882
rect 13346 16830 13358 16882
rect 13410 16830 13422 16882
rect 10222 16818 10274 16830
rect 11566 16818 11618 16830
rect 13694 16818 13746 16830
rect 15710 16882 15762 16894
rect 17950 16882 18002 16894
rect 16146 16830 16158 16882
rect 16210 16830 16222 16882
rect 15710 16818 15762 16830
rect 17950 16818 18002 16830
rect 33182 16882 33234 16894
rect 40462 16882 40514 16894
rect 33506 16830 33518 16882
rect 33570 16830 33582 16882
rect 33182 16818 33234 16830
rect 40462 16818 40514 16830
rect 16606 16770 16658 16782
rect 6514 16718 6526 16770
rect 6578 16718 6590 16770
rect 38098 16718 38110 16770
rect 38162 16718 38174 16770
rect 41570 16718 41582 16770
rect 41634 16718 41646 16770
rect 16606 16706 16658 16718
rect 11454 16658 11506 16670
rect 11454 16594 11506 16606
rect 13022 16658 13074 16670
rect 13022 16594 13074 16606
rect 1344 16490 44576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 44576 16490
rect 1344 16404 44576 16438
rect 9538 16270 9550 16322
rect 9602 16270 9614 16322
rect 5742 16210 5794 16222
rect 2594 16158 2606 16210
rect 2658 16158 2670 16210
rect 4722 16158 4734 16210
rect 4786 16158 4798 16210
rect 5742 16146 5794 16158
rect 9102 16210 9154 16222
rect 9102 16146 9154 16158
rect 12350 16210 12402 16222
rect 12350 16146 12402 16158
rect 19294 16210 19346 16222
rect 19294 16146 19346 16158
rect 23214 16210 23266 16222
rect 23214 16146 23266 16158
rect 24222 16210 24274 16222
rect 31938 16158 31950 16210
rect 32002 16158 32014 16210
rect 24222 16146 24274 16158
rect 8990 16098 9042 16110
rect 12126 16098 12178 16110
rect 1922 16046 1934 16098
rect 1986 16046 1998 16098
rect 9762 16046 9774 16098
rect 9826 16046 9838 16098
rect 8990 16034 9042 16046
rect 12126 16034 12178 16046
rect 12462 16098 12514 16110
rect 25006 16098 25058 16110
rect 12674 16046 12686 16098
rect 12738 16046 12750 16098
rect 17266 16046 17278 16098
rect 17330 16046 17342 16098
rect 29362 16046 29374 16098
rect 29426 16046 29438 16098
rect 12462 16034 12514 16046
rect 25006 16034 25058 16046
rect 12238 15986 12290 15998
rect 23326 15986 23378 15998
rect 9202 15934 9214 15986
rect 9266 15934 9278 15986
rect 15810 15934 15822 15986
rect 15874 15934 15886 15986
rect 12238 15922 12290 15934
rect 23326 15922 23378 15934
rect 23550 15986 23602 15998
rect 23550 15922 23602 15934
rect 24558 15986 24610 15998
rect 24558 15922 24610 15934
rect 24670 15986 24722 15998
rect 24670 15922 24722 15934
rect 24894 15986 24946 15998
rect 24894 15922 24946 15934
rect 25454 15986 25506 15998
rect 25454 15922 25506 15934
rect 25678 15986 25730 15998
rect 25678 15922 25730 15934
rect 26350 15986 26402 15998
rect 26350 15922 26402 15934
rect 22990 15874 23042 15886
rect 22990 15810 23042 15822
rect 23102 15874 23154 15886
rect 23102 15810 23154 15822
rect 25342 15874 25394 15886
rect 25342 15810 25394 15822
rect 26014 15874 26066 15886
rect 26014 15810 26066 15822
rect 28702 15874 28754 15886
rect 28702 15810 28754 15822
rect 1344 15706 44576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 44576 15706
rect 1344 15620 44576 15654
rect 9886 15538 9938 15550
rect 9886 15474 9938 15486
rect 9998 15538 10050 15550
rect 9998 15474 10050 15486
rect 12910 15538 12962 15550
rect 12910 15474 12962 15486
rect 17726 15538 17778 15550
rect 17726 15474 17778 15486
rect 17838 15538 17890 15550
rect 23102 15538 23154 15550
rect 19506 15486 19518 15538
rect 19570 15486 19582 15538
rect 20850 15486 20862 15538
rect 20914 15486 20926 15538
rect 22418 15486 22430 15538
rect 22482 15486 22494 15538
rect 17838 15474 17890 15486
rect 23102 15474 23154 15486
rect 24446 15538 24498 15550
rect 24446 15474 24498 15486
rect 24558 15538 24610 15550
rect 24558 15474 24610 15486
rect 29262 15538 29314 15550
rect 29262 15474 29314 15486
rect 33406 15538 33458 15550
rect 33406 15474 33458 15486
rect 9774 15426 9826 15438
rect 9774 15362 9826 15374
rect 17390 15426 17442 15438
rect 17390 15362 17442 15374
rect 18846 15426 18898 15438
rect 18846 15362 18898 15374
rect 19966 15426 20018 15438
rect 19966 15362 20018 15374
rect 21870 15426 21922 15438
rect 28018 15374 28030 15426
rect 28082 15374 28094 15426
rect 33058 15374 33070 15426
rect 33122 15374 33134 15426
rect 21870 15362 21922 15374
rect 10110 15314 10162 15326
rect 9538 15262 9550 15314
rect 9602 15262 9614 15314
rect 10110 15250 10162 15262
rect 17614 15314 17666 15326
rect 19182 15314 19234 15326
rect 22094 15314 22146 15326
rect 18050 15262 18062 15314
rect 18114 15262 18126 15314
rect 18610 15262 18622 15314
rect 18674 15262 18686 15314
rect 21074 15262 21086 15314
rect 21138 15262 21150 15314
rect 17614 15250 17666 15262
rect 19182 15250 19234 15262
rect 22094 15250 22146 15262
rect 22766 15314 22818 15326
rect 22766 15250 22818 15262
rect 23102 15314 23154 15326
rect 23102 15250 23154 15262
rect 23326 15314 23378 15326
rect 23326 15250 23378 15262
rect 23886 15314 23938 15326
rect 24210 15262 24222 15314
rect 24274 15262 24286 15314
rect 28802 15262 28814 15314
rect 28866 15262 28878 15314
rect 29586 15262 29598 15314
rect 29650 15262 29662 15314
rect 34850 15262 34862 15314
rect 34914 15262 34926 15314
rect 23886 15250 23938 15262
rect 38110 15202 38162 15214
rect 20402 15150 20414 15202
rect 20466 15150 20478 15202
rect 25890 15150 25902 15202
rect 25954 15150 25966 15202
rect 30370 15150 30382 15202
rect 30434 15150 30446 15202
rect 32498 15150 32510 15202
rect 32562 15150 32574 15202
rect 35522 15150 35534 15202
rect 35586 15150 35598 15202
rect 37650 15150 37662 15202
rect 37714 15150 37726 15202
rect 38110 15138 38162 15150
rect 1344 14922 44576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 44576 14922
rect 1344 14836 44576 14870
rect 16270 14754 16322 14766
rect 16270 14690 16322 14702
rect 23550 14754 23602 14766
rect 23550 14690 23602 14702
rect 23886 14754 23938 14766
rect 23886 14690 23938 14702
rect 11006 14642 11058 14654
rect 11006 14578 11058 14590
rect 16494 14642 16546 14654
rect 16494 14578 16546 14590
rect 17054 14642 17106 14654
rect 17054 14578 17106 14590
rect 18062 14642 18114 14654
rect 18062 14578 18114 14590
rect 18846 14642 18898 14654
rect 18846 14578 18898 14590
rect 19294 14642 19346 14654
rect 19294 14578 19346 14590
rect 31502 14642 31554 14654
rect 31502 14578 31554 14590
rect 32734 14642 32786 14654
rect 32734 14578 32786 14590
rect 11342 14530 11394 14542
rect 11342 14466 11394 14478
rect 14926 14530 14978 14542
rect 17726 14530 17778 14542
rect 15474 14478 15486 14530
rect 15538 14478 15550 14530
rect 15922 14478 15934 14530
rect 15986 14478 15998 14530
rect 14926 14466 14978 14478
rect 17726 14466 17778 14478
rect 18174 14530 18226 14542
rect 31726 14530 31778 14542
rect 23874 14478 23886 14530
rect 23938 14478 23950 14530
rect 18174 14466 18226 14478
rect 31726 14466 31778 14478
rect 36430 14530 36482 14542
rect 41246 14530 41298 14542
rect 37538 14478 37550 14530
rect 37602 14478 37614 14530
rect 36430 14466 36482 14478
rect 41246 14466 41298 14478
rect 8654 14418 8706 14430
rect 8654 14354 8706 14366
rect 11678 14418 11730 14430
rect 31390 14418 31442 14430
rect 14578 14366 14590 14418
rect 14642 14366 14654 14418
rect 11678 14354 11730 14366
rect 31390 14354 31442 14366
rect 31950 14418 32002 14430
rect 37650 14366 37662 14418
rect 37714 14366 37726 14418
rect 41346 14366 41358 14418
rect 41410 14366 41422 14418
rect 31950 14354 32002 14366
rect 8766 14306 8818 14318
rect 36094 14306 36146 14318
rect 15250 14254 15262 14306
rect 15314 14254 15326 14306
rect 17378 14254 17390 14306
rect 17442 14254 17454 14306
rect 38994 14254 39006 14306
rect 39058 14254 39070 14306
rect 8766 14242 8818 14254
rect 36094 14242 36146 14254
rect 1344 14138 44576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 44576 14138
rect 1344 14052 44576 14086
rect 14814 13970 14866 13982
rect 14814 13906 14866 13918
rect 15598 13970 15650 13982
rect 15598 13906 15650 13918
rect 16718 13970 16770 13982
rect 31950 13970 32002 13982
rect 27234 13918 27246 13970
rect 27298 13918 27310 13970
rect 16718 13906 16770 13918
rect 31950 13906 32002 13918
rect 36094 13970 36146 13982
rect 36094 13906 36146 13918
rect 39902 13970 39954 13982
rect 39902 13906 39954 13918
rect 8542 13858 8594 13870
rect 8542 13794 8594 13806
rect 9550 13858 9602 13870
rect 9550 13794 9602 13806
rect 21534 13858 21586 13870
rect 21534 13794 21586 13806
rect 21646 13858 21698 13870
rect 21646 13794 21698 13806
rect 23998 13858 24050 13870
rect 23998 13794 24050 13806
rect 24110 13858 24162 13870
rect 28814 13858 28866 13870
rect 26338 13806 26350 13858
rect 26402 13806 26414 13858
rect 24110 13794 24162 13806
rect 28814 13794 28866 13806
rect 37438 13858 37490 13870
rect 37438 13794 37490 13806
rect 8654 13746 8706 13758
rect 24222 13746 24274 13758
rect 28366 13746 28418 13758
rect 9762 13694 9774 13746
rect 9826 13694 9838 13746
rect 10210 13694 10222 13746
rect 10274 13694 10286 13746
rect 26226 13694 26238 13746
rect 26290 13694 26302 13746
rect 8654 13682 8706 13694
rect 24222 13682 24274 13694
rect 28366 13682 28418 13694
rect 31614 13746 31666 13758
rect 31614 13682 31666 13694
rect 31838 13746 31890 13758
rect 31838 13682 31890 13694
rect 32062 13746 32114 13758
rect 35758 13746 35810 13758
rect 32386 13694 32398 13746
rect 32450 13694 32462 13746
rect 32062 13682 32114 13694
rect 35758 13682 35810 13694
rect 35870 13746 35922 13758
rect 35870 13682 35922 13694
rect 36206 13746 36258 13758
rect 36206 13682 36258 13694
rect 36542 13746 36594 13758
rect 36542 13682 36594 13694
rect 36766 13746 36818 13758
rect 36766 13682 36818 13694
rect 37214 13746 37266 13758
rect 37214 13682 37266 13694
rect 37326 13746 37378 13758
rect 41010 13694 41022 13746
rect 41074 13694 41086 13746
rect 37326 13682 37378 13694
rect 9662 13634 9714 13646
rect 40350 13634 40402 13646
rect 15138 13582 15150 13634
rect 15202 13582 15214 13634
rect 41794 13582 41806 13634
rect 41858 13582 41870 13634
rect 43922 13582 43934 13634
rect 43986 13582 43998 13634
rect 9662 13570 9714 13582
rect 40350 13570 40402 13582
rect 8542 13522 8594 13534
rect 8542 13458 8594 13470
rect 9998 13522 10050 13534
rect 9998 13458 10050 13470
rect 21646 13522 21698 13534
rect 40238 13522 40290 13534
rect 24658 13470 24670 13522
rect 24722 13470 24734 13522
rect 31378 13470 31390 13522
rect 31442 13519 31454 13522
rect 31602 13519 31614 13522
rect 31442 13473 31614 13519
rect 31442 13470 31454 13473
rect 31602 13470 31614 13473
rect 31666 13470 31678 13522
rect 21646 13458 21698 13470
rect 40238 13458 40290 13470
rect 1344 13354 44576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 44576 13354
rect 1344 13268 44576 13302
rect 10434 13134 10446 13186
rect 10498 13134 10510 13186
rect 9202 13022 9214 13074
rect 9266 13022 9278 13074
rect 11106 13022 11118 13074
rect 11170 13022 11182 13074
rect 40114 13022 40126 13074
rect 40178 13022 40190 13074
rect 10222 12962 10274 12974
rect 21870 12962 21922 12974
rect 7970 12910 7982 12962
rect 8034 12910 8046 12962
rect 8642 12910 8654 12962
rect 8706 12910 8718 12962
rect 10434 12910 10446 12962
rect 10498 12910 10510 12962
rect 10222 12898 10274 12910
rect 21870 12898 21922 12910
rect 22094 12962 22146 12974
rect 22094 12898 22146 12910
rect 40798 12962 40850 12974
rect 40798 12898 40850 12910
rect 41022 12962 41074 12974
rect 41022 12898 41074 12910
rect 8878 12850 8930 12862
rect 8878 12786 8930 12798
rect 9886 12850 9938 12862
rect 9886 12786 9938 12798
rect 11454 12850 11506 12862
rect 11454 12786 11506 12798
rect 11678 12850 11730 12862
rect 11678 12786 11730 12798
rect 21646 12850 21698 12862
rect 40238 12850 40290 12862
rect 23202 12798 23214 12850
rect 23266 12798 23278 12850
rect 21646 12786 21698 12798
rect 40238 12786 40290 12798
rect 40462 12850 40514 12862
rect 41694 12850 41746 12862
rect 41346 12798 41358 12850
rect 41410 12798 41422 12850
rect 40462 12786 40514 12798
rect 41694 12786 41746 12798
rect 42030 12850 42082 12862
rect 42030 12786 42082 12798
rect 8094 12738 8146 12750
rect 8094 12674 8146 12686
rect 9102 12738 9154 12750
rect 9102 12674 9154 12686
rect 9214 12738 9266 12750
rect 11118 12738 11170 12750
rect 10210 12686 10222 12738
rect 10274 12686 10286 12738
rect 9214 12674 9266 12686
rect 11118 12674 11170 12686
rect 11230 12738 11282 12750
rect 11230 12674 11282 12686
rect 21982 12738 22034 12750
rect 21982 12674 22034 12686
rect 22878 12738 22930 12750
rect 22878 12674 22930 12686
rect 1344 12570 44576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 44576 12570
rect 1344 12484 44576 12518
rect 13134 12402 13186 12414
rect 37662 12402 37714 12414
rect 6402 12350 6414 12402
rect 6466 12350 6478 12402
rect 22754 12350 22766 12402
rect 22818 12350 22830 12402
rect 13134 12338 13186 12350
rect 37662 12338 37714 12350
rect 38446 12402 38498 12414
rect 38446 12338 38498 12350
rect 40798 12402 40850 12414
rect 40798 12338 40850 12350
rect 41022 12402 41074 12414
rect 41022 12338 41074 12350
rect 8878 12290 8930 12302
rect 21534 12290 21586 12302
rect 4162 12238 4174 12290
rect 4226 12238 4238 12290
rect 10098 12238 10110 12290
rect 10162 12238 10174 12290
rect 11106 12238 11118 12290
rect 11170 12238 11182 12290
rect 21298 12238 21310 12290
rect 21362 12238 21374 12290
rect 8878 12226 8930 12238
rect 21534 12226 21586 12238
rect 21646 12290 21698 12302
rect 21646 12226 21698 12238
rect 21758 12290 21810 12302
rect 38098 12238 38110 12290
rect 38162 12238 38174 12290
rect 21758 12226 21810 12238
rect 21870 12178 21922 12190
rect 3490 12126 3502 12178
rect 3554 12126 3566 12178
rect 8530 12126 8542 12178
rect 8594 12126 8606 12178
rect 9538 12126 9550 12178
rect 9602 12126 9614 12178
rect 11218 12126 11230 12178
rect 11282 12126 11294 12178
rect 21870 12114 21922 12126
rect 22206 12178 22258 12190
rect 41134 12178 41186 12190
rect 37426 12126 37438 12178
rect 37490 12126 37502 12178
rect 22206 12114 22258 12126
rect 41134 12114 41186 12126
rect 6974 12066 7026 12078
rect 6974 12002 7026 12014
rect 8766 12066 8818 12078
rect 13694 12066 13746 12078
rect 12898 12014 12910 12066
rect 12962 12014 12974 12066
rect 8766 12002 8818 12014
rect 13694 12002 13746 12014
rect 37102 12066 37154 12078
rect 37102 12002 37154 12014
rect 22430 11954 22482 11966
rect 22430 11890 22482 11902
rect 37774 11954 37826 11966
rect 37774 11890 37826 11902
rect 1344 11786 44576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 44576 11786
rect 1344 11700 44576 11734
rect 25566 11618 25618 11630
rect 12786 11566 12798 11618
rect 12850 11615 12862 11618
rect 13010 11615 13022 11618
rect 12850 11569 13022 11615
rect 12850 11566 12862 11569
rect 13010 11566 13022 11569
rect 13074 11566 13086 11618
rect 25566 11554 25618 11566
rect 5742 11506 5794 11518
rect 22206 11506 22258 11518
rect 4834 11454 4846 11506
rect 4898 11454 4910 11506
rect 21298 11454 21310 11506
rect 21362 11454 21374 11506
rect 5742 11442 5794 11454
rect 22206 11442 22258 11454
rect 24558 11506 24610 11518
rect 24558 11442 24610 11454
rect 8766 11394 8818 11406
rect 1922 11342 1934 11394
rect 1986 11342 1998 11394
rect 2594 11342 2606 11394
rect 2658 11342 2670 11394
rect 8766 11330 8818 11342
rect 9102 11394 9154 11406
rect 9102 11330 9154 11342
rect 17166 11394 17218 11406
rect 25454 11394 25506 11406
rect 17714 11342 17726 11394
rect 17778 11342 17790 11394
rect 17166 11330 17218 11342
rect 25454 11330 25506 11342
rect 31614 11394 31666 11406
rect 31614 11330 31666 11342
rect 31838 11394 31890 11406
rect 31838 11330 31890 11342
rect 32734 11394 32786 11406
rect 35870 11394 35922 11406
rect 32946 11342 32958 11394
rect 33010 11342 33022 11394
rect 32734 11330 32786 11342
rect 35870 11330 35922 11342
rect 36206 11394 36258 11406
rect 36206 11330 36258 11342
rect 36430 11394 36482 11406
rect 36430 11330 36482 11342
rect 37438 11394 37490 11406
rect 37438 11330 37490 11342
rect 37550 11394 37602 11406
rect 37550 11330 37602 11342
rect 37662 11394 37714 11406
rect 37662 11330 37714 11342
rect 21422 11282 21474 11294
rect 12114 11230 12126 11282
rect 12178 11230 12190 11282
rect 21422 11218 21474 11230
rect 21646 11282 21698 11294
rect 21646 11218 21698 11230
rect 25118 11282 25170 11294
rect 25118 11218 25170 11230
rect 26014 11282 26066 11294
rect 26014 11218 26066 11230
rect 26350 11282 26402 11294
rect 26350 11218 26402 11230
rect 31278 11282 31330 11294
rect 31278 11218 31330 11230
rect 32622 11282 32674 11294
rect 32622 11218 32674 11230
rect 8878 11170 8930 11182
rect 8878 11106 8930 11118
rect 11790 11170 11842 11182
rect 11790 11106 11842 11118
rect 17278 11170 17330 11182
rect 17278 11106 17330 11118
rect 17390 11170 17442 11182
rect 17390 11106 17442 11118
rect 17502 11170 17554 11182
rect 17502 11106 17554 11118
rect 24782 11170 24834 11182
rect 24782 11106 24834 11118
rect 25006 11170 25058 11182
rect 25006 11106 25058 11118
rect 25566 11170 25618 11182
rect 25566 11106 25618 11118
rect 26126 11170 26178 11182
rect 26126 11106 26178 11118
rect 31502 11170 31554 11182
rect 34526 11170 34578 11182
rect 32162 11118 32174 11170
rect 32226 11118 32238 11170
rect 34178 11118 34190 11170
rect 34242 11118 34254 11170
rect 31502 11106 31554 11118
rect 34526 11106 34578 11118
rect 35982 11170 36034 11182
rect 36978 11118 36990 11170
rect 37042 11118 37054 11170
rect 35982 11106 36034 11118
rect 1344 11002 44576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 44576 11002
rect 1344 10916 44576 10950
rect 8430 10834 8482 10846
rect 8430 10770 8482 10782
rect 9886 10834 9938 10846
rect 9886 10770 9938 10782
rect 9998 10834 10050 10846
rect 9998 10770 10050 10782
rect 10670 10834 10722 10846
rect 10670 10770 10722 10782
rect 12462 10834 12514 10846
rect 12462 10770 12514 10782
rect 13022 10834 13074 10846
rect 13022 10770 13074 10782
rect 16270 10834 16322 10846
rect 16270 10770 16322 10782
rect 17614 10834 17666 10846
rect 17614 10770 17666 10782
rect 24446 10834 24498 10846
rect 24446 10770 24498 10782
rect 24670 10834 24722 10846
rect 24670 10770 24722 10782
rect 25566 10834 25618 10846
rect 25566 10770 25618 10782
rect 25790 10834 25842 10846
rect 25790 10770 25842 10782
rect 26686 10834 26738 10846
rect 26686 10770 26738 10782
rect 33182 10834 33234 10846
rect 33182 10770 33234 10782
rect 35086 10834 35138 10846
rect 35086 10770 35138 10782
rect 35870 10834 35922 10846
rect 35870 10770 35922 10782
rect 9550 10722 9602 10734
rect 9550 10658 9602 10670
rect 12574 10722 12626 10734
rect 12574 10658 12626 10670
rect 13582 10722 13634 10734
rect 20862 10722 20914 10734
rect 18386 10670 18398 10722
rect 18450 10670 18462 10722
rect 13582 10658 13634 10670
rect 20862 10658 20914 10670
rect 24222 10722 24274 10734
rect 24222 10658 24274 10670
rect 25342 10722 25394 10734
rect 25342 10658 25394 10670
rect 27022 10722 27074 10734
rect 27022 10658 27074 10670
rect 8206 10610 8258 10622
rect 7858 10558 7870 10610
rect 7922 10558 7934 10610
rect 8206 10546 8258 10558
rect 9774 10610 9826 10622
rect 12238 10610 12290 10622
rect 35534 10610 35586 10622
rect 10210 10558 10222 10610
rect 10274 10558 10286 10610
rect 13906 10558 13918 10610
rect 13970 10558 13982 10610
rect 18274 10558 18286 10610
rect 18338 10558 18350 10610
rect 20290 10558 20302 10610
rect 20354 10558 20366 10610
rect 29698 10558 29710 10610
rect 29762 10558 29774 10610
rect 9774 10546 9826 10558
rect 12238 10546 12290 10558
rect 35534 10546 35586 10558
rect 35758 10610 35810 10622
rect 35970 10558 35982 10610
rect 36034 10558 36046 10610
rect 35758 10546 35810 10558
rect 8318 10498 8370 10510
rect 8318 10434 8370 10446
rect 8878 10498 8930 10510
rect 8878 10434 8930 10446
rect 15262 10498 15314 10510
rect 25454 10498 25506 10510
rect 21634 10446 21646 10498
rect 21698 10446 21710 10498
rect 24658 10446 24670 10498
rect 24722 10446 24734 10498
rect 30370 10446 30382 10498
rect 30434 10446 30446 10498
rect 32498 10446 32510 10498
rect 32562 10446 32574 10498
rect 15262 10434 15314 10446
rect 25454 10434 25506 10446
rect 13918 10386 13970 10398
rect 8642 10334 8654 10386
rect 8706 10383 8718 10386
rect 9090 10383 9102 10386
rect 8706 10337 9102 10383
rect 8706 10334 8718 10337
rect 9090 10334 9102 10337
rect 9154 10334 9166 10386
rect 17266 10334 17278 10386
rect 17330 10383 17342 10386
rect 18050 10383 18062 10386
rect 17330 10337 18062 10383
rect 17330 10334 17342 10337
rect 18050 10334 18062 10337
rect 18114 10334 18126 10386
rect 13918 10322 13970 10334
rect 1344 10218 44576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 44576 10218
rect 1344 10132 44576 10166
rect 8430 10050 8482 10062
rect 17838 10050 17890 10062
rect 20414 10050 20466 10062
rect 17154 9998 17166 10050
rect 17218 9998 17230 10050
rect 19842 9998 19854 10050
rect 19906 9998 19918 10050
rect 8430 9986 8482 9998
rect 17838 9986 17890 9998
rect 20414 9986 20466 9998
rect 31278 10050 31330 10062
rect 31278 9986 31330 9998
rect 31614 10050 31666 10062
rect 31614 9986 31666 9998
rect 8094 9938 8146 9950
rect 8094 9874 8146 9886
rect 12686 9938 12738 9950
rect 12686 9874 12738 9886
rect 24894 9938 24946 9950
rect 29262 9938 29314 9950
rect 26450 9886 26462 9938
rect 26514 9886 26526 9938
rect 28578 9886 28590 9938
rect 28642 9886 28654 9938
rect 24894 9874 24946 9886
rect 29262 9874 29314 9886
rect 7534 9826 7586 9838
rect 12462 9826 12514 9838
rect 12226 9774 12238 9826
rect 12290 9774 12302 9826
rect 7534 9762 7586 9774
rect 12462 9762 12514 9774
rect 12910 9826 12962 9838
rect 12910 9762 12962 9774
rect 14366 9826 14418 9838
rect 14366 9762 14418 9774
rect 15038 9826 15090 9838
rect 15038 9762 15090 9774
rect 15486 9826 15538 9838
rect 15486 9762 15538 9774
rect 15598 9826 15650 9838
rect 15598 9762 15650 9774
rect 16606 9826 16658 9838
rect 16606 9762 16658 9774
rect 16942 9826 16994 9838
rect 17614 9826 17666 9838
rect 17378 9774 17390 9826
rect 17442 9774 17454 9826
rect 16942 9762 16994 9774
rect 17614 9762 17666 9774
rect 19070 9826 19122 9838
rect 19070 9762 19122 9774
rect 19294 9826 19346 9838
rect 19294 9762 19346 9774
rect 19630 9826 19682 9838
rect 24782 9826 24834 9838
rect 19842 9774 19854 9826
rect 19906 9774 19918 9826
rect 19630 9762 19682 9774
rect 24782 9762 24834 9774
rect 25118 9826 25170 9838
rect 25118 9762 25170 9774
rect 25342 9826 25394 9838
rect 31390 9826 31442 9838
rect 25778 9774 25790 9826
rect 25842 9774 25854 9826
rect 31826 9774 31838 9826
rect 31890 9774 31902 9826
rect 25342 9762 25394 9774
rect 31390 9762 31442 9774
rect 8654 9714 8706 9726
rect 8654 9650 8706 9662
rect 12014 9714 12066 9726
rect 12014 9650 12066 9662
rect 16046 9714 16098 9726
rect 16046 9650 16098 9662
rect 20526 9714 20578 9726
rect 20526 9650 20578 9662
rect 8542 9602 8594 9614
rect 13582 9602 13634 9614
rect 12338 9550 12350 9602
rect 12402 9550 12414 9602
rect 8542 9538 8594 9550
rect 13582 9538 13634 9550
rect 14814 9602 14866 9614
rect 14814 9538 14866 9550
rect 14926 9602 14978 9614
rect 14926 9538 14978 9550
rect 15710 9602 15762 9614
rect 15710 9538 15762 9550
rect 15822 9602 15874 9614
rect 17950 9602 18002 9614
rect 16818 9550 16830 9602
rect 16882 9550 16894 9602
rect 15822 9538 15874 9550
rect 17950 9538 18002 9550
rect 18174 9602 18226 9614
rect 30942 9602 30994 9614
rect 19618 9550 19630 9602
rect 19682 9550 19694 9602
rect 18174 9538 18226 9550
rect 30942 9538 30994 9550
rect 1344 9434 44576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 44576 9434
rect 1344 9348 44576 9382
rect 12238 9266 12290 9278
rect 12238 9202 12290 9214
rect 12350 9266 12402 9278
rect 17390 9266 17442 9278
rect 12350 9202 12402 9214
rect 16494 9210 16546 9222
rect 14814 9154 14866 9166
rect 14814 9090 14866 9102
rect 15598 9154 15650 9166
rect 15598 9090 15650 9102
rect 15710 9154 15762 9166
rect 17390 9202 17442 9214
rect 18174 9266 18226 9278
rect 18174 9202 18226 9214
rect 20190 9266 20242 9278
rect 20190 9202 20242 9214
rect 21086 9266 21138 9278
rect 21086 9202 21138 9214
rect 23998 9266 24050 9278
rect 23998 9202 24050 9214
rect 16494 9146 16546 9158
rect 17950 9154 18002 9166
rect 15710 9090 15762 9102
rect 17950 9090 18002 9102
rect 20078 9154 20130 9166
rect 20078 9090 20130 9102
rect 24334 9154 24386 9166
rect 24334 9090 24386 9102
rect 24558 9154 24610 9166
rect 24558 9090 24610 9102
rect 26126 9154 26178 9166
rect 26126 9090 26178 9102
rect 26462 9154 26514 9166
rect 26462 9090 26514 9102
rect 26574 9154 26626 9166
rect 35746 9102 35758 9154
rect 35810 9102 35822 9154
rect 26574 9090 26626 9102
rect 12126 9042 12178 9054
rect 12126 8978 12178 8990
rect 12798 9042 12850 9054
rect 17838 9042 17890 9054
rect 15138 8990 15150 9042
rect 15202 8990 15214 9042
rect 16706 8990 16718 9042
rect 16770 8990 16782 9042
rect 12798 8978 12850 8990
rect 17838 8978 17890 8990
rect 20414 9042 20466 9054
rect 20414 8978 20466 8990
rect 20638 9042 20690 9054
rect 20638 8978 20690 8990
rect 25118 9042 25170 9054
rect 25678 9042 25730 9054
rect 25442 8990 25454 9042
rect 25506 8990 25518 9042
rect 25118 8978 25170 8990
rect 25678 8978 25730 8990
rect 25902 9042 25954 9054
rect 38334 9042 38386 9054
rect 35074 8990 35086 9042
rect 35138 8990 35150 9042
rect 25902 8978 25954 8990
rect 38334 8978 38386 8990
rect 14926 8930 14978 8942
rect 14926 8866 14978 8878
rect 17502 8930 17554 8942
rect 26014 8930 26066 8942
rect 24658 8878 24670 8930
rect 24722 8878 24734 8930
rect 37874 8878 37886 8930
rect 37938 8878 37950 8930
rect 17502 8866 17554 8878
rect 26014 8866 26066 8878
rect 15710 8818 15762 8830
rect 15710 8754 15762 8766
rect 1344 8650 44576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 44576 8650
rect 1344 8564 44576 8598
rect 9102 8370 9154 8382
rect 5618 8318 5630 8370
rect 5682 8318 5694 8370
rect 7746 8318 7758 8370
rect 7810 8318 7822 8370
rect 9102 8306 9154 8318
rect 25006 8370 25058 8382
rect 25006 8306 25058 8318
rect 8530 8206 8542 8258
rect 8594 8206 8606 8258
rect 1344 7866 44576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 44576 7866
rect 1344 7780 44576 7814
rect 1344 7082 44576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 44576 7082
rect 1344 6996 44576 7030
rect 9650 6750 9662 6802
rect 9714 6750 9726 6802
rect 21646 6690 21698 6702
rect 11778 6638 11790 6690
rect 11842 6638 11854 6690
rect 12562 6638 12574 6690
rect 12626 6638 12638 6690
rect 21646 6626 21698 6638
rect 18062 6578 18114 6590
rect 18062 6514 18114 6526
rect 18398 6578 18450 6590
rect 18398 6514 18450 6526
rect 13582 6466 13634 6478
rect 13582 6402 13634 6414
rect 21758 6466 21810 6478
rect 21758 6402 21810 6414
rect 1344 6298 44576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 44576 6298
rect 1344 6212 44576 6246
rect 28590 6130 28642 6142
rect 18610 6078 18622 6130
rect 18674 6078 18686 6130
rect 28590 6066 28642 6078
rect 19070 6018 19122 6030
rect 19070 5954 19122 5966
rect 21086 6018 21138 6030
rect 26002 5966 26014 6018
rect 26066 5966 26078 6018
rect 21086 5954 21138 5966
rect 22206 5906 22258 5918
rect 18498 5854 18510 5906
rect 18562 5854 18574 5906
rect 25330 5854 25342 5906
rect 25394 5854 25406 5906
rect 22206 5842 22258 5854
rect 28130 5742 28142 5794
rect 28194 5742 28206 5794
rect 1344 5514 44576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 44576 5514
rect 1344 5428 44576 5462
rect 24782 5234 24834 5246
rect 16482 5182 16494 5234
rect 16546 5182 16558 5234
rect 18610 5182 18622 5234
rect 18674 5182 18686 5234
rect 21298 5182 21310 5234
rect 21362 5182 21374 5234
rect 23426 5182 23438 5234
rect 23490 5182 23502 5234
rect 24782 5170 24834 5182
rect 15374 5122 15426 5134
rect 15810 5070 15822 5122
rect 15874 5070 15886 5122
rect 24098 5070 24110 5122
rect 24162 5070 24174 5122
rect 15374 5058 15426 5070
rect 1344 4730 44576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 44576 4730
rect 1344 4644 44576 4678
rect 16830 4562 16882 4574
rect 16830 4498 16882 4510
rect 18734 4562 18786 4574
rect 18734 4498 18786 4510
rect 14242 4398 14254 4450
rect 14306 4398 14318 4450
rect 19842 4398 19854 4450
rect 19906 4398 19918 4450
rect 13570 4286 13582 4338
rect 13634 4286 13646 4338
rect 19170 4286 19182 4338
rect 19234 4286 19246 4338
rect 16370 4174 16382 4226
rect 16434 4174 16446 4226
rect 21970 4174 21982 4226
rect 22034 4174 22046 4226
rect 1344 3946 44576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 44576 3946
rect 1344 3860 44576 3894
rect 1344 3162 44576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 44576 3162
rect 1344 3076 44576 3110
<< via1 >>
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 18286 42142 18338 42194
rect 33518 42142 33570 42194
rect 6190 42030 6242 42082
rect 9998 42030 10050 42082
rect 5070 41918 5122 41970
rect 5854 41918 5906 41970
rect 8878 41918 8930 41970
rect 9662 41918 9714 41970
rect 13470 41918 13522 41970
rect 17278 41918 17330 41970
rect 21086 41918 21138 41970
rect 24894 41918 24946 41970
rect 28702 41918 28754 41970
rect 32510 41918 32562 41970
rect 36318 41918 36370 41970
rect 40126 41918 40178 41970
rect 14478 41806 14530 41858
rect 22094 41806 22146 41858
rect 25902 41806 25954 41858
rect 29710 41806 29762 41858
rect 37326 41806 37378 41858
rect 41134 41806 41186 41858
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 43598 41246 43650 41298
rect 41582 41134 41634 41186
rect 13918 40910 13970 40962
rect 28478 40910 28530 40962
rect 39790 40910 39842 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 6302 40574 6354 40626
rect 10446 40574 10498 40626
rect 32622 40574 32674 40626
rect 10222 40462 10274 40514
rect 34190 40462 34242 40514
rect 3054 40350 3106 40402
rect 10110 40350 10162 40402
rect 10782 40350 10834 40402
rect 14030 40350 14082 40402
rect 17614 40350 17666 40402
rect 20078 40350 20130 40402
rect 20302 40350 20354 40402
rect 25342 40350 25394 40402
rect 28478 40350 28530 40402
rect 29262 40350 29314 40402
rect 31838 40350 31890 40402
rect 33406 40350 33458 40402
rect 36878 40350 36930 40402
rect 3726 40238 3778 40290
rect 5854 40238 5906 40290
rect 11454 40238 11506 40290
rect 13582 40238 13634 40290
rect 14702 40238 14754 40290
rect 16830 40238 16882 40290
rect 21086 40238 21138 40290
rect 23214 40238 23266 40290
rect 26014 40238 26066 40290
rect 28142 40238 28194 40290
rect 31390 40238 31442 40290
rect 36318 40238 36370 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 9102 39790 9154 39842
rect 6414 39678 6466 39730
rect 11342 39678 11394 39730
rect 17054 39678 17106 39730
rect 20302 39678 20354 39730
rect 34414 39678 34466 39730
rect 34974 39678 35026 39730
rect 37998 39678 38050 39730
rect 38334 39678 38386 39730
rect 6974 39566 7026 39618
rect 7758 39566 7810 39618
rect 7982 39566 8034 39618
rect 9214 39566 9266 39618
rect 9662 39566 9714 39618
rect 10222 39566 10274 39618
rect 10782 39566 10834 39618
rect 11230 39566 11282 39618
rect 11790 39566 11842 39618
rect 17502 39566 17554 39618
rect 31502 39566 31554 39618
rect 41134 39566 41186 39618
rect 41470 39566 41522 39618
rect 41806 39566 41858 39618
rect 7646 39454 7698 39506
rect 9774 39454 9826 39506
rect 11902 39454 11954 39506
rect 13918 39454 13970 39506
rect 14254 39454 14306 39506
rect 18174 39454 18226 39506
rect 32174 39454 32226 39506
rect 40462 39454 40514 39506
rect 41694 39454 41746 39506
rect 42142 39454 42194 39506
rect 6302 39342 6354 39394
rect 6526 39342 6578 39394
rect 7310 39342 7362 39394
rect 7534 39342 7586 39394
rect 8318 39342 8370 39394
rect 8542 39342 8594 39394
rect 8654 39342 8706 39394
rect 9102 39342 9154 39394
rect 9886 39342 9938 39394
rect 11454 39342 11506 39394
rect 12126 39342 12178 39394
rect 28254 39342 28306 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 5182 39006 5234 39058
rect 7982 39006 8034 39058
rect 9550 39006 9602 39058
rect 12126 39006 12178 39058
rect 39230 39006 39282 39058
rect 40350 39006 40402 39058
rect 2606 38894 2658 38946
rect 7646 38894 7698 38946
rect 7758 38894 7810 38946
rect 8878 38894 8930 38946
rect 10782 38894 10834 38946
rect 11566 38894 11618 38946
rect 40126 38894 40178 38946
rect 1934 38782 1986 38834
rect 8990 38782 9042 38834
rect 9886 38782 9938 38834
rect 10222 38782 10274 38834
rect 11790 38782 11842 38834
rect 40014 38782 40066 38834
rect 41134 38782 41186 38834
rect 4734 38670 4786 38722
rect 39678 38670 39730 38722
rect 41918 38670 41970 38722
rect 44046 38670 44098 38722
rect 10446 38558 10498 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 37886 38222 37938 38274
rect 10110 38110 10162 38162
rect 38334 38110 38386 38162
rect 42030 38110 42082 38162
rect 9662 37998 9714 38050
rect 10222 37998 10274 38050
rect 10558 37998 10610 38050
rect 25566 37998 25618 38050
rect 25790 37998 25842 38050
rect 38110 37998 38162 38050
rect 40798 37998 40850 38050
rect 41022 37998 41074 38050
rect 41358 37998 41410 38050
rect 41806 37998 41858 38050
rect 11454 37886 11506 37938
rect 24894 37886 24946 37938
rect 40462 37886 40514 37938
rect 41582 37886 41634 37938
rect 42142 37886 42194 37938
rect 42366 37886 42418 37938
rect 42702 37886 42754 37938
rect 43150 37886 43202 37938
rect 12126 37774 12178 37826
rect 26350 37774 26402 37826
rect 39790 37774 39842 37826
rect 40238 37774 40290 37826
rect 40574 37774 40626 37826
rect 41134 37774 41186 37826
rect 42590 37774 42642 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 6862 37438 6914 37490
rect 19742 37438 19794 37490
rect 25566 37326 25618 37378
rect 30830 37326 30882 37378
rect 7086 37214 7138 37266
rect 20078 37214 20130 37266
rect 24334 37214 24386 37266
rect 25230 37214 25282 37266
rect 27582 37214 27634 37266
rect 34638 37214 34690 37266
rect 37774 37214 37826 37266
rect 20862 37102 20914 37154
rect 22990 37102 23042 37154
rect 23662 37102 23714 37154
rect 24558 37102 24610 37154
rect 28254 37102 28306 37154
rect 30382 37102 30434 37154
rect 35310 37102 35362 37154
rect 37438 37102 37490 37154
rect 38222 37102 38274 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 21534 36654 21586 36706
rect 21870 36654 21922 36706
rect 24222 36654 24274 36706
rect 27918 36654 27970 36706
rect 27134 36542 27186 36594
rect 37662 36542 37714 36594
rect 17278 36430 17330 36482
rect 17502 36430 17554 36482
rect 24334 36430 24386 36482
rect 26798 36430 26850 36482
rect 29486 36430 29538 36482
rect 30830 36430 30882 36482
rect 31278 36430 31330 36482
rect 7086 36318 7138 36370
rect 15598 36318 15650 36370
rect 16942 36318 16994 36370
rect 18062 36318 18114 36370
rect 26910 36318 26962 36370
rect 27246 36318 27298 36370
rect 27582 36318 27634 36370
rect 27806 36318 27858 36370
rect 29150 36318 29202 36370
rect 30382 36318 30434 36370
rect 7198 36206 7250 36258
rect 10446 36206 10498 36258
rect 15486 36206 15538 36258
rect 17726 36206 17778 36258
rect 17950 36206 18002 36258
rect 20862 36206 20914 36258
rect 21646 36206 21698 36258
rect 24222 36206 24274 36258
rect 28366 36206 28418 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 10670 35870 10722 35922
rect 19070 35870 19122 35922
rect 41358 35870 41410 35922
rect 2606 35758 2658 35810
rect 7646 35758 7698 35810
rect 11118 35758 11170 35810
rect 11230 35758 11282 35810
rect 14702 35758 14754 35810
rect 17950 35758 18002 35810
rect 18622 35758 18674 35810
rect 19630 35758 19682 35810
rect 41806 35758 41858 35810
rect 41918 35758 41970 35810
rect 1934 35646 1986 35698
rect 7982 35646 8034 35698
rect 11342 35646 11394 35698
rect 14926 35646 14978 35698
rect 15262 35646 15314 35698
rect 15710 35646 15762 35698
rect 16382 35646 16434 35698
rect 17390 35646 17442 35698
rect 17838 35646 17890 35698
rect 18174 35646 18226 35698
rect 18734 35646 18786 35698
rect 19182 35646 19234 35698
rect 20078 35646 20130 35698
rect 20526 35646 20578 35698
rect 41582 35646 41634 35698
rect 4734 35534 4786 35586
rect 5182 35534 5234 35586
rect 10334 35534 10386 35586
rect 16270 35534 16322 35586
rect 9774 35422 9826 35474
rect 10110 35422 10162 35474
rect 14590 35422 14642 35474
rect 15934 35422 15986 35474
rect 16494 35422 16546 35474
rect 18622 35422 18674 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 17166 35086 17218 35138
rect 17726 35086 17778 35138
rect 18062 35086 18114 35138
rect 9886 34974 9938 35026
rect 10782 34974 10834 35026
rect 11342 34974 11394 35026
rect 15598 34974 15650 35026
rect 16830 34974 16882 35026
rect 33070 34974 33122 35026
rect 40574 34974 40626 35026
rect 43822 34974 43874 35026
rect 8766 34862 8818 34914
rect 9326 34862 9378 34914
rect 10222 34862 10274 34914
rect 11118 34862 11170 34914
rect 11566 34862 11618 34914
rect 11678 34862 11730 34914
rect 14702 34862 14754 34914
rect 15374 34862 15426 34914
rect 25566 34862 25618 34914
rect 30270 34862 30322 34914
rect 33518 34862 33570 34914
rect 41022 34862 41074 34914
rect 14366 34750 14418 34802
rect 14926 34750 14978 34802
rect 15934 34750 15986 34802
rect 17390 34750 17442 34802
rect 25790 34750 25842 34802
rect 30942 34750 30994 34802
rect 41694 34750 41746 34802
rect 9102 34638 9154 34690
rect 9774 34638 9826 34690
rect 9998 34638 10050 34690
rect 10670 34638 10722 34690
rect 10894 34638 10946 34690
rect 12350 34638 12402 34690
rect 14142 34638 14194 34690
rect 14478 34638 14530 34690
rect 15710 34638 15762 34690
rect 17838 34638 17890 34690
rect 25678 34638 25730 34690
rect 26014 34638 26066 34690
rect 27134 34638 27186 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 10110 34302 10162 34354
rect 14702 34302 14754 34354
rect 26574 34302 26626 34354
rect 26798 34302 26850 34354
rect 27358 34302 27410 34354
rect 27694 34302 27746 34354
rect 38894 34302 38946 34354
rect 4958 34190 5010 34242
rect 9662 34190 9714 34242
rect 27918 34190 27970 34242
rect 31838 34190 31890 34242
rect 4286 34078 4338 34130
rect 9550 34078 9602 34130
rect 10558 34078 10610 34130
rect 14142 34078 14194 34130
rect 26350 34078 26402 34130
rect 27134 34078 27186 34130
rect 27470 34078 27522 34130
rect 28030 34078 28082 34130
rect 32062 34078 32114 34130
rect 38334 34078 38386 34130
rect 42254 34078 42306 34130
rect 7086 33966 7138 34018
rect 7534 33966 7586 34018
rect 10894 33966 10946 34018
rect 11454 33966 11506 34018
rect 26686 33966 26738 34018
rect 35534 33966 35586 34018
rect 37662 33966 37714 34018
rect 41918 33966 41970 34018
rect 14366 33854 14418 33906
rect 41470 33854 41522 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 30830 33518 30882 33570
rect 10222 33406 10274 33458
rect 23102 33406 23154 33458
rect 25118 33406 25170 33458
rect 35870 33406 35922 33458
rect 37102 33406 37154 33458
rect 41806 33406 41858 33458
rect 11342 33294 11394 33346
rect 23774 33294 23826 33346
rect 27022 33294 27074 33346
rect 30942 33294 30994 33346
rect 31390 33294 31442 33346
rect 32958 33294 33010 33346
rect 36094 33294 36146 33346
rect 37326 33294 37378 33346
rect 37774 33294 37826 33346
rect 41694 33294 41746 33346
rect 42254 33294 42306 33346
rect 24670 33182 24722 33234
rect 26686 33182 26738 33234
rect 30718 33182 30770 33234
rect 31614 33182 31666 33234
rect 31726 33182 31778 33234
rect 32622 33182 32674 33234
rect 32734 33182 32786 33234
rect 35758 33182 35810 33234
rect 36318 33182 36370 33234
rect 36990 33182 37042 33234
rect 37550 33182 37602 33234
rect 38110 33182 38162 33234
rect 42030 33182 42082 33234
rect 11678 33070 11730 33122
rect 26798 33070 26850 33122
rect 27470 33070 27522 33122
rect 31166 33070 31218 33122
rect 34750 33070 34802 33122
rect 35086 33070 35138 33122
rect 35422 33070 35474 33122
rect 37998 33070 38050 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 19630 32734 19682 32786
rect 30830 32734 30882 32786
rect 31054 32734 31106 32786
rect 31502 32734 31554 32786
rect 32398 32734 32450 32786
rect 36878 32734 36930 32786
rect 37102 32734 37154 32786
rect 37214 32734 37266 32786
rect 42142 32734 42194 32786
rect 15486 32622 15538 32674
rect 37438 32622 37490 32674
rect 41918 32622 41970 32674
rect 15262 32510 15314 32562
rect 19966 32510 20018 32562
rect 23886 32510 23938 32562
rect 24110 32510 24162 32562
rect 26574 32510 26626 32562
rect 31166 32510 31218 32562
rect 31726 32510 31778 32562
rect 32062 32510 32114 32562
rect 32286 32510 32338 32562
rect 36766 32510 36818 32562
rect 37550 32510 37602 32562
rect 41806 32510 41858 32562
rect 20750 32398 20802 32450
rect 22878 32398 22930 32450
rect 23214 32398 23266 32450
rect 26126 32398 26178 32450
rect 27022 32398 27074 32450
rect 31838 32398 31890 32450
rect 32398 32286 32450 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 21534 31950 21586 32002
rect 21870 31950 21922 32002
rect 5070 31838 5122 31890
rect 25678 31838 25730 31890
rect 26238 31838 26290 31890
rect 27134 31838 27186 31890
rect 27582 31838 27634 31890
rect 2158 31726 2210 31778
rect 12910 31726 12962 31778
rect 13582 31726 13634 31778
rect 14030 31726 14082 31778
rect 19966 31726 20018 31778
rect 25790 31726 25842 31778
rect 26686 31726 26738 31778
rect 30046 31726 30098 31778
rect 2942 31614 2994 31666
rect 15150 31614 15202 31666
rect 25342 31614 25394 31666
rect 26126 31614 26178 31666
rect 26462 31614 26514 31666
rect 40350 31614 40402 31666
rect 5742 31502 5794 31554
rect 20750 31502 20802 31554
rect 21646 31502 21698 31554
rect 25566 31502 25618 31554
rect 30270 31502 30322 31554
rect 30718 31502 30770 31554
rect 36430 31502 36482 31554
rect 36990 31502 37042 31554
rect 37326 31502 37378 31554
rect 39678 31502 39730 31554
rect 40014 31502 40066 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4174 31166 4226 31218
rect 16270 31166 16322 31218
rect 31726 31166 31778 31218
rect 41470 31166 41522 31218
rect 30718 31054 30770 31106
rect 31502 31054 31554 31106
rect 36654 31054 36706 31106
rect 40014 31054 40066 31106
rect 40126 31054 40178 31106
rect 41806 31054 41858 31106
rect 6078 30942 6130 30994
rect 15934 30942 15986 30994
rect 16494 30942 16546 30994
rect 16830 30942 16882 30994
rect 17950 30942 18002 30994
rect 30606 30942 30658 30994
rect 30942 30942 30994 30994
rect 31390 30942 31442 30994
rect 32510 30942 32562 30994
rect 33406 30942 33458 30994
rect 40350 30942 40402 30994
rect 41134 30942 41186 30994
rect 41582 30942 41634 30994
rect 4286 30830 4338 30882
rect 6862 30830 6914 30882
rect 8990 30830 9042 30882
rect 9662 30830 9714 30882
rect 10894 30830 10946 30882
rect 16382 30830 16434 30882
rect 17502 30830 17554 30882
rect 20190 30830 20242 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 15822 30382 15874 30434
rect 9550 30270 9602 30322
rect 16158 30270 16210 30322
rect 41470 30270 41522 30322
rect 43598 30270 43650 30322
rect 12462 30158 12514 30210
rect 13022 30158 13074 30210
rect 14926 30158 14978 30210
rect 18958 30158 19010 30210
rect 19630 30158 19682 30210
rect 28590 30158 28642 30210
rect 30158 30158 30210 30210
rect 35310 30158 35362 30210
rect 37438 30158 37490 30210
rect 40686 30158 40738 30210
rect 11678 30046 11730 30098
rect 15710 30046 15762 30098
rect 18286 30046 18338 30098
rect 33518 30046 33570 30098
rect 34974 30046 35026 30098
rect 35982 30046 36034 30098
rect 36990 30046 37042 30098
rect 37326 30046 37378 30098
rect 39118 30046 39170 30098
rect 39342 30046 39394 30098
rect 39454 30046 39506 30098
rect 15150 29934 15202 29986
rect 15598 29934 15650 29986
rect 35198 29934 35250 29986
rect 35646 29934 35698 29986
rect 36430 29934 36482 29986
rect 37102 29934 37154 29986
rect 40350 29934 40402 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 5854 29598 5906 29650
rect 11230 29598 11282 29650
rect 11902 29598 11954 29650
rect 22990 29598 23042 29650
rect 24110 29598 24162 29650
rect 32062 29598 32114 29650
rect 38222 29598 38274 29650
rect 41470 29598 41522 29650
rect 23214 29486 23266 29538
rect 36990 29486 37042 29538
rect 41694 29486 41746 29538
rect 41806 29486 41858 29538
rect 1934 29374 1986 29426
rect 11454 29374 11506 29426
rect 14366 29374 14418 29426
rect 23438 29374 23490 29426
rect 28814 29374 28866 29426
rect 37774 29374 37826 29426
rect 2606 29262 2658 29314
rect 4846 29262 4898 29314
rect 5518 29262 5570 29314
rect 23998 29262 24050 29314
rect 29486 29262 29538 29314
rect 31614 29262 31666 29314
rect 34862 29262 34914 29314
rect 11118 29150 11170 29202
rect 13918 29150 13970 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 4510 28814 4562 28866
rect 15934 28814 15986 28866
rect 29262 28814 29314 28866
rect 29822 28814 29874 28866
rect 30382 28814 30434 28866
rect 5742 28702 5794 28754
rect 6974 28702 7026 28754
rect 15150 28702 15202 28754
rect 27022 28702 27074 28754
rect 6414 28590 6466 28642
rect 11566 28590 11618 28642
rect 11902 28590 11954 28642
rect 12350 28590 12402 28642
rect 12462 28590 12514 28642
rect 12686 28590 12738 28642
rect 12910 28590 12962 28642
rect 15710 28590 15762 28642
rect 16270 28590 16322 28642
rect 16494 28590 16546 28642
rect 16718 28590 16770 28642
rect 17278 28590 17330 28642
rect 21310 28590 21362 28642
rect 21534 28590 21586 28642
rect 21982 28590 22034 28642
rect 22318 28590 22370 28642
rect 26574 28590 26626 28642
rect 29598 28590 29650 28642
rect 30942 28590 30994 28642
rect 31950 28590 32002 28642
rect 32510 28590 32562 28642
rect 32846 28590 32898 28642
rect 34638 28590 34690 28642
rect 35982 28590 36034 28642
rect 5070 28478 5122 28530
rect 5854 28478 5906 28530
rect 5966 28478 6018 28530
rect 17390 28478 17442 28530
rect 26238 28478 26290 28530
rect 29374 28478 29426 28530
rect 29934 28478 29986 28530
rect 32286 28478 32338 28530
rect 32734 28478 32786 28530
rect 36318 28478 36370 28530
rect 4622 28366 4674 28418
rect 4846 28366 4898 28418
rect 5630 28366 5682 28418
rect 15150 28366 15202 28418
rect 15374 28366 15426 28418
rect 17166 28366 17218 28418
rect 21758 28366 21810 28418
rect 28590 28366 28642 28418
rect 29262 28366 29314 28418
rect 30158 28366 30210 28418
rect 30494 28366 30546 28418
rect 30718 28366 30770 28418
rect 34974 28366 35026 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 5406 28030 5458 28082
rect 5630 28030 5682 28082
rect 11454 28030 11506 28082
rect 12350 28030 12402 28082
rect 12574 28030 12626 28082
rect 22878 28030 22930 28082
rect 23662 28030 23714 28082
rect 28590 28030 28642 28082
rect 5742 27918 5794 27970
rect 11902 27918 11954 27970
rect 21870 27918 21922 27970
rect 23102 27918 23154 27970
rect 23214 27918 23266 27970
rect 26014 27918 26066 27970
rect 41694 27918 41746 27970
rect 11678 27806 11730 27858
rect 12686 27806 12738 27858
rect 22654 27806 22706 27858
rect 25342 27806 25394 27858
rect 30158 27806 30210 27858
rect 41582 27806 41634 27858
rect 11454 27694 11506 27746
rect 13134 27694 13186 27746
rect 19742 27694 19794 27746
rect 28142 27694 28194 27746
rect 42254 27694 42306 27746
rect 41694 27582 41746 27634
rect 42142 27582 42194 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 5966 27134 6018 27186
rect 11342 27134 11394 27186
rect 12126 27134 12178 27186
rect 16606 27134 16658 27186
rect 41806 27134 41858 27186
rect 43934 27134 43986 27186
rect 9886 27022 9938 27074
rect 10446 27022 10498 27074
rect 10894 27022 10946 27074
rect 11566 27022 11618 27074
rect 17166 27022 17218 27074
rect 30830 27022 30882 27074
rect 31614 27022 31666 27074
rect 31950 27022 32002 27074
rect 37886 27022 37938 27074
rect 41022 27022 41074 27074
rect 30718 26910 30770 26962
rect 37550 26910 37602 26962
rect 40686 26910 40738 26962
rect 5854 26798 5906 26850
rect 6078 26798 6130 26850
rect 6302 26798 6354 26850
rect 11118 26798 11170 26850
rect 11342 26798 11394 26850
rect 30494 26798 30546 26850
rect 31838 26798 31890 26850
rect 37774 26798 37826 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 4062 26462 4114 26514
rect 12238 26462 12290 26514
rect 13022 26462 13074 26514
rect 13134 26462 13186 26514
rect 18734 26462 18786 26514
rect 33070 26462 33122 26514
rect 33294 26462 33346 26514
rect 36990 26462 37042 26514
rect 41694 26462 41746 26514
rect 5294 26350 5346 26402
rect 9886 26350 9938 26402
rect 11118 26350 11170 26402
rect 11902 26350 11954 26402
rect 15374 26350 15426 26402
rect 16606 26350 16658 26402
rect 17726 26350 17778 26402
rect 33518 26350 33570 26402
rect 36654 26350 36706 26402
rect 36766 26350 36818 26402
rect 41806 26350 41858 26402
rect 42030 26350 42082 26402
rect 4510 26238 4562 26290
rect 4622 26238 4674 26290
rect 4846 26238 4898 26290
rect 5406 26238 5458 26290
rect 5518 26238 5570 26290
rect 10558 26238 10610 26290
rect 10782 26238 10834 26290
rect 12910 26238 12962 26290
rect 13582 26238 13634 26290
rect 16270 26238 16322 26290
rect 17390 26238 17442 26290
rect 18398 26238 18450 26290
rect 36206 26238 36258 26290
rect 41470 26238 41522 26290
rect 9550 26126 9602 26178
rect 15150 26126 15202 26178
rect 32510 26126 32562 26178
rect 33182 26126 33234 26178
rect 35870 26126 35922 26178
rect 36654 26126 36706 26178
rect 41134 26126 41186 26178
rect 42254 26126 42306 26178
rect 5966 26014 6018 26066
rect 11006 26014 11058 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 13582 25678 13634 25730
rect 3614 25566 3666 25618
rect 4734 25566 4786 25618
rect 8318 25566 8370 25618
rect 22654 25566 22706 25618
rect 23102 25566 23154 25618
rect 25230 25566 25282 25618
rect 30494 25566 30546 25618
rect 35982 25566 36034 25618
rect 36430 25566 36482 25618
rect 39230 25566 39282 25618
rect 4398 25454 4450 25506
rect 4846 25454 4898 25506
rect 5966 25454 6018 25506
rect 6190 25454 6242 25506
rect 7198 25454 7250 25506
rect 7982 25454 8034 25506
rect 8206 25454 8258 25506
rect 11342 25454 11394 25506
rect 14142 25454 14194 25506
rect 14366 25454 14418 25506
rect 14590 25454 14642 25506
rect 16046 25454 16098 25506
rect 21646 25454 21698 25506
rect 23774 25454 23826 25506
rect 24222 25454 24274 25506
rect 24894 25454 24946 25506
rect 30606 25454 30658 25506
rect 30830 25454 30882 25506
rect 36990 25454 37042 25506
rect 39006 25454 39058 25506
rect 40910 25454 40962 25506
rect 3838 25342 3890 25394
rect 4622 25342 4674 25394
rect 5742 25342 5794 25394
rect 10782 25342 10834 25394
rect 11006 25342 11058 25394
rect 15710 25342 15762 25394
rect 21310 25342 21362 25394
rect 21422 25342 21474 25394
rect 26014 25342 26066 25394
rect 37326 25342 37378 25394
rect 39902 25342 39954 25394
rect 3726 25230 3778 25282
rect 4062 25230 4114 25282
rect 5070 25230 5122 25282
rect 6078 25230 6130 25282
rect 10670 25230 10722 25282
rect 18062 25230 18114 25282
rect 23438 25230 23490 25282
rect 24446 25230 24498 25282
rect 25678 25230 25730 25282
rect 31054 25230 31106 25282
rect 31278 25230 31330 25282
rect 36318 25230 36370 25282
rect 41134 25230 41186 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 4734 24894 4786 24946
rect 5070 24894 5122 24946
rect 5854 24894 5906 24946
rect 7870 24894 7922 24946
rect 8766 24894 8818 24946
rect 11118 24894 11170 24946
rect 15934 24894 15986 24946
rect 16382 24894 16434 24946
rect 25342 24894 25394 24946
rect 26238 24894 26290 24946
rect 27134 24894 27186 24946
rect 41022 24894 41074 24946
rect 4622 24782 4674 24834
rect 5294 24782 5346 24834
rect 7646 24782 7698 24834
rect 10110 24782 10162 24834
rect 10558 24782 10610 24834
rect 23886 24782 23938 24834
rect 31950 24782 32002 24834
rect 36206 24782 36258 24834
rect 40910 24782 40962 24834
rect 5406 24670 5458 24722
rect 8094 24670 8146 24722
rect 8318 24670 8370 24722
rect 16158 24670 16210 24722
rect 16606 24670 16658 24722
rect 16830 24670 16882 24722
rect 17390 24670 17442 24722
rect 24222 24670 24274 24722
rect 25902 24670 25954 24722
rect 31278 24670 31330 24722
rect 31614 24670 31666 24722
rect 35534 24670 35586 24722
rect 38782 24670 38834 24722
rect 41246 24670 41298 24722
rect 17950 24558 18002 24610
rect 23998 24558 24050 24610
rect 24670 24558 24722 24610
rect 26686 24558 26738 24610
rect 27582 24558 27634 24610
rect 31502 24558 31554 24610
rect 38334 24558 38386 24610
rect 4846 24446 4898 24498
rect 7758 24446 7810 24498
rect 10222 24446 10274 24498
rect 10670 24446 10722 24498
rect 17726 24446 17778 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 7198 24110 7250 24162
rect 21534 24110 21586 24162
rect 7758 23998 7810 24050
rect 17950 23998 18002 24050
rect 20862 23998 20914 24050
rect 29934 23998 29986 24050
rect 32062 23998 32114 24050
rect 32398 23998 32450 24050
rect 34526 23998 34578 24050
rect 40910 23998 40962 24050
rect 6190 23886 6242 23938
rect 6750 23886 6802 23938
rect 18286 23886 18338 23938
rect 18510 23886 18562 23938
rect 19630 23886 19682 23938
rect 21534 23886 21586 23938
rect 22094 23886 22146 23938
rect 22430 23886 22482 23938
rect 22542 23886 22594 23938
rect 23102 23886 23154 23938
rect 25454 23886 25506 23938
rect 26014 23886 26066 23938
rect 29262 23886 29314 23938
rect 35310 23886 35362 23938
rect 35870 23886 35922 23938
rect 41246 23886 41298 23938
rect 6526 23774 6578 23826
rect 7086 23774 7138 23826
rect 7198 23774 7250 23826
rect 18734 23774 18786 23826
rect 21870 23774 21922 23826
rect 22654 23774 22706 23826
rect 41470 23774 41522 23826
rect 41582 23774 41634 23826
rect 41694 23774 41746 23826
rect 6302 23662 6354 23714
rect 19966 23662 20018 23714
rect 21982 23662 22034 23714
rect 41358 23662 41410 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 4958 23326 5010 23378
rect 31166 23326 31218 23378
rect 32398 23326 32450 23378
rect 34638 23326 34690 23378
rect 14366 23214 14418 23266
rect 15262 23214 15314 23266
rect 20190 23214 20242 23266
rect 31278 23214 31330 23266
rect 41806 23214 41858 23266
rect 5294 23102 5346 23154
rect 14478 23102 14530 23154
rect 14926 23102 14978 23154
rect 18622 23102 18674 23154
rect 19518 23102 19570 23154
rect 34862 23102 34914 23154
rect 18510 22990 18562 23042
rect 21198 22990 21250 23042
rect 35422 22990 35474 23042
rect 16046 22878 16098 22930
rect 17838 22878 17890 22930
rect 41694 22878 41746 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 16830 22542 16882 22594
rect 2606 22430 2658 22482
rect 4734 22430 4786 22482
rect 9998 22430 10050 22482
rect 16270 22430 16322 22482
rect 16494 22430 16546 22482
rect 17166 22430 17218 22482
rect 41582 22430 41634 22482
rect 43710 22430 43762 22482
rect 1934 22318 1986 22370
rect 7086 22318 7138 22370
rect 8654 22318 8706 22370
rect 17726 22318 17778 22370
rect 21534 22318 21586 22370
rect 21758 22318 21810 22370
rect 40910 22318 40962 22370
rect 5742 22206 5794 22258
rect 7870 22206 7922 22258
rect 8766 22206 8818 22258
rect 26798 22206 26850 22258
rect 40462 22094 40514 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 7534 21758 7586 21810
rect 11454 21758 11506 21810
rect 15822 21758 15874 21810
rect 10446 21646 10498 21698
rect 11566 21646 11618 21698
rect 12686 21646 12738 21698
rect 13694 21646 13746 21698
rect 22206 21646 22258 21698
rect 6414 21534 6466 21586
rect 7422 21534 7474 21586
rect 10782 21534 10834 21586
rect 11790 21534 11842 21586
rect 12126 21534 12178 21586
rect 13806 21534 13858 21586
rect 16494 21534 16546 21586
rect 22990 21534 23042 21586
rect 36094 21534 36146 21586
rect 6526 21422 6578 21474
rect 15374 21422 15426 21474
rect 20078 21422 20130 21474
rect 23550 21422 23602 21474
rect 36878 21422 36930 21474
rect 39006 21422 39058 21474
rect 39454 21422 39506 21474
rect 16270 21310 16322 21362
rect 16606 21310 16658 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 34638 20974 34690 21026
rect 8318 20862 8370 20914
rect 13806 20862 13858 20914
rect 37326 20862 37378 20914
rect 8206 20750 8258 20802
rect 9102 20750 9154 20802
rect 9998 20750 10050 20802
rect 10558 20750 10610 20802
rect 11454 20750 11506 20802
rect 12686 20750 12738 20802
rect 13470 20750 13522 20802
rect 14926 20750 14978 20802
rect 16942 20750 16994 20802
rect 17390 20750 17442 20802
rect 37550 20750 37602 20802
rect 7758 20638 7810 20690
rect 9886 20638 9938 20690
rect 11342 20638 11394 20690
rect 13918 20638 13970 20690
rect 15374 20638 15426 20690
rect 17950 20638 18002 20690
rect 34974 20638 35026 20690
rect 35198 20638 35250 20690
rect 35422 20638 35474 20690
rect 37214 20638 37266 20690
rect 8990 20526 9042 20578
rect 10558 20526 10610 20578
rect 10670 20526 10722 20578
rect 12350 20526 12402 20578
rect 12574 20526 12626 20578
rect 14702 20526 14754 20578
rect 16942 20526 16994 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 5406 20190 5458 20242
rect 34974 20190 35026 20242
rect 3166 20078 3218 20130
rect 5966 20078 6018 20130
rect 7758 20078 7810 20130
rect 16718 20078 16770 20130
rect 22654 20078 22706 20130
rect 35422 20078 35474 20130
rect 35646 20078 35698 20130
rect 2382 19966 2434 20018
rect 7086 19966 7138 20018
rect 7534 19966 7586 20018
rect 12126 19966 12178 20018
rect 12910 19966 12962 20018
rect 13806 19966 13858 20018
rect 14254 19966 14306 20018
rect 22878 19966 22930 20018
rect 25790 19966 25842 20018
rect 29934 19966 29986 20018
rect 31390 19966 31442 20018
rect 35982 19966 36034 20018
rect 9998 19854 10050 19906
rect 11790 19854 11842 19906
rect 15262 19854 15314 19906
rect 16158 19854 16210 19906
rect 26574 19854 26626 19906
rect 28702 19854 28754 19906
rect 30046 19854 30098 19906
rect 31950 19854 32002 19906
rect 10110 19742 10162 19794
rect 22878 19742 22930 19794
rect 23214 19742 23266 19794
rect 29262 19742 29314 19794
rect 31726 19742 31778 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 26686 19406 26738 19458
rect 38894 19406 38946 19458
rect 23662 19294 23714 19346
rect 25790 19294 25842 19346
rect 26574 19294 26626 19346
rect 27134 19294 27186 19346
rect 29262 19294 29314 19346
rect 30046 19294 30098 19346
rect 35422 19294 35474 19346
rect 37550 19294 37602 19346
rect 8318 19182 8370 19234
rect 9102 19182 9154 19234
rect 9438 19182 9490 19234
rect 11678 19182 11730 19234
rect 16270 19182 16322 19234
rect 22990 19182 23042 19234
rect 26350 19182 26402 19234
rect 30382 19182 30434 19234
rect 30718 19182 30770 19234
rect 31502 19182 31554 19234
rect 32062 19182 32114 19234
rect 34078 19182 34130 19234
rect 37998 19182 38050 19234
rect 38334 19182 38386 19234
rect 38670 19182 38722 19234
rect 10894 19070 10946 19122
rect 16494 19070 16546 19122
rect 17278 19070 17330 19122
rect 32174 19070 32226 19122
rect 34638 19070 34690 19122
rect 11902 18958 11954 19010
rect 16606 18958 16658 19010
rect 30606 18958 30658 19010
rect 31166 18958 31218 19010
rect 31390 18958 31442 19010
rect 31614 18958 31666 19010
rect 39230 18958 39282 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 16158 18510 16210 18562
rect 16494 18510 16546 18562
rect 31614 18510 31666 18562
rect 14926 18398 14978 18450
rect 15374 18398 15426 18450
rect 21646 18398 21698 18450
rect 22094 18398 22146 18450
rect 32398 18398 32450 18450
rect 35758 18398 35810 18450
rect 39118 18398 39170 18450
rect 41806 18398 41858 18450
rect 10110 18286 10162 18338
rect 18734 18286 18786 18338
rect 20862 18286 20914 18338
rect 26014 18286 26066 18338
rect 29486 18286 29538 18338
rect 33182 18286 33234 18338
rect 36542 18286 36594 18338
rect 38670 18286 38722 18338
rect 41694 18286 41746 18338
rect 41470 18174 41522 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 8878 17838 8930 17890
rect 12350 17838 12402 17890
rect 36990 17838 37042 17890
rect 37326 17838 37378 17890
rect 10558 17726 10610 17778
rect 12238 17726 12290 17778
rect 19518 17726 19570 17778
rect 20190 17726 20242 17778
rect 39566 17726 39618 17778
rect 40014 17726 40066 17778
rect 41694 17726 41746 17778
rect 43822 17726 43874 17778
rect 9662 17614 9714 17666
rect 9886 17614 9938 17666
rect 10110 17614 10162 17666
rect 16158 17614 16210 17666
rect 19742 17614 19794 17666
rect 37102 17614 37154 17666
rect 37550 17614 37602 17666
rect 40686 17614 40738 17666
rect 40910 17614 40962 17666
rect 8990 17502 9042 17554
rect 9998 17502 10050 17554
rect 10670 17502 10722 17554
rect 19406 17502 19458 17554
rect 40350 17502 40402 17554
rect 40462 17502 40514 17554
rect 9214 17390 9266 17442
rect 15822 17390 15874 17442
rect 17054 17390 17106 17442
rect 36430 17390 36482 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 6974 17054 7026 17106
rect 9886 17054 9938 17106
rect 10334 17054 10386 17106
rect 11118 17054 11170 17106
rect 13134 17054 13186 17106
rect 40238 17054 40290 17106
rect 41470 17054 41522 17106
rect 4398 16942 4450 16994
rect 11902 16942 11954 16994
rect 13806 16942 13858 16994
rect 14030 16942 14082 16994
rect 14142 16942 14194 16994
rect 17390 16942 17442 16994
rect 40126 16942 40178 16994
rect 41246 16942 41298 16994
rect 3614 16830 3666 16882
rect 9550 16830 9602 16882
rect 10222 16830 10274 16882
rect 11118 16830 11170 16882
rect 11566 16830 11618 16882
rect 13358 16830 13410 16882
rect 13694 16830 13746 16882
rect 15710 16830 15762 16882
rect 16158 16830 16210 16882
rect 17950 16830 18002 16882
rect 33182 16830 33234 16882
rect 33518 16830 33570 16882
rect 40462 16830 40514 16882
rect 6526 16718 6578 16770
rect 16606 16718 16658 16770
rect 38110 16718 38162 16770
rect 41582 16718 41634 16770
rect 11454 16606 11506 16658
rect 13022 16606 13074 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 9550 16270 9602 16322
rect 2606 16158 2658 16210
rect 4734 16158 4786 16210
rect 5742 16158 5794 16210
rect 9102 16158 9154 16210
rect 12350 16158 12402 16210
rect 19294 16158 19346 16210
rect 23214 16158 23266 16210
rect 24222 16158 24274 16210
rect 31950 16158 32002 16210
rect 1934 16046 1986 16098
rect 8990 16046 9042 16098
rect 9774 16046 9826 16098
rect 12126 16046 12178 16098
rect 12462 16046 12514 16098
rect 12686 16046 12738 16098
rect 17278 16046 17330 16098
rect 25006 16046 25058 16098
rect 29374 16046 29426 16098
rect 9214 15934 9266 15986
rect 12238 15934 12290 15986
rect 15822 15934 15874 15986
rect 23326 15934 23378 15986
rect 23550 15934 23602 15986
rect 24558 15934 24610 15986
rect 24670 15934 24722 15986
rect 24894 15934 24946 15986
rect 25454 15934 25506 15986
rect 25678 15934 25730 15986
rect 26350 15934 26402 15986
rect 22990 15822 23042 15874
rect 23102 15822 23154 15874
rect 25342 15822 25394 15874
rect 26014 15822 26066 15874
rect 28702 15822 28754 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 9886 15486 9938 15538
rect 9998 15486 10050 15538
rect 12910 15486 12962 15538
rect 17726 15486 17778 15538
rect 17838 15486 17890 15538
rect 19518 15486 19570 15538
rect 20862 15486 20914 15538
rect 22430 15486 22482 15538
rect 23102 15486 23154 15538
rect 24446 15486 24498 15538
rect 24558 15486 24610 15538
rect 29262 15486 29314 15538
rect 33406 15486 33458 15538
rect 9774 15374 9826 15426
rect 17390 15374 17442 15426
rect 18846 15374 18898 15426
rect 19966 15374 20018 15426
rect 21870 15374 21922 15426
rect 28030 15374 28082 15426
rect 33070 15374 33122 15426
rect 9550 15262 9602 15314
rect 10110 15262 10162 15314
rect 17614 15262 17666 15314
rect 18062 15262 18114 15314
rect 18622 15262 18674 15314
rect 19182 15262 19234 15314
rect 21086 15262 21138 15314
rect 22094 15262 22146 15314
rect 22766 15262 22818 15314
rect 23102 15262 23154 15314
rect 23326 15262 23378 15314
rect 23886 15262 23938 15314
rect 24222 15262 24274 15314
rect 28814 15262 28866 15314
rect 29598 15262 29650 15314
rect 34862 15262 34914 15314
rect 20414 15150 20466 15202
rect 25902 15150 25954 15202
rect 30382 15150 30434 15202
rect 32510 15150 32562 15202
rect 35534 15150 35586 15202
rect 37662 15150 37714 15202
rect 38110 15150 38162 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 16270 14702 16322 14754
rect 23550 14702 23602 14754
rect 23886 14702 23938 14754
rect 11006 14590 11058 14642
rect 16494 14590 16546 14642
rect 17054 14590 17106 14642
rect 18062 14590 18114 14642
rect 18846 14590 18898 14642
rect 19294 14590 19346 14642
rect 31502 14590 31554 14642
rect 32734 14590 32786 14642
rect 11342 14478 11394 14530
rect 14926 14478 14978 14530
rect 15486 14478 15538 14530
rect 15934 14478 15986 14530
rect 17726 14478 17778 14530
rect 18174 14478 18226 14530
rect 23886 14478 23938 14530
rect 31726 14478 31778 14530
rect 36430 14478 36482 14530
rect 37550 14478 37602 14530
rect 41246 14478 41298 14530
rect 8654 14366 8706 14418
rect 11678 14366 11730 14418
rect 14590 14366 14642 14418
rect 31390 14366 31442 14418
rect 31950 14366 32002 14418
rect 37662 14366 37714 14418
rect 41358 14366 41410 14418
rect 8766 14254 8818 14306
rect 15262 14254 15314 14306
rect 17390 14254 17442 14306
rect 36094 14254 36146 14306
rect 39006 14254 39058 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 14814 13918 14866 13970
rect 15598 13918 15650 13970
rect 16718 13918 16770 13970
rect 27246 13918 27298 13970
rect 31950 13918 32002 13970
rect 36094 13918 36146 13970
rect 39902 13918 39954 13970
rect 8542 13806 8594 13858
rect 9550 13806 9602 13858
rect 21534 13806 21586 13858
rect 21646 13806 21698 13858
rect 23998 13806 24050 13858
rect 24110 13806 24162 13858
rect 26350 13806 26402 13858
rect 28814 13806 28866 13858
rect 37438 13806 37490 13858
rect 8654 13694 8706 13746
rect 9774 13694 9826 13746
rect 10222 13694 10274 13746
rect 24222 13694 24274 13746
rect 26238 13694 26290 13746
rect 28366 13694 28418 13746
rect 31614 13694 31666 13746
rect 31838 13694 31890 13746
rect 32062 13694 32114 13746
rect 32398 13694 32450 13746
rect 35758 13694 35810 13746
rect 35870 13694 35922 13746
rect 36206 13694 36258 13746
rect 36542 13694 36594 13746
rect 36766 13694 36818 13746
rect 37214 13694 37266 13746
rect 37326 13694 37378 13746
rect 41022 13694 41074 13746
rect 9662 13582 9714 13634
rect 15150 13582 15202 13634
rect 40350 13582 40402 13634
rect 41806 13582 41858 13634
rect 43934 13582 43986 13634
rect 8542 13470 8594 13522
rect 9998 13470 10050 13522
rect 21646 13470 21698 13522
rect 24670 13470 24722 13522
rect 31390 13470 31442 13522
rect 31614 13470 31666 13522
rect 40238 13470 40290 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 10446 13134 10498 13186
rect 9214 13022 9266 13074
rect 11118 13022 11170 13074
rect 40126 13022 40178 13074
rect 7982 12910 8034 12962
rect 8654 12910 8706 12962
rect 10222 12910 10274 12962
rect 10446 12910 10498 12962
rect 21870 12910 21922 12962
rect 22094 12910 22146 12962
rect 40798 12910 40850 12962
rect 41022 12910 41074 12962
rect 8878 12798 8930 12850
rect 9886 12798 9938 12850
rect 11454 12798 11506 12850
rect 11678 12798 11730 12850
rect 21646 12798 21698 12850
rect 23214 12798 23266 12850
rect 40238 12798 40290 12850
rect 40462 12798 40514 12850
rect 41358 12798 41410 12850
rect 41694 12798 41746 12850
rect 42030 12798 42082 12850
rect 8094 12686 8146 12738
rect 9102 12686 9154 12738
rect 9214 12686 9266 12738
rect 10222 12686 10274 12738
rect 11118 12686 11170 12738
rect 11230 12686 11282 12738
rect 21982 12686 22034 12738
rect 22878 12686 22930 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 6414 12350 6466 12402
rect 13134 12350 13186 12402
rect 22766 12350 22818 12402
rect 37662 12350 37714 12402
rect 38446 12350 38498 12402
rect 40798 12350 40850 12402
rect 41022 12350 41074 12402
rect 4174 12238 4226 12290
rect 8878 12238 8930 12290
rect 10110 12238 10162 12290
rect 11118 12238 11170 12290
rect 21310 12238 21362 12290
rect 21534 12238 21586 12290
rect 21646 12238 21698 12290
rect 21758 12238 21810 12290
rect 38110 12238 38162 12290
rect 3502 12126 3554 12178
rect 8542 12126 8594 12178
rect 9550 12126 9602 12178
rect 11230 12126 11282 12178
rect 21870 12126 21922 12178
rect 22206 12126 22258 12178
rect 37438 12126 37490 12178
rect 41134 12126 41186 12178
rect 6974 12014 7026 12066
rect 8766 12014 8818 12066
rect 12910 12014 12962 12066
rect 13694 12014 13746 12066
rect 37102 12014 37154 12066
rect 22430 11902 22482 11954
rect 37774 11902 37826 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 12798 11566 12850 11618
rect 13022 11566 13074 11618
rect 25566 11566 25618 11618
rect 4846 11454 4898 11506
rect 5742 11454 5794 11506
rect 21310 11454 21362 11506
rect 22206 11454 22258 11506
rect 24558 11454 24610 11506
rect 1934 11342 1986 11394
rect 2606 11342 2658 11394
rect 8766 11342 8818 11394
rect 9102 11342 9154 11394
rect 17166 11342 17218 11394
rect 17726 11342 17778 11394
rect 25454 11342 25506 11394
rect 31614 11342 31666 11394
rect 31838 11342 31890 11394
rect 32734 11342 32786 11394
rect 32958 11342 33010 11394
rect 35870 11342 35922 11394
rect 36206 11342 36258 11394
rect 36430 11342 36482 11394
rect 37438 11342 37490 11394
rect 37550 11342 37602 11394
rect 37662 11342 37714 11394
rect 12126 11230 12178 11282
rect 21422 11230 21474 11282
rect 21646 11230 21698 11282
rect 25118 11230 25170 11282
rect 26014 11230 26066 11282
rect 26350 11230 26402 11282
rect 31278 11230 31330 11282
rect 32622 11230 32674 11282
rect 8878 11118 8930 11170
rect 11790 11118 11842 11170
rect 17278 11118 17330 11170
rect 17390 11118 17442 11170
rect 17502 11118 17554 11170
rect 24782 11118 24834 11170
rect 25006 11118 25058 11170
rect 25566 11118 25618 11170
rect 26126 11118 26178 11170
rect 31502 11118 31554 11170
rect 32174 11118 32226 11170
rect 34190 11118 34242 11170
rect 34526 11118 34578 11170
rect 35982 11118 36034 11170
rect 36990 11118 37042 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 8430 10782 8482 10834
rect 9886 10782 9938 10834
rect 9998 10782 10050 10834
rect 10670 10782 10722 10834
rect 12462 10782 12514 10834
rect 13022 10782 13074 10834
rect 16270 10782 16322 10834
rect 17614 10782 17666 10834
rect 24446 10782 24498 10834
rect 24670 10782 24722 10834
rect 25566 10782 25618 10834
rect 25790 10782 25842 10834
rect 26686 10782 26738 10834
rect 33182 10782 33234 10834
rect 35086 10782 35138 10834
rect 35870 10782 35922 10834
rect 9550 10670 9602 10722
rect 12574 10670 12626 10722
rect 13582 10670 13634 10722
rect 18398 10670 18450 10722
rect 20862 10670 20914 10722
rect 24222 10670 24274 10722
rect 25342 10670 25394 10722
rect 27022 10670 27074 10722
rect 7870 10558 7922 10610
rect 8206 10558 8258 10610
rect 9774 10558 9826 10610
rect 10222 10558 10274 10610
rect 12238 10558 12290 10610
rect 13918 10558 13970 10610
rect 18286 10558 18338 10610
rect 20302 10558 20354 10610
rect 29710 10558 29762 10610
rect 35534 10558 35586 10610
rect 35758 10558 35810 10610
rect 35982 10558 36034 10610
rect 8318 10446 8370 10498
rect 8878 10446 8930 10498
rect 15262 10446 15314 10498
rect 21646 10446 21698 10498
rect 24670 10446 24722 10498
rect 25454 10446 25506 10498
rect 30382 10446 30434 10498
rect 32510 10446 32562 10498
rect 8654 10334 8706 10386
rect 9102 10334 9154 10386
rect 13918 10334 13970 10386
rect 17278 10334 17330 10386
rect 18062 10334 18114 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 8430 9998 8482 10050
rect 17166 9998 17218 10050
rect 17838 9998 17890 10050
rect 19854 9998 19906 10050
rect 20414 9998 20466 10050
rect 31278 9998 31330 10050
rect 31614 9998 31666 10050
rect 8094 9886 8146 9938
rect 12686 9886 12738 9938
rect 24894 9886 24946 9938
rect 26462 9886 26514 9938
rect 28590 9886 28642 9938
rect 29262 9886 29314 9938
rect 7534 9774 7586 9826
rect 12238 9774 12290 9826
rect 12462 9774 12514 9826
rect 12910 9774 12962 9826
rect 14366 9774 14418 9826
rect 15038 9774 15090 9826
rect 15486 9774 15538 9826
rect 15598 9774 15650 9826
rect 16606 9774 16658 9826
rect 16942 9774 16994 9826
rect 17390 9774 17442 9826
rect 17614 9774 17666 9826
rect 19070 9774 19122 9826
rect 19294 9774 19346 9826
rect 19630 9774 19682 9826
rect 19854 9774 19906 9826
rect 24782 9774 24834 9826
rect 25118 9774 25170 9826
rect 25342 9774 25394 9826
rect 25790 9774 25842 9826
rect 31390 9774 31442 9826
rect 31838 9774 31890 9826
rect 8654 9662 8706 9714
rect 12014 9662 12066 9714
rect 16046 9662 16098 9714
rect 20526 9662 20578 9714
rect 8542 9550 8594 9602
rect 12350 9550 12402 9602
rect 13582 9550 13634 9602
rect 14814 9550 14866 9602
rect 14926 9550 14978 9602
rect 15710 9550 15762 9602
rect 15822 9550 15874 9602
rect 16830 9550 16882 9602
rect 17950 9550 18002 9602
rect 18174 9550 18226 9602
rect 19630 9550 19682 9602
rect 30942 9550 30994 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 12238 9214 12290 9266
rect 12350 9214 12402 9266
rect 14814 9102 14866 9154
rect 15598 9102 15650 9154
rect 15710 9102 15762 9154
rect 16494 9158 16546 9210
rect 17390 9214 17442 9266
rect 18174 9214 18226 9266
rect 20190 9214 20242 9266
rect 21086 9214 21138 9266
rect 23998 9214 24050 9266
rect 17950 9102 18002 9154
rect 20078 9102 20130 9154
rect 24334 9102 24386 9154
rect 24558 9102 24610 9154
rect 26126 9102 26178 9154
rect 26462 9102 26514 9154
rect 26574 9102 26626 9154
rect 35758 9102 35810 9154
rect 12126 8990 12178 9042
rect 12798 8990 12850 9042
rect 15150 8990 15202 9042
rect 16718 8990 16770 9042
rect 17838 8990 17890 9042
rect 20414 8990 20466 9042
rect 20638 8990 20690 9042
rect 25118 8990 25170 9042
rect 25454 8990 25506 9042
rect 25678 8990 25730 9042
rect 25902 8990 25954 9042
rect 35086 8990 35138 9042
rect 38334 8990 38386 9042
rect 14926 8878 14978 8930
rect 17502 8878 17554 8930
rect 24670 8878 24722 8930
rect 26014 8878 26066 8930
rect 37886 8878 37938 8930
rect 15710 8766 15762 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 5630 8318 5682 8370
rect 7758 8318 7810 8370
rect 9102 8318 9154 8370
rect 25006 8318 25058 8370
rect 8542 8206 8594 8258
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 9662 6750 9714 6802
rect 11790 6638 11842 6690
rect 12574 6638 12626 6690
rect 21646 6638 21698 6690
rect 18062 6526 18114 6578
rect 18398 6526 18450 6578
rect 13582 6414 13634 6466
rect 21758 6414 21810 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 18622 6078 18674 6130
rect 28590 6078 28642 6130
rect 19070 5966 19122 6018
rect 21086 5966 21138 6018
rect 26014 5966 26066 6018
rect 18510 5854 18562 5906
rect 22206 5854 22258 5906
rect 25342 5854 25394 5906
rect 28142 5742 28194 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 16494 5182 16546 5234
rect 18622 5182 18674 5234
rect 21310 5182 21362 5234
rect 23438 5182 23490 5234
rect 24782 5182 24834 5234
rect 15374 5070 15426 5122
rect 15822 5070 15874 5122
rect 24110 5070 24162 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 16830 4510 16882 4562
rect 18734 4510 18786 4562
rect 14254 4398 14306 4450
rect 19854 4398 19906 4450
rect 13582 4286 13634 4338
rect 19182 4286 19234 4338
rect 16382 4174 16434 4226
rect 21982 4174 22034 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 1792 45200 1904 46000
rect 5600 45200 5712 46000
rect 9408 45200 9520 46000
rect 13216 45200 13328 46000
rect 17024 45200 17136 46000
rect 17388 45276 17892 45332
rect 1820 43708 1876 45200
rect 1820 43652 2324 43708
rect 1932 38834 1988 38846
rect 1932 38782 1934 38834
rect 1986 38782 1988 38834
rect 1932 35698 1988 38782
rect 1932 35646 1934 35698
rect 1986 35646 1988 35698
rect 1932 34020 1988 35646
rect 1932 33954 1988 33964
rect 2156 31778 2212 31790
rect 2156 31726 2158 31778
rect 2210 31726 2212 31778
rect 2156 31556 2212 31726
rect 1932 29428 1988 29438
rect 2156 29428 2212 31500
rect 1932 29426 2212 29428
rect 1932 29374 1934 29426
rect 1986 29374 2212 29426
rect 1932 29372 2212 29374
rect 1932 29362 1988 29372
rect 1932 22370 1988 22382
rect 1932 22318 1934 22370
rect 1986 22318 1988 22370
rect 1932 22260 1988 22318
rect 1932 20020 1988 22204
rect 2268 22148 2324 43652
rect 5628 43092 5684 45200
rect 5628 43036 5908 43092
rect 5068 41972 5124 41982
rect 5852 41972 5908 43036
rect 5068 41970 5908 41972
rect 5068 41918 5070 41970
rect 5122 41918 5854 41970
rect 5906 41918 5908 41970
rect 5068 41916 5908 41918
rect 5068 41906 5124 41916
rect 5852 41906 5908 41916
rect 6188 42082 6244 42094
rect 6188 42030 6190 42082
rect 6242 42030 6244 42082
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 5180 40964 5236 40974
rect 3052 40404 3108 40414
rect 3276 40404 3332 40414
rect 3052 40402 3276 40404
rect 3052 40350 3054 40402
rect 3106 40350 3276 40402
rect 3052 40348 3276 40350
rect 3052 40338 3108 40348
rect 3276 40338 3332 40348
rect 5180 40404 5236 40908
rect 3724 40292 3780 40302
rect 3724 40198 3780 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5180 39058 5236 40348
rect 6188 40404 6244 42030
rect 8876 41972 8932 41982
rect 9436 41972 9492 45200
rect 9996 42082 10052 42094
rect 9996 42030 9998 42082
rect 10050 42030 10052 42082
rect 9660 41972 9716 41982
rect 8876 41970 9716 41972
rect 8876 41918 8878 41970
rect 8930 41918 9662 41970
rect 9714 41918 9716 41970
rect 8876 41916 9716 41918
rect 8876 41906 8932 41916
rect 9660 41906 9716 41916
rect 6300 40964 6356 40974
rect 6300 40626 6356 40908
rect 6300 40574 6302 40626
rect 6354 40574 6356 40626
rect 6300 40562 6356 40574
rect 6188 40338 6244 40348
rect 8092 40516 8148 40526
rect 5852 40290 5908 40302
rect 5852 40238 5854 40290
rect 5906 40238 5908 40290
rect 5852 40180 5908 40238
rect 5852 40114 5908 40124
rect 6412 40292 6468 40302
rect 6412 39730 6468 40236
rect 6412 39678 6414 39730
rect 6466 39678 6468 39730
rect 6412 39666 6468 39678
rect 6972 39618 7028 39630
rect 6972 39566 6974 39618
rect 7026 39566 7028 39618
rect 6972 39508 7028 39566
rect 7756 39620 7812 39630
rect 7980 39620 8036 39630
rect 7756 39618 8036 39620
rect 7756 39566 7758 39618
rect 7810 39566 7982 39618
rect 8034 39566 8036 39618
rect 7756 39564 8036 39566
rect 6972 39442 7028 39452
rect 7644 39508 7700 39518
rect 7644 39414 7700 39452
rect 6300 39396 6356 39406
rect 6300 39302 6356 39340
rect 6524 39394 6580 39406
rect 6524 39342 6526 39394
rect 6578 39342 6580 39394
rect 5180 39006 5182 39058
rect 5234 39006 5236 39058
rect 2604 38948 2660 38958
rect 2604 38854 2660 38892
rect 4732 38724 4788 38734
rect 4732 38722 4900 38724
rect 4732 38670 4734 38722
rect 4786 38670 4900 38722
rect 4732 38668 4900 38670
rect 4732 38658 4788 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 2604 35812 2660 35822
rect 2604 35718 2660 35756
rect 4732 35586 4788 35598
rect 4732 35534 4734 35586
rect 4786 35534 4788 35586
rect 4732 35476 4788 35534
rect 4732 35410 4788 35420
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4844 35028 4900 38668
rect 4844 34962 4900 34972
rect 4956 36260 5012 36270
rect 4956 34242 5012 36204
rect 4956 34190 4958 34242
rect 5010 34190 5012 34242
rect 4956 34178 5012 34190
rect 5180 35586 5236 39006
rect 6524 38668 6580 39342
rect 7308 39394 7364 39406
rect 7308 39342 7310 39394
rect 7362 39342 7364 39394
rect 7308 39060 7364 39342
rect 7532 39396 7588 39406
rect 7532 39302 7588 39340
rect 7756 39172 7812 39564
rect 7980 39554 8036 39564
rect 7308 38668 7364 39004
rect 6524 38612 7364 38668
rect 7644 39116 7812 39172
rect 7644 38946 7700 39116
rect 7868 39060 7924 39070
rect 7644 38894 7646 38946
rect 7698 38894 7700 38946
rect 6860 37490 6916 38612
rect 6860 37438 6862 37490
rect 6914 37438 6916 37490
rect 6860 37426 6916 37438
rect 5180 35534 5182 35586
rect 5234 35534 5236 35586
rect 4284 34130 4340 34142
rect 4284 34078 4286 34130
rect 4338 34078 4340 34130
rect 4284 34020 4340 34078
rect 4284 33954 4340 33964
rect 5180 34020 5236 35534
rect 7084 37266 7140 37278
rect 7084 37214 7086 37266
rect 7138 37214 7140 37266
rect 7084 36370 7140 37214
rect 7084 36318 7086 36370
rect 7138 36318 7140 36370
rect 7084 34804 7140 36318
rect 7196 36260 7252 36270
rect 7196 36166 7252 36204
rect 7644 35812 7700 38894
rect 7756 38948 7812 38958
rect 7868 38948 7924 39004
rect 7980 39060 8036 39070
rect 8092 39060 8148 40460
rect 8764 40404 8820 40414
rect 9996 40404 10052 42030
rect 13244 41972 13300 45200
rect 17052 45108 17108 45200
rect 17388 45108 17444 45276
rect 17052 45052 17444 45108
rect 17836 43708 17892 45276
rect 20832 45200 20944 46000
rect 24640 45200 24752 46000
rect 28448 45200 28560 46000
rect 32256 45200 32368 46000
rect 32620 45276 33124 45332
rect 17836 43652 18340 43708
rect 18284 42194 18340 43652
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 18284 42142 18286 42194
rect 18338 42142 18340 42194
rect 18284 42130 18340 42142
rect 13244 41906 13300 41916
rect 13468 41970 13524 41982
rect 13468 41918 13470 41970
rect 13522 41918 13524 41970
rect 10780 40964 10836 40974
rect 10444 40628 10500 40638
rect 10444 40534 10500 40572
rect 10220 40516 10276 40526
rect 10220 40422 10276 40460
rect 8316 39396 8372 39406
rect 8316 39302 8372 39340
rect 8540 39394 8596 39406
rect 8540 39342 8542 39394
rect 8594 39342 8596 39394
rect 7980 39058 8148 39060
rect 7980 39006 7982 39058
rect 8034 39006 8148 39058
rect 7980 39004 8148 39006
rect 8540 39060 8596 39342
rect 8652 39396 8708 39406
rect 8652 39302 8708 39340
rect 7980 38994 8036 39004
rect 8540 38994 8596 39004
rect 7756 38946 7924 38948
rect 7756 38894 7758 38946
rect 7810 38894 7924 38946
rect 7756 38892 7924 38894
rect 7756 38882 7812 38892
rect 7644 35718 7700 35756
rect 7980 35698 8036 35710
rect 7980 35646 7982 35698
rect 8034 35646 8036 35698
rect 7980 35140 8036 35646
rect 7980 35074 8036 35084
rect 8764 34916 8820 40348
rect 9436 40348 10052 40404
rect 10108 40402 10164 40414
rect 10108 40350 10110 40402
rect 10162 40350 10164 40402
rect 9100 39842 9156 39854
rect 9100 39790 9102 39842
rect 9154 39790 9156 39842
rect 9100 39732 9156 39790
rect 9100 39666 9156 39676
rect 9212 39620 9268 39630
rect 9212 39526 9268 39564
rect 9100 39394 9156 39406
rect 9100 39342 9102 39394
rect 9154 39342 9156 39394
rect 9100 39172 9156 39342
rect 9100 39106 9156 39116
rect 8876 38948 8932 38958
rect 8876 38854 8932 38892
rect 8988 38836 9044 38846
rect 8988 38742 9044 38780
rect 9324 35476 9380 35486
rect 8764 34914 9268 34916
rect 8764 34862 8766 34914
rect 8818 34862 9268 34914
rect 8764 34860 9268 34862
rect 8764 34850 8820 34860
rect 7084 34738 7140 34748
rect 9100 34690 9156 34702
rect 9100 34638 9102 34690
rect 9154 34638 9156 34690
rect 9100 34580 9156 34638
rect 9100 34514 9156 34524
rect 9212 34356 9268 34860
rect 9324 34914 9380 35420
rect 9324 34862 9326 34914
rect 9378 34862 9380 34914
rect 9324 34850 9380 34862
rect 9436 34580 9492 40348
rect 10108 39844 10164 40350
rect 10780 40402 10836 40908
rect 10780 40350 10782 40402
rect 10834 40350 10836 40402
rect 10780 40338 10836 40350
rect 11452 40292 11508 40302
rect 11340 40290 11508 40292
rect 11340 40238 11454 40290
rect 11506 40238 11508 40290
rect 11340 40236 11508 40238
rect 10108 39778 10164 39788
rect 11228 39844 11284 39854
rect 9660 39618 9716 39630
rect 9660 39566 9662 39618
rect 9714 39566 9716 39618
rect 9548 39172 9604 39182
rect 9548 39058 9604 39116
rect 9548 39006 9550 39058
rect 9602 39006 9604 39058
rect 9548 38994 9604 39006
rect 9660 38948 9716 39566
rect 10220 39620 10276 39630
rect 10276 39564 10388 39620
rect 10220 39526 10276 39564
rect 9660 38882 9716 38892
rect 9772 39506 9828 39518
rect 9772 39454 9774 39506
rect 9826 39454 9828 39506
rect 9772 38668 9828 39454
rect 9884 39396 9940 39406
rect 9884 39302 9940 39340
rect 9884 38836 9940 38846
rect 10220 38836 10276 38846
rect 9940 38834 10276 38836
rect 9940 38782 10222 38834
rect 10274 38782 10276 38834
rect 9940 38780 10276 38782
rect 9884 38742 9940 38780
rect 10220 38770 10276 38780
rect 9660 38612 9828 38668
rect 10108 38612 10164 38622
rect 9660 38050 9716 38612
rect 10108 38162 10164 38556
rect 10108 38110 10110 38162
rect 10162 38110 10164 38162
rect 10108 38098 10164 38110
rect 10332 38612 10388 39564
rect 10780 39618 10836 39630
rect 10780 39566 10782 39618
rect 10834 39566 10836 39618
rect 10780 39508 10836 39566
rect 10780 39442 10836 39452
rect 11228 39618 11284 39788
rect 11340 39730 11396 40236
rect 11452 40226 11508 40236
rect 13468 40180 13524 41918
rect 14476 41972 14532 41982
rect 17276 41972 17332 41982
rect 14476 41858 14532 41916
rect 14476 41806 14478 41858
rect 14530 41806 14532 41858
rect 14476 41794 14532 41806
rect 16828 41970 17332 41972
rect 16828 41918 17278 41970
rect 17330 41918 17332 41970
rect 16828 41916 17332 41918
rect 13916 40964 13972 40974
rect 13916 40870 13972 40908
rect 14028 40404 14084 40414
rect 14028 40310 14084 40348
rect 13580 40292 13636 40302
rect 14700 40292 14756 40302
rect 13580 40198 13636 40236
rect 14252 40290 14756 40292
rect 14252 40238 14702 40290
rect 14754 40238 14756 40290
rect 14252 40236 14756 40238
rect 13468 40114 13524 40124
rect 11900 39844 11956 39854
rect 11340 39678 11342 39730
rect 11394 39678 11396 39730
rect 11340 39666 11396 39678
rect 11788 39732 11844 39742
rect 11228 39566 11230 39618
rect 11282 39566 11284 39618
rect 11228 39172 11284 39566
rect 11788 39618 11844 39676
rect 11788 39566 11790 39618
rect 11842 39566 11844 39618
rect 11788 39554 11844 39566
rect 11900 39506 11956 39788
rect 11900 39454 11902 39506
rect 11954 39454 11956 39506
rect 11900 39442 11956 39454
rect 13916 39506 13972 39518
rect 13916 39454 13918 39506
rect 13970 39454 13972 39506
rect 11452 39396 11508 39406
rect 12124 39396 12180 39406
rect 11452 39394 11732 39396
rect 11452 39342 11454 39394
rect 11506 39342 11732 39394
rect 11452 39340 11732 39342
rect 11452 39330 11508 39340
rect 11228 39116 11620 39172
rect 10780 38948 10836 38958
rect 10780 38854 10836 38892
rect 10556 38836 10612 38846
rect 10444 38612 10500 38622
rect 10332 38610 10500 38612
rect 10332 38558 10446 38610
rect 10498 38558 10500 38610
rect 10332 38556 10500 38558
rect 9660 37998 9662 38050
rect 9714 37998 9716 38050
rect 9660 36260 9716 37998
rect 10220 38052 10276 38062
rect 10332 38052 10388 38556
rect 10444 38546 10500 38556
rect 10220 38050 10388 38052
rect 10220 37998 10222 38050
rect 10274 37998 10388 38050
rect 10220 37996 10388 37998
rect 10556 38050 10612 38780
rect 11228 38836 11284 39116
rect 11564 38946 11620 39116
rect 11564 38894 11566 38946
rect 11618 38894 11620 38946
rect 11564 38882 11620 38894
rect 11676 38948 11732 39340
rect 12124 39302 12180 39340
rect 12124 39060 12180 39070
rect 12124 38966 12180 39004
rect 13916 39060 13972 39454
rect 14252 39506 14308 40236
rect 14700 40226 14756 40236
rect 16828 40290 16884 41916
rect 17276 41906 17332 41916
rect 20860 41860 20916 45200
rect 21084 41972 21140 41982
rect 20860 41794 20916 41804
rect 20972 41970 21140 41972
rect 20972 41918 21086 41970
rect 21138 41918 21140 41970
rect 20972 41916 21140 41918
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20076 40460 20356 40516
rect 16828 40238 16830 40290
rect 16882 40238 16884 40290
rect 16828 40226 16884 40238
rect 17052 40404 17108 40414
rect 17612 40404 17668 40414
rect 19740 40404 19796 40414
rect 17052 39730 17108 40348
rect 17052 39678 17054 39730
rect 17106 39678 17108 39730
rect 17052 39666 17108 39678
rect 17500 40348 17612 40404
rect 17500 39618 17556 40348
rect 17612 40310 17668 40348
rect 19628 40348 19740 40404
rect 17500 39566 17502 39618
rect 17554 39566 17556 39618
rect 17500 39554 17556 39566
rect 14252 39454 14254 39506
rect 14306 39454 14308 39506
rect 14252 39442 14308 39454
rect 18172 39506 18228 39518
rect 18172 39454 18174 39506
rect 18226 39454 18228 39506
rect 18172 39284 18228 39454
rect 18172 39218 18228 39228
rect 13916 38994 13972 39004
rect 11676 38836 11732 38892
rect 11788 38836 11844 38846
rect 11676 38834 11844 38836
rect 11676 38782 11790 38834
rect 11842 38782 11844 38834
rect 11676 38780 11844 38782
rect 11228 38770 11284 38780
rect 11788 38770 11844 38780
rect 10556 37998 10558 38050
rect 10610 37998 10612 38050
rect 10220 37716 10276 37996
rect 9660 36194 9716 36204
rect 9996 37660 10276 37716
rect 9772 35476 9828 35486
rect 9996 35476 10052 37660
rect 10444 36258 10500 36270
rect 10444 36206 10446 36258
rect 10498 36206 10500 36258
rect 10332 35586 10388 35598
rect 10332 35534 10334 35586
rect 10386 35534 10388 35586
rect 9772 35474 10052 35476
rect 9772 35422 9774 35474
rect 9826 35422 10052 35474
rect 9772 35420 10052 35422
rect 10108 35474 10164 35486
rect 10108 35422 10110 35474
rect 10162 35422 10164 35474
rect 9772 35410 9828 35420
rect 9884 35028 9940 35038
rect 10108 35028 10164 35422
rect 10332 35476 10388 35534
rect 10332 35410 10388 35420
rect 10444 35252 10500 36206
rect 10556 35924 10612 37998
rect 11452 37938 11508 37950
rect 11452 37886 11454 37938
rect 11506 37886 11508 37938
rect 11452 37828 11508 37886
rect 10668 35924 10724 35934
rect 10556 35922 10724 35924
rect 10556 35870 10670 35922
rect 10722 35870 10724 35922
rect 10556 35868 10724 35870
rect 10668 35858 10724 35868
rect 11116 35812 11172 35822
rect 9884 35026 10164 35028
rect 9884 34974 9886 35026
rect 9938 34974 10164 35026
rect 9884 34972 10164 34974
rect 9884 34962 9940 34972
rect 10108 34916 10164 34972
rect 10108 34850 10164 34860
rect 10220 35028 10276 35038
rect 10220 34914 10276 34972
rect 10220 34862 10222 34914
rect 10274 34862 10276 34914
rect 10220 34850 10276 34862
rect 9772 34692 9828 34702
rect 9996 34692 10052 34702
rect 10108 34692 10164 34702
rect 9772 34690 9940 34692
rect 9772 34638 9774 34690
rect 9826 34638 9940 34690
rect 9772 34636 9940 34638
rect 9772 34626 9828 34636
rect 9436 34524 9716 34580
rect 9660 34468 9716 34524
rect 9660 34412 9828 34468
rect 9548 34356 9604 34366
rect 9212 34300 9492 34356
rect 5180 33954 5236 33964
rect 7084 34132 7140 34142
rect 9436 34132 9492 34300
rect 9604 34300 9716 34356
rect 9548 34290 9604 34300
rect 9660 34242 9716 34300
rect 9660 34190 9662 34242
rect 9714 34190 9716 34242
rect 9660 34178 9716 34190
rect 9548 34132 9604 34142
rect 9436 34130 9604 34132
rect 9436 34078 9550 34130
rect 9602 34078 9604 34130
rect 9436 34076 9604 34078
rect 7084 34018 7140 34076
rect 9548 34066 9604 34076
rect 7084 33966 7086 34018
rect 7138 33966 7140 34018
rect 7084 33954 7140 33966
rect 7532 34020 7588 34030
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 5068 31890 5124 31902
rect 5068 31838 5070 31890
rect 5122 31838 5124 31890
rect 2940 31668 2996 31678
rect 2940 31574 2996 31612
rect 4172 31668 4228 31678
rect 4172 31218 4228 31612
rect 4172 31166 4174 31218
rect 4226 31166 4228 31218
rect 4172 31154 4228 31166
rect 4284 30882 4340 30894
rect 4284 30830 4286 30882
rect 4338 30830 4340 30882
rect 2604 29314 2660 29326
rect 2604 29262 2606 29314
rect 2658 29262 2660 29314
rect 2604 28868 2660 29262
rect 2604 28802 2660 28812
rect 4284 28756 4340 30830
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5068 29540 5124 31838
rect 5740 31556 5796 31566
rect 7532 31556 7588 33964
rect 5796 31500 5908 31556
rect 5740 31462 5796 31500
rect 5852 30996 5908 31500
rect 6076 30996 6132 31006
rect 5852 30994 6132 30996
rect 5852 30942 6078 30994
rect 6130 30942 6132 30994
rect 5852 30940 6132 30942
rect 5852 29650 5908 30940
rect 6076 30930 6132 30940
rect 5852 29598 5854 29650
rect 5906 29598 5908 29650
rect 5852 29586 5908 29598
rect 6860 30882 6916 30894
rect 6860 30830 6862 30882
rect 6914 30830 6916 30882
rect 6860 29652 6916 30830
rect 7532 30884 7588 31500
rect 7532 30818 7588 30828
rect 8988 30882 9044 30894
rect 8988 30830 8990 30882
rect 9042 30830 9044 30882
rect 6860 29586 6916 29596
rect 5068 29484 5684 29540
rect 5628 29428 5684 29484
rect 5628 29372 5908 29428
rect 4844 29314 4900 29326
rect 4844 29262 4846 29314
rect 4898 29262 4900 29314
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4508 28868 4564 28878
rect 4508 28774 4564 28812
rect 4284 28690 4340 28700
rect 4844 28644 4900 29262
rect 4732 28588 4900 28644
rect 5516 29314 5572 29326
rect 5516 29262 5518 29314
rect 5570 29262 5572 29314
rect 4060 28420 4116 28430
rect 4060 26514 4116 28364
rect 4620 28418 4676 28430
rect 4620 28366 4622 28418
rect 4674 28366 4676 28418
rect 4620 28308 4676 28366
rect 4620 27636 4676 28252
rect 4732 28084 4788 28588
rect 5068 28532 5124 28542
rect 5068 28438 5124 28476
rect 4844 28420 4900 28430
rect 4844 28418 5012 28420
rect 4844 28366 4846 28418
rect 4898 28366 5012 28418
rect 4844 28364 5012 28366
rect 4844 28354 4900 28364
rect 4956 28196 5012 28364
rect 5516 28308 5572 29262
rect 5740 28756 5796 28766
rect 5740 28662 5796 28700
rect 5852 28756 5908 29372
rect 6412 28756 6468 28766
rect 5852 28700 6132 28756
rect 5852 28530 5908 28700
rect 5852 28478 5854 28530
rect 5906 28478 5908 28530
rect 5852 28466 5908 28478
rect 5964 28530 6020 28542
rect 5964 28478 5966 28530
rect 6018 28478 6020 28530
rect 5628 28420 5684 28430
rect 5628 28326 5684 28364
rect 5516 28242 5572 28252
rect 4956 28130 5012 28140
rect 5404 28196 5460 28206
rect 4844 28084 4900 28094
rect 4732 28028 4844 28084
rect 4844 28018 4900 28028
rect 5404 28082 5460 28140
rect 5404 28030 5406 28082
rect 5458 28030 5460 28082
rect 5404 28018 5460 28030
rect 5628 28084 5684 28094
rect 5964 28084 6020 28478
rect 5628 27990 5684 28028
rect 5740 28028 6020 28084
rect 5740 27970 5796 28028
rect 5740 27918 5742 27970
rect 5794 27918 5796 27970
rect 5740 27906 5796 27918
rect 4060 26462 4062 26514
rect 4114 26462 4116 26514
rect 4060 26450 4116 26462
rect 4284 27580 4676 27636
rect 4284 26068 4340 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 5964 27186 6020 28028
rect 5964 27134 5966 27186
rect 6018 27134 6020 27186
rect 5964 27122 6020 27134
rect 6076 27076 6132 28700
rect 6412 28642 6468 28700
rect 6972 28756 7028 28766
rect 6972 28662 7028 28700
rect 6412 28590 6414 28642
rect 6466 28590 6468 28642
rect 6412 28578 6468 28590
rect 7756 28532 7812 28542
rect 6076 27020 6468 27076
rect 6412 26908 6468 27020
rect 5852 26852 5908 26862
rect 5852 26850 6020 26852
rect 5852 26798 5854 26850
rect 5906 26798 6020 26850
rect 5852 26796 6020 26798
rect 5852 26786 5908 26796
rect 5292 26516 5348 26526
rect 5292 26402 5348 26460
rect 5292 26350 5294 26402
rect 5346 26350 5348 26402
rect 5292 26338 5348 26350
rect 5852 26404 5908 26414
rect 3836 26012 4284 26068
rect 4508 26290 4564 26302
rect 4508 26238 4510 26290
rect 4562 26238 4564 26290
rect 4508 26068 4564 26238
rect 4620 26292 4676 26302
rect 4620 26198 4676 26236
rect 4844 26292 4900 26302
rect 4844 26290 5012 26292
rect 4844 26238 4846 26290
rect 4898 26238 5012 26290
rect 4844 26236 5012 26238
rect 4844 26226 4900 26236
rect 4956 26180 5012 26236
rect 5404 26290 5460 26302
rect 5404 26238 5406 26290
rect 5458 26238 5460 26290
rect 5404 26180 5460 26238
rect 4956 26124 5460 26180
rect 5516 26290 5572 26302
rect 5516 26238 5518 26290
rect 5570 26238 5572 26290
rect 4508 26012 4900 26068
rect 3612 25620 3668 25630
rect 3836 25620 3892 26012
rect 4284 26002 4340 26012
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4732 25620 4788 25630
rect 3612 25618 3892 25620
rect 3612 25566 3614 25618
rect 3666 25566 3892 25618
rect 3612 25564 3892 25566
rect 3612 25554 3668 25564
rect 3836 25394 3892 25564
rect 4396 25618 4788 25620
rect 4396 25566 4734 25618
rect 4786 25566 4788 25618
rect 4396 25564 4788 25566
rect 4396 25506 4452 25564
rect 4732 25554 4788 25564
rect 4396 25454 4398 25506
rect 4450 25454 4452 25506
rect 4396 25442 4452 25454
rect 4844 25508 4900 26012
rect 4844 25414 4900 25452
rect 3836 25342 3838 25394
rect 3890 25342 3892 25394
rect 3836 25330 3892 25342
rect 4620 25396 4676 25406
rect 4620 25394 4788 25396
rect 4620 25342 4622 25394
rect 4674 25342 4788 25394
rect 4620 25340 4788 25342
rect 4620 25330 4676 25340
rect 3724 25282 3780 25294
rect 3724 25230 3726 25282
rect 3778 25230 3780 25282
rect 2604 23716 2660 23726
rect 2604 22482 2660 23660
rect 3724 23716 3780 25230
rect 4060 25282 4116 25294
rect 4060 25230 4062 25282
rect 4114 25230 4116 25282
rect 4060 24948 4116 25230
rect 4060 24882 4116 24892
rect 4732 24946 4788 25340
rect 4732 24894 4734 24946
rect 4786 24894 4788 24946
rect 4732 24882 4788 24894
rect 4844 25284 4900 25294
rect 4620 24834 4676 24846
rect 4620 24782 4622 24834
rect 4674 24782 4676 24834
rect 4620 24724 4676 24782
rect 4620 24658 4676 24668
rect 4844 24498 4900 25228
rect 4844 24446 4846 24498
rect 4898 24446 4900 24498
rect 4844 24434 4900 24446
rect 4956 24724 5012 26124
rect 5516 25508 5572 26238
rect 5516 25442 5572 25452
rect 5852 25508 5908 26348
rect 5964 26066 6020 26796
rect 6076 26850 6132 26862
rect 6076 26798 6078 26850
rect 6130 26798 6132 26850
rect 6076 26404 6132 26798
rect 6076 26338 6132 26348
rect 6300 26850 6356 26862
rect 6300 26798 6302 26850
rect 6354 26798 6356 26850
rect 5964 26014 5966 26066
rect 6018 26014 6020 26066
rect 5964 25844 6020 26014
rect 6300 26292 6356 26798
rect 6412 26852 6692 26908
rect 6412 26516 6468 26852
rect 6412 26450 6468 26460
rect 6300 25956 6356 26236
rect 6300 25900 6468 25956
rect 5964 25788 6356 25844
rect 5964 25508 6020 25518
rect 5852 25506 6020 25508
rect 5852 25454 5966 25506
rect 6018 25454 6020 25506
rect 5852 25452 6020 25454
rect 5740 25396 5796 25406
rect 5740 25302 5796 25340
rect 5068 25284 5124 25294
rect 5852 25284 5908 25452
rect 5964 25442 6020 25452
rect 6188 25508 6244 25518
rect 6188 25414 6244 25452
rect 5068 25282 5236 25284
rect 5068 25230 5070 25282
rect 5122 25230 5236 25282
rect 5068 25228 5236 25230
rect 5068 25218 5124 25228
rect 5180 25060 5236 25228
rect 5852 25218 5908 25228
rect 6076 25282 6132 25294
rect 6076 25230 6078 25282
rect 6130 25230 6132 25282
rect 5292 25060 5348 25070
rect 5180 25004 5292 25060
rect 5292 24994 5348 25004
rect 5068 24948 5124 24958
rect 5068 24854 5124 24892
rect 5852 24948 5908 24958
rect 5852 24854 5908 24892
rect 5292 24834 5348 24846
rect 5292 24782 5294 24834
rect 5346 24782 5348 24834
rect 5292 24724 5348 24782
rect 5012 24668 5348 24724
rect 5404 24724 5460 24734
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 3724 23650 3780 23660
rect 2604 22430 2606 22482
rect 2658 22430 2660 22482
rect 2604 22418 2660 22430
rect 3164 23604 3220 23614
rect 2268 22082 2324 22092
rect 3164 20130 3220 23548
rect 4956 23378 5012 24668
rect 5404 24630 5460 24668
rect 6076 24724 6132 25230
rect 6076 23828 6132 24668
rect 6188 25284 6244 25294
rect 6188 23938 6244 25228
rect 6300 24836 6356 25788
rect 6412 25396 6468 25900
rect 6412 25330 6468 25340
rect 6300 24770 6356 24780
rect 6188 23886 6190 23938
rect 6242 23886 6244 23938
rect 6188 23874 6244 23886
rect 6076 23762 6132 23772
rect 6524 23826 6580 23838
rect 6524 23774 6526 23826
rect 6578 23774 6580 23826
rect 6300 23716 6356 23726
rect 6300 23622 6356 23660
rect 4956 23326 4958 23378
rect 5010 23326 5012 23378
rect 4956 23314 5012 23326
rect 6524 23492 6580 23774
rect 5292 23154 5348 23166
rect 5292 23102 5294 23154
rect 5346 23102 5348 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4732 22482 4788 22494
rect 4732 22430 4734 22482
rect 4786 22430 4788 22482
rect 4732 22372 4788 22430
rect 4732 22306 4788 22316
rect 5292 22372 5348 23102
rect 5292 22306 5348 22316
rect 5516 22260 5572 22270
rect 5740 22260 5796 22270
rect 5572 22258 6020 22260
rect 5572 22206 5742 22258
rect 5794 22206 6020 22258
rect 5572 22204 6020 22206
rect 5516 22194 5572 22204
rect 5740 22194 5796 22204
rect 5404 21476 5460 21486
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 5404 20242 5460 21420
rect 5404 20190 5406 20242
rect 5458 20190 5460 20242
rect 5404 20178 5460 20190
rect 3164 20078 3166 20130
rect 3218 20078 3220 20130
rect 3164 20066 3220 20078
rect 5964 20130 6020 22204
rect 6412 21586 6468 21598
rect 6412 21534 6414 21586
rect 6466 21534 6468 21586
rect 6412 21476 6468 21534
rect 6412 21410 6468 21420
rect 6524 21474 6580 23436
rect 6636 21588 6692 26852
rect 7196 25508 7252 25518
rect 7196 25414 7252 25452
rect 7644 24836 7700 24846
rect 7644 24742 7700 24780
rect 7756 24498 7812 28476
rect 8764 27188 8820 27198
rect 8316 25620 8372 25630
rect 8316 25526 8372 25564
rect 7980 25506 8036 25518
rect 7980 25454 7982 25506
rect 8034 25454 8036 25506
rect 7868 24948 7924 24958
rect 7868 24854 7924 24892
rect 7756 24446 7758 24498
rect 7810 24446 7812 24498
rect 7756 24434 7812 24446
rect 7196 24162 7252 24174
rect 7196 24110 7198 24162
rect 7250 24110 7252 24162
rect 7196 24052 7252 24110
rect 7756 24164 7812 24174
rect 7756 24052 7812 24108
rect 6972 23996 7252 24052
rect 7308 24050 7812 24052
rect 7308 23998 7758 24050
rect 7810 23998 7812 24050
rect 7308 23996 7812 23998
rect 6748 23940 6804 23950
rect 6972 23940 7028 23996
rect 6748 23938 7028 23940
rect 6748 23886 6750 23938
rect 6802 23886 7028 23938
rect 6748 23884 7028 23886
rect 6748 23874 6804 23884
rect 7084 23828 7140 23838
rect 7084 23734 7140 23772
rect 7196 23828 7252 23838
rect 7308 23828 7364 23996
rect 7196 23826 7364 23828
rect 7196 23774 7198 23826
rect 7250 23774 7364 23826
rect 7196 23772 7364 23774
rect 7196 23762 7252 23772
rect 7084 22372 7140 22382
rect 6748 21588 6804 21598
rect 6636 21532 6748 21588
rect 6748 21522 6804 21532
rect 6524 21422 6526 21474
rect 6578 21422 6580 21474
rect 6524 21410 6580 21422
rect 5964 20078 5966 20130
rect 6018 20078 6020 20130
rect 5964 20066 6020 20078
rect 2380 20020 2436 20030
rect 1932 20018 2436 20020
rect 1932 19966 2382 20018
rect 2434 19966 2436 20018
rect 1932 19964 2436 19966
rect 1932 16884 1988 19964
rect 2380 19954 2436 19964
rect 7084 20018 7140 22316
rect 7644 22372 7700 22382
rect 7532 21812 7588 21822
rect 7644 21812 7700 22316
rect 7756 21924 7812 23996
rect 7980 23492 8036 25454
rect 8204 25508 8260 25518
rect 8204 25414 8260 25452
rect 8764 24948 8820 27132
rect 8988 27076 9044 30830
rect 9660 30884 9716 30894
rect 9660 30790 9716 30828
rect 9548 30322 9604 30334
rect 9548 30270 9550 30322
rect 9602 30270 9604 30322
rect 9548 28644 9604 30270
rect 9548 28578 9604 28588
rect 9772 28084 9828 34412
rect 9884 34132 9940 34636
rect 9996 34690 10108 34692
rect 9996 34638 9998 34690
rect 10050 34638 10108 34690
rect 9996 34636 10108 34638
rect 9996 34626 10052 34636
rect 10108 34354 10164 34636
rect 10444 34580 10500 35196
rect 10780 35810 11172 35812
rect 10780 35758 11118 35810
rect 11170 35758 11172 35810
rect 10780 35756 11172 35758
rect 10780 35026 10836 35756
rect 11116 35746 11172 35756
rect 11228 35812 11284 35822
rect 11228 35718 11284 35756
rect 11340 35698 11396 35710
rect 11340 35646 11342 35698
rect 11394 35646 11396 35698
rect 11340 35588 11396 35646
rect 11116 35532 11396 35588
rect 11116 35252 11172 35532
rect 11452 35476 11508 37772
rect 12124 37828 12180 37838
rect 12124 37734 12180 37772
rect 19628 37492 19684 40348
rect 19740 40338 19796 40348
rect 20076 40404 20132 40460
rect 20076 40310 20132 40348
rect 20300 40402 20356 40460
rect 20300 40350 20302 40402
rect 20354 40350 20356 40402
rect 20300 40338 20356 40350
rect 20972 39956 21028 41916
rect 21084 41906 21140 41916
rect 23212 41972 23268 41982
rect 22092 41860 22148 41870
rect 22092 41766 22148 41804
rect 20300 39900 21028 39956
rect 21084 40290 21140 40302
rect 21084 40238 21086 40290
rect 21138 40238 21140 40290
rect 20300 39730 20356 39900
rect 20300 39678 20302 39730
rect 20354 39678 20356 39730
rect 20300 39666 20356 39678
rect 21084 39508 21140 40238
rect 23212 40290 23268 41916
rect 24668 41860 24724 45200
rect 24668 41794 24724 41804
rect 24892 41970 24948 41982
rect 24892 41918 24894 41970
rect 24946 41918 24948 41970
rect 23212 40238 23214 40290
rect 23266 40238 23268 40290
rect 23212 40226 23268 40238
rect 24892 40292 24948 41918
rect 25900 41860 25956 41870
rect 25900 41766 25956 41804
rect 28476 41860 28532 45200
rect 32284 45108 32340 45200
rect 32620 45108 32676 45276
rect 32284 45052 32676 45108
rect 33068 43708 33124 45276
rect 36064 45200 36176 46000
rect 39872 45200 39984 46000
rect 43680 45200 43792 46000
rect 33068 43652 33572 43708
rect 33516 42194 33572 43652
rect 33516 42142 33518 42194
rect 33570 42142 33572 42194
rect 33516 42130 33572 42142
rect 28700 41972 28756 41982
rect 28700 41878 28756 41916
rect 31388 41972 31444 41982
rect 28476 41794 28532 41804
rect 29708 41860 29764 41870
rect 29708 41766 29764 41804
rect 28476 40962 28532 40974
rect 28476 40910 28478 40962
rect 28530 40910 28532 40962
rect 25340 40404 25396 40414
rect 25340 40310 25396 40348
rect 28476 40404 28532 40910
rect 26012 40292 26068 40302
rect 24892 40226 24948 40236
rect 25900 40290 26068 40292
rect 25900 40238 26014 40290
rect 26066 40238 26068 40290
rect 25900 40236 26068 40238
rect 21084 39442 21140 39452
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 25564 38050 25620 38062
rect 25564 37998 25566 38050
rect 25618 37998 25620 38050
rect 21868 37940 21924 37950
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19740 37492 19796 37502
rect 19516 37490 20132 37492
rect 19516 37438 19742 37490
rect 19794 37438 20132 37490
rect 19516 37436 20132 37438
rect 17276 36484 17332 36494
rect 17276 36390 17332 36428
rect 17500 36482 17556 36494
rect 17500 36430 17502 36482
rect 17554 36430 17556 36482
rect 15596 36372 15652 36382
rect 15484 36260 15540 36270
rect 15260 36258 15540 36260
rect 15260 36206 15486 36258
rect 15538 36206 15540 36258
rect 15260 36204 15540 36206
rect 14700 35810 14756 35822
rect 14700 35758 14702 35810
rect 14754 35758 14756 35810
rect 11116 35186 11172 35196
rect 11228 35420 11508 35476
rect 11564 35476 11620 35486
rect 10780 34974 10782 35026
rect 10834 34974 10836 35026
rect 10780 34962 10836 34974
rect 11116 34916 11172 34926
rect 11116 34822 11172 34860
rect 10444 34514 10500 34524
rect 10668 34690 10724 34702
rect 10668 34638 10670 34690
rect 10722 34638 10724 34690
rect 10108 34302 10110 34354
rect 10162 34302 10164 34354
rect 10108 34290 10164 34302
rect 10556 34356 10612 34366
rect 9884 34076 10164 34132
rect 10108 33572 10164 34076
rect 10556 34130 10612 34300
rect 10556 34078 10558 34130
rect 10610 34078 10612 34130
rect 10556 34066 10612 34078
rect 10220 33572 10276 33582
rect 10108 33516 10220 33572
rect 10220 33458 10276 33516
rect 10668 33572 10724 34638
rect 10892 34692 10948 34702
rect 10892 34598 10948 34636
rect 10892 34020 10948 34030
rect 11228 34020 11284 35420
rect 11340 35028 11396 35038
rect 11340 34934 11396 34972
rect 11564 34914 11620 35420
rect 14588 35476 14644 35486
rect 14700 35476 14756 35758
rect 14924 35700 14980 35710
rect 14924 35698 15092 35700
rect 14924 35646 14926 35698
rect 14978 35646 15092 35698
rect 14924 35644 15092 35646
rect 14924 35634 14980 35644
rect 14924 35476 14980 35486
rect 14700 35420 14924 35476
rect 14588 35382 14644 35420
rect 14924 35410 14980 35420
rect 14140 35252 14196 35262
rect 11564 34862 11566 34914
rect 11618 34862 11620 34914
rect 11564 34850 11620 34862
rect 11676 34914 11732 34926
rect 11676 34862 11678 34914
rect 11730 34862 11732 34914
rect 10668 33506 10724 33516
rect 10780 34018 11284 34020
rect 10780 33966 10894 34018
rect 10946 33966 11284 34018
rect 10780 33964 11284 33966
rect 11340 34356 11396 34366
rect 10220 33406 10222 33458
rect 10274 33406 10276 33458
rect 10220 33394 10276 33406
rect 10332 28644 10388 28654
rect 8988 27010 9044 27020
rect 9660 28028 9828 28084
rect 9996 28084 10052 28094
rect 9548 26178 9604 26190
rect 9548 26126 9550 26178
rect 9602 26126 9604 26178
rect 8764 24854 8820 24892
rect 9212 25732 9268 25742
rect 8092 24722 8148 24734
rect 8092 24670 8094 24722
rect 8146 24670 8148 24722
rect 8092 24276 8148 24670
rect 8316 24722 8372 24734
rect 8316 24670 8318 24722
rect 8370 24670 8372 24722
rect 8316 24500 8372 24670
rect 8316 24434 8372 24444
rect 8092 24210 8148 24220
rect 7868 23436 7980 23492
rect 7868 22258 7924 23436
rect 7980 23426 8036 23436
rect 8764 23604 8820 23614
rect 8652 22372 8708 22382
rect 8652 22278 8708 22316
rect 7868 22206 7870 22258
rect 7922 22206 7924 22258
rect 7868 22194 7924 22206
rect 8764 22258 8820 23548
rect 8764 22206 8766 22258
rect 8818 22206 8820 22258
rect 8764 22194 8820 22206
rect 9100 23268 9156 23278
rect 7756 21868 7924 21924
rect 7532 21810 7812 21812
rect 7532 21758 7534 21810
rect 7586 21758 7812 21810
rect 7532 21756 7812 21758
rect 7532 21746 7588 21756
rect 7420 21588 7476 21598
rect 7420 20692 7476 21532
rect 7420 20626 7476 20636
rect 7756 20690 7812 21756
rect 7756 20638 7758 20690
rect 7810 20638 7812 20690
rect 7756 20626 7812 20638
rect 7756 20132 7812 20142
rect 7756 20038 7812 20076
rect 7084 19966 7086 20018
rect 7138 19966 7140 20018
rect 7084 19954 7140 19966
rect 7532 20018 7588 20030
rect 7532 19966 7534 20018
rect 7586 19966 7588 20018
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 6972 18340 7028 18350
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 6972 17106 7028 18284
rect 6972 17054 6974 17106
rect 7026 17054 7028 17106
rect 4396 16996 4452 17006
rect 4396 16902 4452 16940
rect 1932 16098 1988 16828
rect 3612 16884 3668 16894
rect 3612 16790 3668 16828
rect 4844 16884 4900 16894
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 2604 16212 2660 16222
rect 2604 16118 2660 16156
rect 4732 16212 4788 16222
rect 4844 16212 4900 16828
rect 6524 16772 6580 16782
rect 6524 16678 6580 16716
rect 4732 16210 4900 16212
rect 4732 16158 4734 16210
rect 4786 16158 4900 16210
rect 4732 16156 4900 16158
rect 5740 16212 5796 16222
rect 4732 16146 4788 16156
rect 5740 16118 5796 16156
rect 6972 16212 7028 17054
rect 1932 16046 1934 16098
rect 1986 16046 1988 16098
rect 1932 11956 1988 16046
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4172 13636 4228 13646
rect 4172 12290 4228 13580
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 6412 12404 6468 12414
rect 6412 12310 6468 12348
rect 4172 12238 4174 12290
rect 4226 12238 4228 12290
rect 4172 12226 4228 12238
rect 4844 12292 4900 12302
rect 1932 11394 1988 11900
rect 3500 12178 3556 12190
rect 3500 12126 3502 12178
rect 3554 12126 3556 12178
rect 3500 11956 3556 12126
rect 3500 11890 3556 11900
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11506 4900 12236
rect 6972 12066 7028 16156
rect 6972 12014 6974 12066
rect 7026 12014 7028 12066
rect 4844 11454 4846 11506
rect 4898 11454 4900 11506
rect 4844 11442 4900 11454
rect 5740 11956 5796 11966
rect 5740 11508 5796 11900
rect 5740 11414 5796 11452
rect 6972 11508 7028 12014
rect 1932 11342 1934 11394
rect 1986 11342 1988 11394
rect 1932 11330 1988 11342
rect 2604 11396 2660 11406
rect 2604 11302 2660 11340
rect 6972 10388 7028 11452
rect 6972 10322 7028 10332
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 7532 9826 7588 19966
rect 7868 10612 7924 21868
rect 8316 21700 8372 21710
rect 8316 20914 8372 21644
rect 8316 20862 8318 20914
rect 8370 20862 8372 20914
rect 8316 20850 8372 20862
rect 8204 20802 8260 20814
rect 8204 20750 8206 20802
rect 8258 20750 8260 20802
rect 8204 18564 8260 20750
rect 9100 20802 9156 23212
rect 9100 20750 9102 20802
rect 9154 20750 9156 20802
rect 9100 20738 9156 20750
rect 8988 20578 9044 20590
rect 8988 20526 8990 20578
rect 9042 20526 9044 20578
rect 8204 18498 8260 18508
rect 8316 19234 8372 19246
rect 8316 19182 8318 19234
rect 8370 19182 8372 19234
rect 8316 18004 8372 19182
rect 8316 17948 8932 18004
rect 8876 17890 8932 17948
rect 8876 17838 8878 17890
rect 8930 17838 8932 17890
rect 8876 15876 8932 17838
rect 8988 17556 9044 20526
rect 9100 19236 9156 19246
rect 9212 19236 9268 25676
rect 9548 25508 9604 26126
rect 9548 23268 9604 25452
rect 9660 25060 9716 28028
rect 9884 27076 9940 27086
rect 9884 26402 9940 27020
rect 9884 26350 9886 26402
rect 9938 26350 9940 26402
rect 9884 26338 9940 26350
rect 9660 24994 9716 25004
rect 9996 24836 10052 28028
rect 10108 24836 10164 24846
rect 9996 24834 10164 24836
rect 9996 24782 10110 24834
rect 10162 24782 10164 24834
rect 9996 24780 10164 24782
rect 9996 23604 10052 24780
rect 10108 24770 10164 24780
rect 9548 23202 9604 23212
rect 9884 23548 9996 23604
rect 10220 24500 10276 24510
rect 10220 23604 10276 24444
rect 10332 23828 10388 28588
rect 10444 27074 10500 27086
rect 10444 27022 10446 27074
rect 10498 27022 10500 27074
rect 10444 25732 10500 27022
rect 10780 26908 10836 33964
rect 10892 33954 10948 33964
rect 11340 33346 11396 34300
rect 11676 34356 11732 34862
rect 12348 34692 12404 34702
rect 12348 34598 12404 34636
rect 14140 34690 14196 35196
rect 14700 35028 14756 35038
rect 15036 35028 15092 35644
rect 15260 35698 15316 36204
rect 15484 36194 15540 36204
rect 15260 35646 15262 35698
rect 15314 35646 15316 35698
rect 15260 35634 15316 35646
rect 15596 35700 15652 36316
rect 16940 36372 16996 36382
rect 16940 36278 16996 36316
rect 16156 36260 16212 36270
rect 16044 36204 16156 36260
rect 15708 35700 15764 35710
rect 15596 35698 15764 35700
rect 15596 35646 15710 35698
rect 15762 35646 15764 35698
rect 15596 35644 15764 35646
rect 15708 35634 15764 35644
rect 15708 35476 15764 35486
rect 15596 35028 15652 35038
rect 15036 34972 15428 35028
rect 14700 34914 14756 34972
rect 14700 34862 14702 34914
rect 14754 34862 14756 34914
rect 14700 34850 14756 34862
rect 15372 34916 15428 34972
rect 15596 34934 15652 34972
rect 15372 34822 15428 34860
rect 14364 34804 14420 34814
rect 14924 34804 14980 34814
rect 14364 34710 14420 34748
rect 14812 34802 14980 34804
rect 14812 34750 14926 34802
rect 14978 34750 14980 34802
rect 14812 34748 14980 34750
rect 14140 34638 14142 34690
rect 14194 34638 14196 34690
rect 14140 34580 14196 34638
rect 14476 34690 14532 34702
rect 14476 34638 14478 34690
rect 14530 34638 14532 34690
rect 14476 34580 14532 34638
rect 14140 34524 14532 34580
rect 11676 34290 11732 34300
rect 14140 34132 14196 34142
rect 14140 34038 14196 34076
rect 11452 34018 11508 34030
rect 11452 33966 11454 34018
rect 11506 33966 11508 34018
rect 11452 33572 11508 33966
rect 14364 33908 14420 33918
rect 14364 33814 14420 33852
rect 11452 33506 11508 33516
rect 11340 33294 11342 33346
rect 11394 33294 11396 33346
rect 11340 33282 11396 33294
rect 11676 33124 11732 33134
rect 11676 33030 11732 33068
rect 12908 33124 12964 33134
rect 12908 31780 12964 33068
rect 12908 31686 12964 31724
rect 13580 31780 13636 31790
rect 13580 31686 13636 31724
rect 14028 31778 14084 31790
rect 14028 31726 14030 31778
rect 14082 31726 14084 31778
rect 13020 31668 13076 31678
rect 10892 30884 10948 30894
rect 10892 30790 10948 30828
rect 12460 30212 12516 30222
rect 13020 30212 13076 31612
rect 12460 30210 13076 30212
rect 12460 30158 12462 30210
rect 12514 30158 13022 30210
rect 13074 30158 13076 30210
rect 12460 30156 13076 30158
rect 12460 30146 12516 30156
rect 13020 30146 13076 30156
rect 14028 31556 14084 31726
rect 11676 30098 11732 30110
rect 11676 30046 11678 30098
rect 11730 30046 11732 30098
rect 11228 29652 11284 29662
rect 11228 29558 11284 29596
rect 11452 29652 11508 29662
rect 11452 29426 11508 29596
rect 11452 29374 11454 29426
rect 11506 29374 11508 29426
rect 11452 29362 11508 29374
rect 11116 29204 11172 29214
rect 11116 29202 11396 29204
rect 11116 29150 11118 29202
rect 11170 29150 11396 29202
rect 11116 29148 11396 29150
rect 11116 29138 11172 29148
rect 10892 27188 10948 27198
rect 10892 27074 10948 27132
rect 11340 27186 11396 29148
rect 11676 28756 11732 30046
rect 11900 29652 11956 29662
rect 11900 29558 11956 29596
rect 14028 29652 14084 31500
rect 14028 29586 14084 29596
rect 14364 30324 14420 30334
rect 14364 29426 14420 30268
rect 14364 29374 14366 29426
rect 14418 29374 14420 29426
rect 14364 29362 14420 29374
rect 13916 29202 13972 29214
rect 13916 29150 13918 29202
rect 13970 29150 13972 29202
rect 11676 28690 11732 28700
rect 12572 28756 12628 28766
rect 11452 28644 11508 28654
rect 11564 28644 11620 28654
rect 11508 28642 11620 28644
rect 11508 28590 11566 28642
rect 11618 28590 11620 28642
rect 11508 28588 11620 28590
rect 11452 28082 11508 28588
rect 11564 28578 11620 28588
rect 11900 28642 11956 28654
rect 11900 28590 11902 28642
rect 11954 28590 11956 28642
rect 11900 28420 11956 28590
rect 11900 28354 11956 28364
rect 12348 28642 12404 28654
rect 12348 28590 12350 28642
rect 12402 28590 12404 28642
rect 11452 28030 11454 28082
rect 11506 28030 11508 28082
rect 11452 28018 11508 28030
rect 12348 28082 12404 28590
rect 12348 28030 12350 28082
rect 12402 28030 12404 28082
rect 12348 28018 12404 28030
rect 12460 28642 12516 28654
rect 12460 28590 12462 28642
rect 12514 28590 12516 28642
rect 12460 28420 12516 28590
rect 12572 28644 12628 28700
rect 12796 28756 12852 28766
rect 12684 28644 12740 28654
rect 12572 28642 12740 28644
rect 12572 28590 12686 28642
rect 12738 28590 12740 28642
rect 12572 28588 12740 28590
rect 12684 28578 12740 28588
rect 11900 27972 11956 27982
rect 11900 27878 11956 27916
rect 11676 27860 11732 27870
rect 11340 27134 11342 27186
rect 11394 27134 11396 27186
rect 11340 27122 11396 27134
rect 11452 27746 11508 27758
rect 11452 27694 11454 27746
rect 11506 27694 11508 27746
rect 10892 27022 10894 27074
rect 10946 27022 10948 27074
rect 10892 27010 10948 27022
rect 10780 26852 10948 26908
rect 10780 26404 10836 26414
rect 10444 25666 10500 25676
rect 10556 26292 10612 26302
rect 10556 25620 10612 26236
rect 10780 26290 10836 26348
rect 10780 26238 10782 26290
rect 10834 26238 10836 26290
rect 10780 26226 10836 26238
rect 10556 25554 10612 25564
rect 10780 25732 10836 25742
rect 10780 25394 10836 25676
rect 10780 25342 10782 25394
rect 10834 25342 10836 25394
rect 10780 25330 10836 25342
rect 10668 25284 10724 25294
rect 10668 25190 10724 25228
rect 10556 25060 10612 25070
rect 10556 24834 10612 25004
rect 10556 24782 10558 24834
rect 10610 24782 10612 24834
rect 10556 24770 10612 24782
rect 10668 24498 10724 24510
rect 10668 24446 10670 24498
rect 10722 24446 10724 24498
rect 10668 24276 10724 24446
rect 10668 24210 10724 24220
rect 10332 23772 10612 23828
rect 10220 23548 10500 23604
rect 9884 20690 9940 23548
rect 9996 23538 10052 23548
rect 9996 22484 10052 22494
rect 9996 22390 10052 22428
rect 10444 21698 10500 23548
rect 10444 21646 10446 21698
rect 10498 21646 10500 21698
rect 10444 21634 10500 21646
rect 9884 20638 9886 20690
rect 9938 20638 9940 20690
rect 9884 20626 9940 20638
rect 9996 20802 10052 20814
rect 9996 20750 9998 20802
rect 10050 20750 10052 20802
rect 9100 19234 9268 19236
rect 9100 19182 9102 19234
rect 9154 19182 9268 19234
rect 9100 19180 9268 19182
rect 9436 20132 9492 20142
rect 9436 19234 9492 20076
rect 9996 20132 10052 20750
rect 10556 20802 10612 23772
rect 10556 20750 10558 20802
rect 10610 20750 10612 20802
rect 10556 20738 10612 20750
rect 10780 21586 10836 21598
rect 10780 21534 10782 21586
rect 10834 21534 10836 21586
rect 9996 20066 10052 20076
rect 10556 20578 10612 20590
rect 10556 20526 10558 20578
rect 10610 20526 10612 20578
rect 10556 20020 10612 20526
rect 10556 19954 10612 19964
rect 10668 20578 10724 20590
rect 10668 20526 10670 20578
rect 10722 20526 10724 20578
rect 9996 19908 10052 19918
rect 9436 19182 9438 19234
rect 9490 19182 9492 19234
rect 9100 19170 9156 19180
rect 9436 19170 9492 19182
rect 9884 19906 10052 19908
rect 9884 19854 9998 19906
rect 10050 19854 10052 19906
rect 9884 19852 10052 19854
rect 8988 16772 9044 17500
rect 9436 18900 9492 18910
rect 9212 17444 9268 17454
rect 9212 17442 9380 17444
rect 9212 17390 9214 17442
rect 9266 17390 9380 17442
rect 9212 17388 9380 17390
rect 9212 17378 9268 17388
rect 8988 16706 9044 16716
rect 9100 16996 9156 17006
rect 8988 16212 9044 16222
rect 8988 16098 9044 16156
rect 9100 16210 9156 16940
rect 9100 16158 9102 16210
rect 9154 16158 9156 16210
rect 9100 16146 9156 16158
rect 8988 16046 8990 16098
rect 9042 16046 9044 16098
rect 8988 16034 9044 16046
rect 9212 15986 9268 15998
rect 9212 15934 9214 15986
rect 9266 15934 9268 15986
rect 9212 15876 9268 15934
rect 8876 15820 9268 15876
rect 9324 14532 9380 17388
rect 9436 16100 9492 18844
rect 9660 18788 9716 18798
rect 9660 17666 9716 18732
rect 9660 17614 9662 17666
rect 9714 17614 9716 17666
rect 9660 17602 9716 17614
rect 9884 18452 9940 19852
rect 9996 19842 10052 19852
rect 10108 19796 10164 19806
rect 10108 19702 10164 19740
rect 10668 19236 10724 20526
rect 10780 20244 10836 21534
rect 10892 20580 10948 26852
rect 11116 26850 11172 26862
rect 11116 26798 11118 26850
rect 11170 26798 11172 26850
rect 11116 26402 11172 26798
rect 11116 26350 11118 26402
rect 11170 26350 11172 26402
rect 11116 26338 11172 26350
rect 11340 26850 11396 26862
rect 11340 26798 11342 26850
rect 11394 26798 11396 26850
rect 11004 26068 11060 26078
rect 11340 26068 11396 26798
rect 11452 26292 11508 27694
rect 11564 27074 11620 27086
rect 11564 27022 11566 27074
rect 11618 27022 11620 27074
rect 11564 26964 11620 27022
rect 11564 26898 11620 26908
rect 11452 26226 11508 26236
rect 11004 26066 11396 26068
rect 11004 26014 11006 26066
rect 11058 26014 11396 26066
rect 11004 26012 11396 26014
rect 11004 25732 11060 26012
rect 11004 25666 11060 25676
rect 11340 25732 11396 25742
rect 11340 25506 11396 25676
rect 11340 25454 11342 25506
rect 11394 25454 11396 25506
rect 11340 25442 11396 25454
rect 11004 25396 11060 25406
rect 11004 25302 11060 25340
rect 11116 25060 11172 25070
rect 11116 24946 11172 25004
rect 11116 24894 11118 24946
rect 11170 24894 11172 24946
rect 11116 24882 11172 24894
rect 11676 23044 11732 27804
rect 12124 27188 12180 27198
rect 12124 27094 12180 27132
rect 12460 27076 12516 28364
rect 12572 28084 12628 28094
rect 12796 28084 12852 28700
rect 12908 28644 12964 28654
rect 12908 28550 12964 28588
rect 12572 28082 13188 28084
rect 12572 28030 12574 28082
rect 12626 28030 13188 28082
rect 12572 28028 13188 28030
rect 12572 28018 12628 28028
rect 12684 27858 12740 27870
rect 12684 27806 12686 27858
rect 12738 27806 12740 27858
rect 12572 27076 12628 27086
rect 12460 27020 12572 27076
rect 12572 27010 12628 27020
rect 12684 26964 12740 27806
rect 13132 27748 13188 28028
rect 13132 27746 13300 27748
rect 13132 27694 13134 27746
rect 13186 27694 13300 27746
rect 13132 27692 13300 27694
rect 13132 27682 13188 27692
rect 12684 26852 13076 26908
rect 12236 26516 12292 26526
rect 12236 26422 12292 26460
rect 13020 26514 13076 26852
rect 13020 26462 13022 26514
rect 13074 26462 13076 26514
rect 13020 26450 13076 26462
rect 13132 26516 13188 26526
rect 13132 26422 13188 26460
rect 11900 26404 11956 26414
rect 11900 26310 11956 26348
rect 12908 26290 12964 26302
rect 12908 26238 12910 26290
rect 12962 26238 12964 26290
rect 12908 25732 12964 26238
rect 12908 25666 12964 25676
rect 13244 24612 13300 27692
rect 13916 26908 13972 29150
rect 14140 27076 14196 27086
rect 13916 26852 14084 26908
rect 13580 26292 13636 26302
rect 13580 26198 13636 26236
rect 13580 25732 13636 25742
rect 13580 25638 13636 25676
rect 14028 25620 14084 26852
rect 14028 25554 14084 25564
rect 13244 24546 13300 24556
rect 14140 25506 14196 27020
rect 14476 26852 14532 34524
rect 14700 34356 14756 34366
rect 14812 34356 14868 34748
rect 14924 34738 14980 34748
rect 14700 34354 14868 34356
rect 14700 34302 14702 34354
rect 14754 34302 14868 34354
rect 14700 34300 14868 34302
rect 15372 34692 15428 34702
rect 14700 34290 14756 34300
rect 15260 33908 15316 33918
rect 15260 32564 15316 33852
rect 15260 32470 15316 32508
rect 15148 31668 15204 31678
rect 15148 31574 15204 31612
rect 14924 30324 14980 30334
rect 14924 30210 14980 30268
rect 14924 30158 14926 30210
rect 14978 30158 14980 30210
rect 14924 30146 14980 30158
rect 15148 29988 15204 29998
rect 15148 29986 15316 29988
rect 15148 29934 15150 29986
rect 15202 29934 15316 29986
rect 15148 29932 15316 29934
rect 15148 29922 15204 29932
rect 15148 28754 15204 28766
rect 15148 28702 15150 28754
rect 15202 28702 15204 28754
rect 15148 28644 15204 28702
rect 15148 28578 15204 28588
rect 15148 28418 15204 28430
rect 15148 28366 15150 28418
rect 15202 28366 15204 28418
rect 15148 27860 15204 28366
rect 15260 28420 15316 29932
rect 15372 28644 15428 34636
rect 15708 34690 15764 35420
rect 15932 35474 15988 35486
rect 15932 35422 15934 35474
rect 15986 35422 15988 35474
rect 15932 35140 15988 35422
rect 15932 35074 15988 35084
rect 15932 34804 15988 34814
rect 16044 34804 16100 36204
rect 16156 36194 16212 36204
rect 17500 36148 17556 36430
rect 19068 36484 19124 36494
rect 18060 36370 18116 36382
rect 18060 36318 18062 36370
rect 18114 36318 18116 36370
rect 17724 36260 17780 36270
rect 17724 36166 17780 36204
rect 17948 36258 18004 36270
rect 17948 36206 17950 36258
rect 18002 36206 18004 36258
rect 17500 36082 17556 36092
rect 17948 35924 18004 36206
rect 18060 36148 18116 36318
rect 18060 36082 18116 36092
rect 17612 35868 18004 35924
rect 16268 35812 16324 35822
rect 16268 35586 16324 35756
rect 16380 35700 16436 35738
rect 16380 35634 16436 35644
rect 17388 35700 17444 35710
rect 17388 35606 17444 35644
rect 16268 35534 16270 35586
rect 16322 35534 16324 35586
rect 16268 35522 16324 35534
rect 16492 35476 16548 35486
rect 16492 35382 16548 35420
rect 17164 35476 17220 35486
rect 17164 35138 17220 35420
rect 17164 35086 17166 35138
rect 17218 35086 17220 35138
rect 17164 35074 17220 35086
rect 16828 35026 16884 35038
rect 16828 34974 16830 35026
rect 16882 34974 16884 35026
rect 16828 34916 16884 34974
rect 16828 34850 16884 34860
rect 15932 34802 16100 34804
rect 15932 34750 15934 34802
rect 15986 34750 16100 34802
rect 15932 34748 16100 34750
rect 17388 34802 17444 34814
rect 17388 34750 17390 34802
rect 17442 34750 17444 34802
rect 15932 34738 15988 34748
rect 15708 34638 15710 34690
rect 15762 34638 15764 34690
rect 15484 32676 15540 32686
rect 15708 32676 15764 34638
rect 17388 34692 17444 34750
rect 17612 34692 17668 35868
rect 17948 35810 18004 35868
rect 19068 35922 19124 36428
rect 19068 35870 19070 35922
rect 19122 35870 19124 35922
rect 19068 35858 19124 35870
rect 17948 35758 17950 35810
rect 18002 35758 18004 35810
rect 17948 35746 18004 35758
rect 18172 35812 18228 35822
rect 17836 35700 17892 35710
rect 17836 35476 17892 35644
rect 18172 35698 18228 35756
rect 18620 35812 18676 35822
rect 18620 35718 18676 35756
rect 18172 35646 18174 35698
rect 18226 35646 18228 35698
rect 18172 35634 18228 35646
rect 18732 35700 18788 35710
rect 18732 35606 18788 35644
rect 19180 35700 19236 35710
rect 19180 35606 19236 35644
rect 18620 35476 18676 35486
rect 17836 35420 18116 35476
rect 17724 35140 17780 35150
rect 17724 35046 17780 35084
rect 18060 35138 18116 35420
rect 18620 35382 18676 35420
rect 18060 35086 18062 35138
rect 18114 35086 18116 35138
rect 18060 35074 18116 35086
rect 17836 34692 17892 34702
rect 17388 34690 17892 34692
rect 17388 34638 17838 34690
rect 17890 34638 17892 34690
rect 17388 34636 17892 34638
rect 15484 32674 15764 32676
rect 15484 32622 15486 32674
rect 15538 32622 15764 32674
rect 15484 32620 15764 32622
rect 17052 33572 17108 33582
rect 15484 31948 15540 32620
rect 16940 32564 16996 32574
rect 15484 31892 16324 31948
rect 16268 31218 16324 31892
rect 16268 31166 16270 31218
rect 16322 31166 16324 31218
rect 16268 31154 16324 31166
rect 15932 30996 15988 31006
rect 15932 30902 15988 30940
rect 16492 30994 16548 31006
rect 16492 30942 16494 30994
rect 16546 30942 16548 30994
rect 16380 30884 16436 30894
rect 16044 30882 16436 30884
rect 16044 30830 16382 30882
rect 16434 30830 16436 30882
rect 16044 30828 16436 30830
rect 15820 30436 15876 30446
rect 16044 30436 16100 30828
rect 16380 30818 16436 30828
rect 15820 30434 16100 30436
rect 15820 30382 15822 30434
rect 15874 30382 16100 30434
rect 15820 30380 16100 30382
rect 15820 30370 15876 30380
rect 16156 30324 16212 30334
rect 16156 30230 16212 30268
rect 15708 30100 15764 30110
rect 15708 30006 15764 30044
rect 15596 29986 15652 29998
rect 15596 29934 15598 29986
rect 15650 29934 15652 29986
rect 15596 28980 15652 29934
rect 15596 28924 15988 28980
rect 15932 28866 15988 28924
rect 15932 28814 15934 28866
rect 15986 28814 15988 28866
rect 15372 28588 15652 28644
rect 15372 28420 15428 28430
rect 15260 28418 15428 28420
rect 15260 28366 15374 28418
rect 15426 28366 15428 28418
rect 15260 28364 15428 28366
rect 15372 27972 15428 28364
rect 15372 27906 15428 27916
rect 15148 27794 15204 27804
rect 14476 26786 14532 26796
rect 15372 27076 15428 27086
rect 15372 26402 15428 27020
rect 15372 26350 15374 26402
rect 15426 26350 15428 26402
rect 15372 26338 15428 26350
rect 15148 26178 15204 26190
rect 15148 26126 15150 26178
rect 15202 26126 15204 26178
rect 14588 25620 14644 25630
rect 14140 25454 14142 25506
rect 14194 25454 14196 25506
rect 14140 24052 14196 25454
rect 14364 25508 14420 25518
rect 14364 25414 14420 25452
rect 14588 25506 14644 25564
rect 14588 25454 14590 25506
rect 14642 25454 14644 25506
rect 14140 23996 14532 24052
rect 14364 23268 14420 23278
rect 14364 23174 14420 23212
rect 11340 22988 11732 23044
rect 14476 23154 14532 23996
rect 14476 23102 14478 23154
rect 14530 23102 14532 23154
rect 11340 21364 11396 22988
rect 11452 21810 11508 21822
rect 11452 21758 11454 21810
rect 11506 21758 11508 21810
rect 11452 21588 11508 21758
rect 11564 21698 11620 21710
rect 12684 21700 12740 21710
rect 11564 21646 11566 21698
rect 11618 21646 11620 21698
rect 11564 21588 11620 21646
rect 12348 21698 12740 21700
rect 12348 21646 12686 21698
rect 12738 21646 12740 21698
rect 12348 21644 12740 21646
rect 11564 21532 11732 21588
rect 11452 21522 11508 21532
rect 11340 21308 11620 21364
rect 11452 20802 11508 20814
rect 11452 20750 11454 20802
rect 11506 20750 11508 20802
rect 11340 20692 11396 20702
rect 11340 20598 11396 20636
rect 10892 20524 11284 20580
rect 10780 20178 10836 20188
rect 10444 19180 10724 19236
rect 10892 19796 10948 19806
rect 10444 18788 10500 19180
rect 10892 19122 10948 19740
rect 10892 19070 10894 19122
rect 10946 19070 10948 19122
rect 10892 19058 10948 19070
rect 9884 17666 9940 18396
rect 10332 18732 10500 18788
rect 10108 18340 10164 18350
rect 10108 18246 10164 18284
rect 9884 17614 9886 17666
rect 9938 17614 9940 17666
rect 9884 17602 9940 17614
rect 10108 17666 10164 17678
rect 10108 17614 10110 17666
rect 10162 17614 10164 17666
rect 9996 17554 10052 17566
rect 9996 17502 9998 17554
rect 10050 17502 10052 17554
rect 9996 17444 10052 17502
rect 9884 17388 10052 17444
rect 10108 17556 10164 17614
rect 9884 17106 9940 17388
rect 10108 17332 10164 17500
rect 9884 17054 9886 17106
rect 9938 17054 9940 17106
rect 9548 16884 9604 16894
rect 9548 16790 9604 16828
rect 9884 16772 9940 17054
rect 9884 16706 9940 16716
rect 9996 17276 10164 17332
rect 9548 16324 9604 16334
rect 9548 16322 9940 16324
rect 9548 16270 9550 16322
rect 9602 16270 9940 16322
rect 9548 16268 9940 16270
rect 9548 16258 9604 16268
rect 9772 16100 9828 16138
rect 9436 16044 9716 16100
rect 8652 14476 9380 14532
rect 9548 15314 9604 15326
rect 9548 15262 9550 15314
rect 9602 15262 9604 15314
rect 8652 14418 8708 14476
rect 8652 14366 8654 14418
rect 8706 14366 8708 14418
rect 8540 13860 8596 13870
rect 8428 13858 8596 13860
rect 8428 13806 8542 13858
rect 8594 13806 8596 13858
rect 8428 13804 8596 13806
rect 8092 13188 8148 13198
rect 7980 12962 8036 12974
rect 7980 12910 7982 12962
rect 8034 12910 8036 12962
rect 7980 12740 8036 12910
rect 7980 12404 8036 12684
rect 8092 12738 8148 13132
rect 8428 12964 8484 13804
rect 8540 13794 8596 13804
rect 8652 13746 8708 14366
rect 8652 13694 8654 13746
rect 8706 13694 8708 13746
rect 8092 12686 8094 12738
rect 8146 12686 8148 12738
rect 8092 12516 8148 12686
rect 8316 12908 8484 12964
rect 8540 13522 8596 13534
rect 8540 13470 8542 13522
rect 8594 13470 8596 13522
rect 8540 12964 8596 13470
rect 8652 13300 8708 13694
rect 8652 13234 8708 13244
rect 8764 14306 8820 14318
rect 8764 14254 8766 14306
rect 8818 14254 8820 14306
rect 8764 13860 8820 14254
rect 9548 13860 9604 15262
rect 9660 15092 9716 16044
rect 9772 16034 9828 16044
rect 9772 15876 9828 15886
rect 9772 15426 9828 15820
rect 9884 15538 9940 16268
rect 9884 15486 9886 15538
rect 9938 15486 9940 15538
rect 9884 15474 9940 15486
rect 9996 15538 10052 17276
rect 10332 17108 10388 18732
rect 10444 18564 10500 18574
rect 10444 17780 10500 18508
rect 10556 17836 10836 17892
rect 10556 17780 10612 17836
rect 10444 17778 10612 17780
rect 10444 17726 10558 17778
rect 10610 17726 10612 17778
rect 10444 17724 10612 17726
rect 10556 17714 10612 17724
rect 10332 17014 10388 17052
rect 10668 17556 10724 17566
rect 10220 16884 10276 16894
rect 10220 16790 10276 16828
rect 9996 15486 9998 15538
rect 10050 15486 10052 15538
rect 9996 15474 10052 15486
rect 10220 16100 10276 16110
rect 9772 15374 9774 15426
rect 9826 15374 9828 15426
rect 9772 15316 9828 15374
rect 9772 15260 9940 15316
rect 9660 15036 9828 15092
rect 8764 13858 9604 13860
rect 8764 13806 9550 13858
rect 9602 13806 9604 13858
rect 8764 13804 9604 13806
rect 8652 12964 8708 12974
rect 8540 12962 8708 12964
rect 8540 12910 8654 12962
rect 8706 12910 8708 12962
rect 8540 12908 8708 12910
rect 8316 12740 8372 12908
rect 8652 12898 8708 12908
rect 8316 12674 8372 12684
rect 8092 12460 8596 12516
rect 7980 12338 8036 12348
rect 8540 12178 8596 12460
rect 8764 12292 8820 13804
rect 9548 13794 9604 13804
rect 9772 13746 9828 15036
rect 9772 13694 9774 13746
rect 9826 13694 9828 13746
rect 9660 13636 9716 13646
rect 9660 13542 9716 13580
rect 9212 13524 9268 13534
rect 9212 13074 9268 13468
rect 9772 13412 9828 13694
rect 9660 13356 9828 13412
rect 9660 13188 9716 13356
rect 9660 13122 9716 13132
rect 9212 13022 9214 13074
rect 9266 13022 9268 13074
rect 9212 13010 9268 13022
rect 9772 13076 9828 13086
rect 9884 13076 9940 15260
rect 10108 15314 10164 15326
rect 10108 15262 10110 15314
rect 10162 15262 10164 15314
rect 10108 13972 10164 15262
rect 10108 13906 10164 13916
rect 10220 13748 10276 16044
rect 10668 15148 10724 17500
rect 10108 13746 10276 13748
rect 10108 13694 10222 13746
rect 10274 13694 10276 13746
rect 10108 13692 10276 13694
rect 9996 13524 10052 13534
rect 9996 13430 10052 13468
rect 9828 13020 9940 13076
rect 9996 13300 10052 13310
rect 9772 13010 9828 13020
rect 8876 12852 8932 12862
rect 9884 12852 9940 12862
rect 8876 12758 8932 12796
rect 9324 12850 9940 12852
rect 9324 12798 9886 12850
rect 9938 12798 9940 12850
rect 9324 12796 9940 12798
rect 9100 12740 9156 12750
rect 8876 12292 8932 12302
rect 8764 12290 8932 12292
rect 8764 12238 8878 12290
rect 8930 12238 8932 12290
rect 8764 12236 8932 12238
rect 8876 12226 8932 12236
rect 8540 12126 8542 12178
rect 8594 12126 8596 12178
rect 8540 12114 8596 12126
rect 9100 12180 9156 12684
rect 9212 12738 9268 12750
rect 9212 12686 9214 12738
rect 9266 12686 9268 12738
rect 9212 12628 9268 12686
rect 9212 12562 9268 12572
rect 9100 12114 9156 12124
rect 8764 12066 8820 12078
rect 8764 12014 8766 12066
rect 8818 12014 8820 12066
rect 8764 11396 8820 12014
rect 8428 11394 8820 11396
rect 8428 11342 8766 11394
rect 8818 11342 8820 11394
rect 8428 11340 8820 11342
rect 8428 10834 8484 11340
rect 8764 11330 8820 11340
rect 9100 11396 9156 11406
rect 9324 11396 9380 12796
rect 9884 12786 9940 12796
rect 9996 12292 10052 13244
rect 10108 12964 10164 13692
rect 10220 13682 10276 13692
rect 10332 15092 10724 15148
rect 10108 12898 10164 12908
rect 10220 12964 10276 12974
rect 10332 12964 10388 15092
rect 10556 13972 10612 13982
rect 10444 13188 10500 13226
rect 10444 13122 10500 13132
rect 10220 12962 10388 12964
rect 10220 12910 10222 12962
rect 10274 12910 10388 12962
rect 10220 12908 10388 12910
rect 10444 12964 10500 12974
rect 10220 12898 10276 12908
rect 10444 12870 10500 12908
rect 10220 12738 10276 12750
rect 10220 12686 10222 12738
rect 10274 12686 10276 12738
rect 10108 12292 10164 12302
rect 9996 12290 10164 12292
rect 9996 12238 10110 12290
rect 10162 12238 10164 12290
rect 9996 12236 10164 12238
rect 10108 12226 10164 12236
rect 9548 12180 9604 12190
rect 9548 12086 9604 12124
rect 9996 11732 10052 11742
rect 9100 11394 9604 11396
rect 9100 11342 9102 11394
rect 9154 11342 9604 11394
rect 9100 11340 9604 11342
rect 9100 11330 9156 11340
rect 8876 11172 8932 11182
rect 8876 11078 8932 11116
rect 8428 10782 8430 10834
rect 8482 10782 8484 10834
rect 8428 10770 8484 10782
rect 9548 10722 9604 11340
rect 9996 11172 10052 11676
rect 10220 11396 10276 12686
rect 10556 12628 10612 13916
rect 10556 12562 10612 12572
rect 10780 12292 10836 17836
rect 11116 17108 11172 17118
rect 11004 17106 11172 17108
rect 11004 17054 11118 17106
rect 11170 17054 11172 17106
rect 11004 17052 11172 17054
rect 11004 16436 11060 17052
rect 11116 17042 11172 17052
rect 11004 16370 11060 16380
rect 11116 16882 11172 16894
rect 11116 16830 11118 16882
rect 11170 16830 11172 16882
rect 11116 16100 11172 16830
rect 11116 16034 11172 16044
rect 11228 15148 11284 20524
rect 11452 17556 11508 20750
rect 11564 19236 11620 21308
rect 11676 19684 11732 21532
rect 11788 21586 11844 21598
rect 11788 21534 11790 21586
rect 11842 21534 11844 21586
rect 11788 21476 11844 21534
rect 12124 21588 12180 21598
rect 12124 21494 12180 21532
rect 11788 19906 11844 21420
rect 12348 20578 12404 21644
rect 12684 21634 12740 21644
rect 13692 21700 13748 21710
rect 13692 21606 13748 21644
rect 13804 21586 13860 21598
rect 13804 21534 13806 21586
rect 13858 21534 13860 21586
rect 13804 20914 13860 21534
rect 13804 20862 13806 20914
rect 13858 20862 13860 20914
rect 13804 20850 13860 20862
rect 12684 20802 12740 20814
rect 12684 20750 12686 20802
rect 12738 20750 12740 20802
rect 12348 20526 12350 20578
rect 12402 20526 12404 20578
rect 12348 20514 12404 20526
rect 12572 20580 12628 20590
rect 12572 20486 12628 20524
rect 12684 20468 12740 20750
rect 12684 20402 12740 20412
rect 13468 20802 13524 20814
rect 13468 20750 13470 20802
rect 13522 20750 13524 20802
rect 12236 20244 12292 20254
rect 11788 19854 11790 19906
rect 11842 19854 11844 19906
rect 11788 19842 11844 19854
rect 12124 20018 12180 20030
rect 12124 19966 12126 20018
rect 12178 19966 12180 20018
rect 12124 19684 12180 19966
rect 11676 19628 12180 19684
rect 11676 19236 11732 19246
rect 11564 19234 11732 19236
rect 11564 19182 11678 19234
rect 11730 19182 11732 19234
rect 11564 19180 11732 19182
rect 11676 19170 11732 19180
rect 11900 19012 11956 19022
rect 11900 18918 11956 18956
rect 12124 18900 12180 19628
rect 12124 18834 12180 18844
rect 12236 17780 12292 20188
rect 12348 20132 12404 20142
rect 12348 17892 12404 20076
rect 12908 20020 12964 20030
rect 12908 19926 12964 19964
rect 13468 18564 13524 20750
rect 13916 20692 13972 20702
rect 14476 20692 14532 23102
rect 13916 20690 14532 20692
rect 13916 20638 13918 20690
rect 13970 20638 14532 20690
rect 13916 20636 14532 20638
rect 14588 23268 14644 25454
rect 13916 20626 13972 20636
rect 14252 20468 14308 20478
rect 13804 20018 13860 20030
rect 13804 19966 13806 20018
rect 13858 19966 13860 20018
rect 13804 18788 13860 19966
rect 14252 20018 14308 20412
rect 14588 20468 14644 23212
rect 15148 25508 15204 26126
rect 14924 23156 14980 23166
rect 15148 23156 15204 25452
rect 15596 25060 15652 28588
rect 15708 28642 15764 28654
rect 15708 28590 15710 28642
rect 15762 28590 15764 28642
rect 15708 28308 15764 28590
rect 15932 28532 15988 28814
rect 15932 28466 15988 28476
rect 16268 28642 16324 28654
rect 16268 28590 16270 28642
rect 16322 28590 16324 28642
rect 16268 28308 16324 28590
rect 15708 28252 16324 28308
rect 16492 28642 16548 30942
rect 16828 30994 16884 31006
rect 16828 30942 16830 30994
rect 16882 30942 16884 30994
rect 16828 30884 16884 30942
rect 16828 30818 16884 30828
rect 16492 28590 16494 28642
rect 16546 28590 16548 28642
rect 15708 26292 15764 28252
rect 16492 27972 16548 28590
rect 16716 28644 16772 28654
rect 16716 28550 16772 28588
rect 16492 27906 16548 27916
rect 16604 27860 16660 27870
rect 16604 27186 16660 27804
rect 16604 27134 16606 27186
rect 16658 27134 16660 27186
rect 16604 27122 16660 27134
rect 16604 26402 16660 26414
rect 16604 26350 16606 26402
rect 16658 26350 16660 26402
rect 16268 26292 16324 26302
rect 15708 26226 15764 26236
rect 16044 26290 16324 26292
rect 16044 26238 16270 26290
rect 16322 26238 16324 26290
rect 16044 26236 16324 26238
rect 16044 25508 16100 26236
rect 16268 26226 16324 26236
rect 16604 26292 16660 26350
rect 16604 26226 16660 26236
rect 16044 25506 16436 25508
rect 16044 25454 16046 25506
rect 16098 25454 16436 25506
rect 16044 25452 16436 25454
rect 16044 25442 16100 25452
rect 15708 25396 15764 25406
rect 15708 25302 15764 25340
rect 15596 25004 15988 25060
rect 15260 23268 15316 23278
rect 15260 23174 15316 23212
rect 14924 23154 15204 23156
rect 14924 23102 14926 23154
rect 14978 23102 15204 23154
rect 14924 23100 15204 23102
rect 14924 20802 14980 23100
rect 15820 21810 15876 25004
rect 15932 24948 15988 25004
rect 15932 24946 16212 24948
rect 15932 24894 15934 24946
rect 15986 24894 16212 24946
rect 15932 24892 16212 24894
rect 15932 24882 15988 24892
rect 16156 24722 16212 24892
rect 16380 24946 16436 25452
rect 16380 24894 16382 24946
rect 16434 24894 16436 24946
rect 16380 24882 16436 24894
rect 16156 24670 16158 24722
rect 16210 24670 16212 24722
rect 16156 24658 16212 24670
rect 16604 24724 16660 24734
rect 16604 24630 16660 24668
rect 16828 24722 16884 24734
rect 16828 24670 16830 24722
rect 16882 24670 16884 24722
rect 16828 23828 16884 24670
rect 16828 23762 16884 23772
rect 16828 23604 16884 23614
rect 16044 22932 16100 22942
rect 16268 22932 16324 22942
rect 16044 22930 16268 22932
rect 16044 22878 16046 22930
rect 16098 22878 16268 22930
rect 16044 22876 16268 22878
rect 16044 22866 16100 22876
rect 16268 22482 16324 22876
rect 16828 22594 16884 23548
rect 16828 22542 16830 22594
rect 16882 22542 16884 22594
rect 16828 22530 16884 22542
rect 16268 22430 16270 22482
rect 16322 22430 16324 22482
rect 16268 22418 16324 22430
rect 16492 22484 16548 22494
rect 16492 22390 16548 22428
rect 16940 22372 16996 32508
rect 17052 22484 17108 33516
rect 17836 33460 17892 34636
rect 17836 33394 17892 33404
rect 19516 32788 19572 37436
rect 19740 37426 19796 37436
rect 20076 37266 20132 37436
rect 20076 37214 20078 37266
rect 20130 37214 20132 37266
rect 20076 37202 20132 37214
rect 20860 37156 20916 37166
rect 20860 37154 21588 37156
rect 20860 37102 20862 37154
rect 20914 37102 21588 37154
rect 20860 37100 21588 37102
rect 20860 37090 20916 37100
rect 21532 36706 21588 37100
rect 21532 36654 21534 36706
rect 21586 36654 21588 36706
rect 21532 36642 21588 36654
rect 21868 36706 21924 37884
rect 24892 37940 24948 37950
rect 24892 37846 24948 37884
rect 24332 37380 24388 37390
rect 22988 37268 23044 37278
rect 22988 37154 23044 37212
rect 24220 37268 24276 37278
rect 22988 37102 22990 37154
rect 23042 37102 23044 37154
rect 22988 37090 23044 37102
rect 23660 37154 23716 37166
rect 23660 37102 23662 37154
rect 23714 37102 23716 37154
rect 21868 36654 21870 36706
rect 21922 36654 21924 36706
rect 21868 36642 21924 36654
rect 20524 36484 20580 36494
rect 19628 36148 19684 36158
rect 19628 35810 19684 36092
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19628 35758 19630 35810
rect 19682 35758 19684 35810
rect 19628 35746 19684 35758
rect 20076 35812 20132 35822
rect 20076 35698 20132 35756
rect 20076 35646 20078 35698
rect 20130 35646 20132 35698
rect 20076 35634 20132 35646
rect 20524 35698 20580 36428
rect 20860 36260 20916 36270
rect 21644 36260 21700 36270
rect 20860 36258 21700 36260
rect 20860 36206 20862 36258
rect 20914 36206 21646 36258
rect 21698 36206 21700 36258
rect 20860 36204 21700 36206
rect 20860 36194 20916 36204
rect 20524 35646 20526 35698
rect 20578 35646 20580 35698
rect 20524 35634 20580 35646
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32788 19684 32798
rect 19516 32786 20020 32788
rect 19516 32734 19630 32786
rect 19682 32734 20020 32786
rect 19516 32732 20020 32734
rect 18956 31668 19012 31678
rect 17948 30996 18004 31006
rect 17948 30902 18004 30940
rect 17500 30884 17556 30894
rect 17276 28644 17332 28654
rect 17276 28550 17332 28588
rect 17388 28532 17444 28542
rect 17388 28438 17444 28476
rect 17164 28418 17220 28430
rect 17164 28366 17166 28418
rect 17218 28366 17220 28418
rect 17164 27972 17220 28366
rect 17164 27906 17220 27916
rect 17164 27748 17220 27758
rect 17164 27076 17220 27692
rect 17164 26982 17220 27020
rect 17388 26292 17444 26302
rect 17388 26198 17444 26236
rect 17500 24836 17556 30828
rect 18956 30324 19012 31612
rect 18956 30210 19012 30268
rect 18956 30158 18958 30210
rect 19010 30158 19012 30210
rect 18956 30146 19012 30158
rect 19628 30324 19684 32732
rect 19964 32562 20020 32732
rect 19964 32510 19966 32562
rect 20018 32510 20020 32562
rect 19964 32498 20020 32510
rect 20748 32452 20804 32462
rect 20748 32450 21588 32452
rect 20748 32398 20750 32450
rect 20802 32398 21588 32450
rect 20748 32396 21588 32398
rect 20748 32386 20804 32396
rect 21532 32002 21588 32396
rect 21532 31950 21534 32002
rect 21586 31950 21588 32002
rect 21532 31938 21588 31950
rect 19964 31778 20020 31790
rect 19964 31726 19966 31778
rect 20018 31726 20020 31778
rect 19964 31556 20020 31726
rect 20748 31556 20804 31566
rect 19964 31500 20244 31556
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 30884 20244 31500
rect 20748 31462 20804 31500
rect 21644 31556 21700 36204
rect 23660 35700 23716 37102
rect 24220 36932 24276 37212
rect 24332 37266 24388 37324
rect 25564 37380 25620 37998
rect 25788 38050 25844 38062
rect 25788 37998 25790 38050
rect 25842 37998 25844 38050
rect 25788 37828 25844 37998
rect 25788 37762 25844 37772
rect 25620 37324 25732 37380
rect 25564 37286 25620 37324
rect 24332 37214 24334 37266
rect 24386 37214 24388 37266
rect 24332 37202 24388 37214
rect 25228 37268 25284 37278
rect 25228 37174 25284 37212
rect 24556 37154 24612 37166
rect 24556 37102 24558 37154
rect 24610 37102 24612 37154
rect 24556 37044 24612 37102
rect 24108 36876 24276 36932
rect 24332 36988 24556 37044
rect 24108 36260 24164 36876
rect 24220 36706 24276 36718
rect 24220 36654 24222 36706
rect 24274 36654 24276 36706
rect 24220 36484 24276 36654
rect 24220 36418 24276 36428
rect 24332 36482 24388 36988
rect 24556 36978 24612 36988
rect 24332 36430 24334 36482
rect 24386 36430 24388 36482
rect 24332 36418 24388 36430
rect 25564 36484 25620 36494
rect 24220 36260 24276 36270
rect 24108 36258 24276 36260
rect 24108 36206 24222 36258
rect 24274 36206 24276 36258
rect 24108 36204 24276 36206
rect 24220 36194 24276 36204
rect 23660 35634 23716 35644
rect 25564 34914 25620 36428
rect 25676 36260 25732 37324
rect 25676 36194 25732 36204
rect 25564 34862 25566 34914
rect 25618 34862 25620 34914
rect 25564 34850 25620 34862
rect 25788 34804 25844 34814
rect 25788 34710 25844 34748
rect 23772 34692 23828 34702
rect 23100 33460 23156 33470
rect 23100 33366 23156 33404
rect 23772 33346 23828 34636
rect 25676 34692 25732 34702
rect 25676 34598 25732 34636
rect 25900 34468 25956 40236
rect 26012 40226 26068 40236
rect 28140 40292 28196 40302
rect 28140 40290 28420 40292
rect 28140 40238 28142 40290
rect 28194 40238 28420 40290
rect 28140 40236 28420 40238
rect 28140 40226 28196 40236
rect 28364 40180 28420 40236
rect 28252 39396 28308 39406
rect 28252 39302 28308 39340
rect 26348 37828 26404 37838
rect 26124 37772 26348 37828
rect 26012 34692 26068 34702
rect 26012 34598 26068 34636
rect 25676 34412 25956 34468
rect 23772 33294 23774 33346
rect 23826 33294 23828 33346
rect 23772 33282 23828 33294
rect 25116 33458 25172 33470
rect 25116 33406 25118 33458
rect 25170 33406 25172 33458
rect 23884 33236 23940 33246
rect 22876 32564 22932 32574
rect 22876 32450 22932 32508
rect 23884 32564 23940 33180
rect 24668 33236 24724 33246
rect 24668 33142 24724 33180
rect 25116 32788 25172 33406
rect 25116 32722 25172 32732
rect 23884 32470 23940 32508
rect 24108 32564 24164 32574
rect 24108 32470 24164 32508
rect 23212 32452 23268 32462
rect 22876 32398 22878 32450
rect 22930 32398 22932 32450
rect 22876 32386 22932 32398
rect 22988 32450 23268 32452
rect 22988 32398 23214 32450
rect 23266 32398 23268 32450
rect 22988 32396 23268 32398
rect 22988 32228 23044 32396
rect 23212 32386 23268 32396
rect 21868 32172 23044 32228
rect 21868 32002 21924 32172
rect 21868 31950 21870 32002
rect 21922 31950 21924 32002
rect 21868 31938 21924 31950
rect 25564 31892 25620 31902
rect 25340 31836 25564 31892
rect 25340 31666 25396 31836
rect 25564 31826 25620 31836
rect 25676 31890 25732 34412
rect 26124 32450 26180 37772
rect 26348 37734 26404 37772
rect 27580 37380 27636 37390
rect 27580 37266 27636 37324
rect 27580 37214 27582 37266
rect 27634 37214 27636 37266
rect 27580 37202 27636 37214
rect 28252 37156 28308 37166
rect 27916 37154 28308 37156
rect 27916 37102 28254 37154
rect 28306 37102 28308 37154
rect 27916 37100 28308 37102
rect 27916 36706 27972 37100
rect 28252 37090 28308 37100
rect 27916 36654 27918 36706
rect 27970 36654 27972 36706
rect 27916 36642 27972 36654
rect 27132 36596 27188 36606
rect 27132 36594 27860 36596
rect 27132 36542 27134 36594
rect 27186 36542 27860 36594
rect 27132 36540 27860 36542
rect 27132 36530 27188 36540
rect 26796 36482 26852 36494
rect 26796 36430 26798 36482
rect 26850 36430 26852 36482
rect 26796 36372 26852 36430
rect 26572 36260 26628 36270
rect 26572 34354 26628 36204
rect 26572 34302 26574 34354
rect 26626 34302 26628 34354
rect 26572 34290 26628 34302
rect 26796 34356 26852 36316
rect 26908 36370 26964 36382
rect 26908 36318 26910 36370
rect 26962 36318 26964 36370
rect 26908 36260 26964 36318
rect 27244 36370 27300 36382
rect 27244 36318 27246 36370
rect 27298 36318 27300 36370
rect 27244 36260 27300 36318
rect 27580 36370 27636 36382
rect 27580 36318 27582 36370
rect 27634 36318 27636 36370
rect 27468 36260 27524 36270
rect 27244 36204 27468 36260
rect 26908 36194 26964 36204
rect 27468 36194 27524 36204
rect 27356 34804 27412 34814
rect 27132 34692 27188 34702
rect 27132 34690 27300 34692
rect 27132 34638 27134 34690
rect 27186 34638 27300 34690
rect 27132 34636 27300 34638
rect 27132 34626 27188 34636
rect 26796 34354 27188 34356
rect 26796 34302 26798 34354
rect 26850 34302 27188 34354
rect 26796 34300 27188 34302
rect 26796 34290 26852 34300
rect 27132 34244 27188 34300
rect 26348 34132 26404 34142
rect 26348 34038 26404 34076
rect 26908 34132 26964 34142
rect 26684 34018 26740 34030
rect 26684 33966 26686 34018
rect 26738 33966 26740 34018
rect 26684 33234 26740 33966
rect 26684 33182 26686 33234
rect 26738 33182 26740 33234
rect 26124 32398 26126 32450
rect 26178 32398 26180 32450
rect 26124 32386 26180 32398
rect 26572 32562 26628 32574
rect 26572 32510 26574 32562
rect 26626 32510 26628 32562
rect 26572 32452 26628 32510
rect 26684 32564 26740 33182
rect 26796 33124 26852 33134
rect 26796 33030 26852 33068
rect 26684 32498 26740 32508
rect 26572 32386 26628 32396
rect 26908 32116 26964 34076
rect 27132 34130 27188 34188
rect 27132 34078 27134 34130
rect 27186 34078 27188 34130
rect 27132 34066 27188 34078
rect 27244 34132 27300 34636
rect 27356 34354 27412 34748
rect 27356 34302 27358 34354
rect 27410 34302 27412 34354
rect 27356 34290 27412 34302
rect 27244 34066 27300 34076
rect 27468 34132 27524 34142
rect 27468 34038 27524 34076
rect 27580 33684 27636 36318
rect 27804 36370 27860 36540
rect 28364 36484 28420 40124
rect 28476 37380 28532 40348
rect 29260 40402 29316 40414
rect 29260 40350 29262 40402
rect 29314 40350 29316 40402
rect 29260 39396 29316 40350
rect 31388 40290 31444 41916
rect 32508 41972 32564 41982
rect 32508 41878 32564 41916
rect 36092 41860 36148 45200
rect 36092 41794 36148 41804
rect 36316 41970 36372 41982
rect 36316 41918 36318 41970
rect 36370 41918 36372 41970
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 32620 40628 32676 40638
rect 32620 40534 32676 40572
rect 34188 40628 34244 40638
rect 34188 40514 34244 40572
rect 34188 40462 34190 40514
rect 34242 40462 34244 40514
rect 34188 40450 34244 40462
rect 31836 40404 31892 40414
rect 31724 40402 31892 40404
rect 31724 40350 31838 40402
rect 31890 40350 31892 40402
rect 31724 40348 31892 40350
rect 31388 40238 31390 40290
rect 31442 40238 31444 40290
rect 31388 40226 31444 40238
rect 31500 40292 31556 40302
rect 31500 39618 31556 40236
rect 31500 39566 31502 39618
rect 31554 39566 31556 39618
rect 31500 39554 31556 39566
rect 29260 39330 29316 39340
rect 28476 37314 28532 37324
rect 30268 37380 30324 37390
rect 27804 36318 27806 36370
rect 27858 36318 27860 36370
rect 27804 36306 27860 36318
rect 28252 36428 28420 36484
rect 29484 36484 29540 36494
rect 27692 34692 27748 34702
rect 27692 34354 27748 34636
rect 27692 34302 27694 34354
rect 27746 34302 27748 34354
rect 27692 34290 27748 34302
rect 27916 34244 27972 34254
rect 27916 34150 27972 34188
rect 28028 34132 28084 34142
rect 28028 34038 28084 34076
rect 27020 33628 27636 33684
rect 27020 33346 27076 33628
rect 27020 33294 27022 33346
rect 27074 33294 27076 33346
rect 27020 33282 27076 33294
rect 27468 33124 27524 33134
rect 27132 33012 27188 33022
rect 27020 32452 27076 32462
rect 27020 32358 27076 32396
rect 27020 32116 27076 32126
rect 26908 32060 27020 32116
rect 26236 31892 26292 31902
rect 25676 31838 25678 31890
rect 25730 31838 25732 31890
rect 25676 31826 25732 31838
rect 25788 31890 26292 31892
rect 25788 31838 26238 31890
rect 26290 31838 26292 31890
rect 25788 31836 26292 31838
rect 25788 31778 25844 31836
rect 26236 31826 26292 31836
rect 25788 31726 25790 31778
rect 25842 31726 25844 31778
rect 25788 31714 25844 31726
rect 26684 31780 26740 31790
rect 26684 31686 26740 31724
rect 25340 31614 25342 31666
rect 25394 31614 25396 31666
rect 25340 31602 25396 31614
rect 26124 31666 26180 31678
rect 26124 31614 26126 31666
rect 26178 31614 26180 31666
rect 20188 30790 20244 30828
rect 19628 30210 19684 30268
rect 21644 30324 21700 31500
rect 24108 31556 24164 31566
rect 23436 31444 23492 31454
rect 21644 30258 21700 30268
rect 22540 30324 22596 30334
rect 19628 30158 19630 30210
rect 19682 30158 19684 30210
rect 19628 30146 19684 30158
rect 18284 30100 18340 30110
rect 18284 30006 18340 30044
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20300 28756 20356 28766
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19740 27748 19796 27758
rect 19740 27654 19796 27692
rect 17724 27188 17780 27198
rect 17724 26402 17780 27132
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 18732 26516 18788 26526
rect 18732 26422 18788 26460
rect 17724 26350 17726 26402
rect 17778 26350 17780 26402
rect 17724 24948 17780 26350
rect 18396 26290 18452 26302
rect 18396 26238 18398 26290
rect 18450 26238 18452 26290
rect 17724 24882 17780 24892
rect 18060 25284 18116 25294
rect 18396 25284 18452 26238
rect 18060 25282 18452 25284
rect 18060 25230 18062 25282
rect 18114 25230 18452 25282
rect 18060 25228 18452 25230
rect 18060 25060 18116 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 17500 24770 17556 24780
rect 17388 24724 17444 24734
rect 17388 24630 17444 24668
rect 17948 24610 18004 24622
rect 17948 24558 17950 24610
rect 18002 24558 18004 24610
rect 17724 24498 17780 24510
rect 17724 24446 17726 24498
rect 17778 24446 17780 24498
rect 17724 23604 17780 24446
rect 17948 24276 18004 24558
rect 17948 24210 18004 24220
rect 18060 24164 18116 25004
rect 19516 24276 19572 24286
rect 18060 24108 18564 24164
rect 17948 24052 18004 24062
rect 18060 24052 18116 24108
rect 17948 24050 18116 24052
rect 17948 23998 17950 24050
rect 18002 23998 18116 24050
rect 17948 23996 18116 23998
rect 17948 23986 18004 23996
rect 17724 23538 17780 23548
rect 18284 23940 18340 23950
rect 18284 23604 18340 23884
rect 18508 23938 18564 24108
rect 18508 23886 18510 23938
rect 18562 23886 18564 23938
rect 18508 23874 18564 23886
rect 18284 23538 18340 23548
rect 18732 23828 18788 23838
rect 18620 23154 18676 23166
rect 18620 23102 18622 23154
rect 18674 23102 18676 23154
rect 18508 23042 18564 23054
rect 18508 22990 18510 23042
rect 18562 22990 18564 23042
rect 17836 22930 17892 22942
rect 17836 22878 17838 22930
rect 17890 22878 17892 22930
rect 17164 22484 17220 22494
rect 17052 22482 17220 22484
rect 17052 22430 17166 22482
rect 17218 22430 17220 22482
rect 17052 22428 17220 22430
rect 16940 22316 17108 22372
rect 15820 21758 15822 21810
rect 15874 21758 15876 21810
rect 14924 20750 14926 20802
rect 14978 20750 14980 20802
rect 14924 20738 14980 20750
rect 15372 21474 15428 21486
rect 15372 21422 15374 21474
rect 15426 21422 15428 21474
rect 15372 21364 15428 21422
rect 15260 20692 15316 20702
rect 14588 20402 14644 20412
rect 14700 20578 14756 20590
rect 14700 20526 14702 20578
rect 14754 20526 14756 20578
rect 14252 19966 14254 20018
rect 14306 19966 14308 20018
rect 14252 19954 14308 19966
rect 13804 18722 13860 18732
rect 13132 18508 13524 18564
rect 12348 17890 12964 17892
rect 12348 17838 12350 17890
rect 12402 17838 12964 17890
rect 12348 17836 12964 17838
rect 12348 17826 12404 17836
rect 11452 17490 11508 17500
rect 12012 17778 12292 17780
rect 12012 17726 12238 17778
rect 12290 17726 12292 17778
rect 12012 17724 12292 17726
rect 11340 17108 11396 17118
rect 11396 17052 11620 17108
rect 11340 17042 11396 17052
rect 11564 16882 11620 17052
rect 11900 16996 11956 17006
rect 11900 16902 11956 16940
rect 11564 16830 11566 16882
rect 11618 16830 11620 16882
rect 11564 16818 11620 16830
rect 11452 16660 11508 16670
rect 11452 16566 11508 16604
rect 11676 16100 11732 16110
rect 11228 15092 11396 15148
rect 11004 14644 11060 14654
rect 11340 14644 11396 15092
rect 11004 14642 11396 14644
rect 11004 14590 11006 14642
rect 11058 14590 11396 14642
rect 11004 14588 11396 14590
rect 11004 14578 11060 14588
rect 11340 14530 11396 14588
rect 11340 14478 11342 14530
rect 11394 14478 11396 14530
rect 11340 13972 11396 14478
rect 11676 14418 11732 16044
rect 12012 15148 12068 17724
rect 12236 17714 12292 17724
rect 12348 16660 12404 16670
rect 12124 16212 12180 16222
rect 12124 16098 12180 16156
rect 12348 16210 12404 16604
rect 12348 16158 12350 16210
rect 12402 16158 12404 16210
rect 12348 16146 12404 16158
rect 12124 16046 12126 16098
rect 12178 16046 12180 16098
rect 12124 16034 12180 16046
rect 12460 16100 12516 16110
rect 12460 16006 12516 16044
rect 12684 16100 12740 16110
rect 12684 16098 12852 16100
rect 12684 16046 12686 16098
rect 12738 16046 12852 16098
rect 12684 16044 12852 16046
rect 12684 16034 12740 16044
rect 12236 15988 12292 15998
rect 12236 15894 12292 15932
rect 12796 15988 12852 16044
rect 12796 15540 12852 15932
rect 12908 15764 12964 17836
rect 13132 17106 13188 18508
rect 14700 18452 14756 20526
rect 15260 19906 15316 20636
rect 15372 20690 15428 21308
rect 15372 20638 15374 20690
rect 15426 20638 15428 20690
rect 15372 20626 15428 20638
rect 15820 20188 15876 21758
rect 16492 21588 16548 21598
rect 16492 21586 16772 21588
rect 16492 21534 16494 21586
rect 16546 21534 16772 21586
rect 16492 21532 16772 21534
rect 16492 21522 16548 21532
rect 16268 21364 16324 21374
rect 16268 21270 16324 21308
rect 16604 21362 16660 21374
rect 16604 21310 16606 21362
rect 16658 21310 16660 21362
rect 16604 20804 16660 21310
rect 15820 20132 16100 20188
rect 15260 19854 15262 19906
rect 15314 19854 15316 19906
rect 15260 19842 15316 19854
rect 15708 18564 15764 18574
rect 14700 18386 14756 18396
rect 14924 18452 14980 18462
rect 15372 18452 15428 18462
rect 14924 18450 15372 18452
rect 14924 18398 14926 18450
rect 14978 18398 15372 18450
rect 14924 18396 15372 18398
rect 14924 18386 14980 18396
rect 15372 18358 15428 18396
rect 14140 18228 14196 18238
rect 14140 17220 14196 18172
rect 13132 17054 13134 17106
rect 13186 17054 13188 17106
rect 13132 16772 13188 17054
rect 13692 17164 14196 17220
rect 13356 16884 13412 16894
rect 13356 16790 13412 16828
rect 13692 16882 13748 17164
rect 13804 16996 13860 17006
rect 13804 16902 13860 16940
rect 14028 16994 14084 17006
rect 14028 16942 14030 16994
rect 14082 16942 14084 16994
rect 13692 16830 13694 16882
rect 13746 16830 13748 16882
rect 13692 16818 13748 16830
rect 14028 16884 14084 16942
rect 14140 16994 14196 17164
rect 14140 16942 14142 16994
rect 14194 16942 14196 16994
rect 14140 16930 14196 16942
rect 14028 16818 14084 16828
rect 15708 16882 15764 18508
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15708 16818 15764 16830
rect 15820 17442 15876 17454
rect 15820 17390 15822 17442
rect 15874 17390 15876 17442
rect 15820 16884 15876 17390
rect 16044 17108 16100 20132
rect 16156 19906 16212 19918
rect 16156 19854 16158 19906
rect 16210 19854 16212 19906
rect 16156 18564 16212 19854
rect 16268 19234 16324 19246
rect 16268 19182 16270 19234
rect 16322 19182 16324 19234
rect 16268 19012 16324 19182
rect 16492 19124 16548 19134
rect 16268 18946 16324 18956
rect 16380 19122 16548 19124
rect 16380 19070 16494 19122
rect 16546 19070 16548 19122
rect 16380 19068 16548 19070
rect 16156 18470 16212 18508
rect 16156 18340 16212 18350
rect 16156 17666 16212 18284
rect 16156 17614 16158 17666
rect 16210 17614 16212 17666
rect 16156 17602 16212 17614
rect 16044 17052 16324 17108
rect 16156 16884 16212 16894
rect 15820 16828 16156 16884
rect 16156 16790 16212 16828
rect 13020 16658 13076 16670
rect 13020 16606 13022 16658
rect 13074 16606 13076 16658
rect 13020 16212 13076 16606
rect 13020 16146 13076 16156
rect 13132 16100 13188 16716
rect 13132 16034 13188 16044
rect 15820 15986 15876 15998
rect 15820 15934 15822 15986
rect 15874 15934 15876 15986
rect 14588 15876 14644 15886
rect 12908 15708 13188 15764
rect 12908 15540 12964 15550
rect 12796 15538 13076 15540
rect 12796 15486 12910 15538
rect 12962 15486 13076 15538
rect 12796 15484 13076 15486
rect 12908 15474 12964 15484
rect 12012 15092 12404 15148
rect 11676 14366 11678 14418
rect 11730 14366 11732 14418
rect 11676 14354 11732 14366
rect 11340 13906 11396 13916
rect 11116 13188 11172 13198
rect 11116 13074 11172 13132
rect 11116 13022 11118 13074
rect 11170 13022 11172 13074
rect 11116 13010 11172 13022
rect 11452 12852 11508 12862
rect 11452 12758 11508 12796
rect 11676 12850 11732 12862
rect 11676 12798 11678 12850
rect 11730 12798 11732 12850
rect 11116 12740 11172 12750
rect 11116 12646 11172 12684
rect 11228 12738 11284 12750
rect 11228 12686 11230 12738
rect 11282 12686 11284 12738
rect 11228 12516 11284 12686
rect 10780 12226 10836 12236
rect 11116 12460 11284 12516
rect 11116 12292 11172 12460
rect 11116 12198 11172 12236
rect 11228 12178 11284 12190
rect 11228 12126 11230 12178
rect 11282 12126 11284 12178
rect 11228 11732 11284 12126
rect 11228 11666 11284 11676
rect 11676 11396 11732 12798
rect 11676 11340 12180 11396
rect 10220 11330 10276 11340
rect 9884 10836 9940 10846
rect 9548 10670 9550 10722
rect 9602 10670 9604 10722
rect 9548 10658 9604 10670
rect 9660 10834 9940 10836
rect 9660 10782 9886 10834
rect 9938 10782 9940 10834
rect 9660 10780 9940 10782
rect 7868 10518 7924 10556
rect 8204 10612 8260 10622
rect 8092 9940 8148 9950
rect 8204 9940 8260 10556
rect 8316 10498 8372 10510
rect 8316 10446 8318 10498
rect 8370 10446 8372 10498
rect 8316 10052 8372 10446
rect 8876 10500 8932 10510
rect 8876 10406 8932 10444
rect 8652 10386 8708 10398
rect 8652 10334 8654 10386
rect 8706 10334 8708 10386
rect 8428 10052 8484 10062
rect 8316 10050 8484 10052
rect 8316 9998 8430 10050
rect 8482 9998 8484 10050
rect 8316 9996 8484 9998
rect 8428 9986 8484 9996
rect 8092 9938 8260 9940
rect 8092 9886 8094 9938
rect 8146 9886 8260 9938
rect 8092 9884 8260 9886
rect 8092 9874 8148 9884
rect 7532 9774 7534 9826
rect 7586 9774 7588 9826
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 5628 8372 5684 8382
rect 5628 8278 5684 8316
rect 7532 8372 7588 9774
rect 8652 9714 8708 10334
rect 8652 9662 8654 9714
rect 8706 9662 8708 9714
rect 8652 9650 8708 9662
rect 8764 10388 8820 10398
rect 7532 8306 7588 8316
rect 7756 9604 7812 9614
rect 7756 8370 7812 9548
rect 8540 9604 8596 9614
rect 8540 9510 8596 9548
rect 8764 8372 8820 10332
rect 9100 10388 9156 10398
rect 9660 10388 9716 10780
rect 9884 10770 9940 10780
rect 9996 10834 10052 11116
rect 11788 11172 11844 11182
rect 11788 11078 11844 11116
rect 9996 10782 9998 10834
rect 10050 10782 10052 10834
rect 9996 10770 10052 10782
rect 10220 10836 10276 10846
rect 9100 10386 9716 10388
rect 9100 10334 9102 10386
rect 9154 10334 9716 10386
rect 9100 10332 9716 10334
rect 9772 10610 9828 10622
rect 9772 10558 9774 10610
rect 9826 10558 9828 10610
rect 9100 10322 9156 10332
rect 9772 9492 9828 10558
rect 10220 10610 10276 10780
rect 10668 10836 10724 10846
rect 10668 10742 10724 10780
rect 10220 10558 10222 10610
rect 10274 10558 10276 10610
rect 10220 10546 10276 10558
rect 11900 9492 11956 11340
rect 12124 11284 12180 11340
rect 12124 11190 12180 11228
rect 12348 10836 12404 15092
rect 12908 12066 12964 12078
rect 12908 12014 12910 12066
rect 12962 12014 12964 12066
rect 12796 11620 12852 11630
rect 12572 11618 12852 11620
rect 12572 11566 12798 11618
rect 12850 11566 12852 11618
rect 12572 11564 12852 11566
rect 12460 10836 12516 10846
rect 12348 10834 12516 10836
rect 12348 10782 12462 10834
rect 12514 10782 12516 10834
rect 12348 10780 12516 10782
rect 12236 10610 12292 10622
rect 12236 10558 12238 10610
rect 12290 10558 12292 10610
rect 12236 9826 12292 10558
rect 12460 10500 12516 10780
rect 12572 10722 12628 11564
rect 12796 11554 12852 11564
rect 12572 10670 12574 10722
rect 12626 10670 12628 10722
rect 12572 10658 12628 10670
rect 12684 11284 12740 11294
rect 12684 10724 12740 11228
rect 12460 10444 12628 10500
rect 12236 9774 12238 9826
rect 12290 9774 12292 9826
rect 12236 9762 12292 9774
rect 12460 9828 12516 9838
rect 12460 9734 12516 9772
rect 12012 9716 12068 9726
rect 12012 9714 12180 9716
rect 12012 9662 12014 9714
rect 12066 9662 12180 9714
rect 12012 9660 12180 9662
rect 12012 9650 12068 9660
rect 11900 9436 12068 9492
rect 9772 9426 9828 9436
rect 12012 9044 12068 9436
rect 12124 9268 12180 9660
rect 12348 9604 12404 9614
rect 12348 9602 12516 9604
rect 12348 9550 12350 9602
rect 12402 9550 12516 9602
rect 12348 9548 12516 9550
rect 12348 9538 12404 9548
rect 12236 9268 12292 9278
rect 12124 9266 12292 9268
rect 12124 9214 12238 9266
rect 12290 9214 12292 9266
rect 12124 9212 12292 9214
rect 12236 9202 12292 9212
rect 12348 9268 12404 9278
rect 12348 9174 12404 9212
rect 12124 9044 12180 9054
rect 12012 9042 12180 9044
rect 12012 8990 12126 9042
rect 12178 8990 12180 9042
rect 12012 8988 12180 8990
rect 12124 8978 12180 8988
rect 12460 8428 12516 9548
rect 9100 8372 9156 8382
rect 7756 8318 7758 8370
rect 7810 8318 7812 8370
rect 7756 8306 7812 8318
rect 8540 8370 9156 8372
rect 8540 8318 9102 8370
rect 9154 8318 9156 8370
rect 8540 8316 9156 8318
rect 8540 8258 8596 8316
rect 9100 8306 9156 8316
rect 11788 8372 12516 8428
rect 8540 8206 8542 8258
rect 8594 8206 8596 8258
rect 8540 8194 8596 8206
rect 9660 7588 9716 7598
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 9660 6802 9716 7532
rect 9660 6750 9662 6802
rect 9714 6750 9716 6802
rect 9660 6738 9716 6750
rect 11788 6690 11844 8372
rect 12572 7588 12628 10444
rect 12684 9938 12740 10668
rect 12908 11172 12964 12014
rect 12908 10612 12964 11116
rect 13020 11618 13076 15484
rect 13132 12402 13188 15708
rect 14588 14418 14644 15820
rect 15260 15204 15316 15214
rect 14924 14532 14980 14542
rect 14924 14438 14980 14476
rect 14588 14366 14590 14418
rect 14642 14366 14644 14418
rect 14588 14354 14644 14366
rect 15260 14306 15316 15148
rect 15484 14532 15540 14542
rect 15484 14438 15540 14476
rect 15260 14254 15262 14306
rect 15314 14254 15316 14306
rect 14812 13972 14868 13982
rect 14812 13878 14868 13916
rect 13132 12350 13134 12402
rect 13186 12350 13188 12402
rect 13132 12338 13188 12350
rect 15148 13634 15204 13646
rect 15148 13582 15150 13634
rect 15202 13582 15204 13634
rect 13020 11566 13022 11618
rect 13074 11566 13076 11618
rect 13020 10834 13076 11566
rect 13020 10782 13022 10834
rect 13074 10782 13076 10834
rect 13020 10770 13076 10782
rect 13692 12066 13748 12078
rect 13692 12014 13694 12066
rect 13746 12014 13748 12066
rect 13580 10724 13636 10734
rect 13580 10630 13636 10668
rect 13692 10724 13748 12014
rect 13916 10724 13972 10734
rect 13692 10668 13916 10724
rect 12908 10546 12964 10556
rect 12684 9886 12686 9938
rect 12738 9886 12740 9938
rect 12684 9874 12740 9886
rect 12908 10388 12964 10398
rect 12908 9826 12964 10332
rect 13692 10388 13748 10668
rect 13916 10610 13972 10668
rect 13916 10558 13918 10610
rect 13970 10558 13972 10610
rect 13916 10546 13972 10558
rect 14364 10500 14420 10510
rect 13692 10322 13748 10332
rect 13916 10386 13972 10398
rect 13916 10334 13918 10386
rect 13970 10334 13972 10386
rect 12908 9774 12910 9826
rect 12962 9774 12964 9826
rect 12796 9492 12852 9502
rect 12796 9042 12852 9436
rect 12908 9268 12964 9774
rect 12908 9202 12964 9212
rect 13580 9828 13636 9838
rect 13580 9602 13636 9772
rect 13916 9828 13972 10334
rect 13916 9762 13972 9772
rect 14364 9826 14420 10444
rect 15148 10052 15204 13582
rect 15260 12180 15316 14254
rect 15596 13972 15652 13982
rect 15596 13878 15652 13916
rect 15260 12124 15764 12180
rect 15260 10500 15316 10510
rect 15260 10406 15316 10444
rect 14924 9996 15204 10052
rect 14924 9940 14980 9996
rect 14364 9774 14366 9826
rect 14418 9774 14420 9826
rect 14364 9762 14420 9774
rect 14700 9884 14980 9940
rect 13580 9550 13582 9602
rect 13634 9550 13636 9602
rect 13580 9156 13636 9550
rect 13580 9090 13636 9100
rect 14700 9156 14756 9884
rect 15036 9828 15092 9838
rect 15036 9734 15092 9772
rect 15484 9828 15540 9866
rect 15484 9762 15540 9772
rect 15596 9826 15652 9838
rect 15596 9774 15598 9826
rect 15650 9774 15652 9826
rect 15372 9716 15428 9726
rect 14812 9604 14868 9614
rect 14812 9510 14868 9548
rect 14924 9602 14980 9614
rect 14924 9550 14926 9602
rect 14978 9550 14980 9602
rect 14700 9090 14756 9100
rect 14812 9156 14868 9166
rect 14924 9156 14980 9550
rect 14812 9154 14980 9156
rect 14812 9102 14814 9154
rect 14866 9102 14980 9154
rect 14812 9100 14980 9102
rect 15148 9380 15204 9390
rect 14812 9090 14868 9100
rect 12796 8990 12798 9042
rect 12850 8990 12852 9042
rect 12796 8978 12852 8990
rect 15148 9042 15204 9324
rect 15372 9268 15428 9660
rect 15596 9716 15652 9774
rect 15708 9828 15764 12124
rect 15820 9828 15876 15934
rect 16156 15540 16212 15550
rect 15932 14532 15988 14542
rect 15932 14438 15988 14476
rect 16156 11788 16212 15484
rect 16268 14756 16324 17052
rect 16380 15148 16436 19068
rect 16492 19058 16548 19068
rect 16604 19010 16660 20748
rect 16716 20804 16772 21532
rect 16940 20804 16996 20814
rect 16716 20802 16996 20804
rect 16716 20750 16942 20802
rect 16994 20750 16996 20802
rect 16716 20748 16996 20750
rect 16716 20692 16772 20748
rect 16940 20738 16996 20748
rect 16716 20626 16772 20636
rect 16940 20580 16996 20590
rect 17052 20580 17108 22316
rect 16940 20578 17108 20580
rect 16940 20526 16942 20578
rect 16994 20526 17108 20578
rect 16940 20524 17108 20526
rect 16940 20514 16996 20524
rect 16716 20468 16772 20478
rect 16716 20130 16772 20412
rect 16716 20078 16718 20130
rect 16770 20078 16772 20130
rect 16716 20066 16772 20078
rect 16604 18958 16606 19010
rect 16658 18958 16660 19010
rect 16604 18946 16660 18958
rect 16492 18562 16548 18574
rect 16492 18510 16494 18562
rect 16546 18510 16548 18562
rect 16492 18228 16548 18510
rect 16492 18162 16548 18172
rect 17052 17444 17108 17454
rect 16940 17442 17108 17444
rect 16940 17390 17054 17442
rect 17106 17390 17108 17442
rect 16940 17388 17108 17390
rect 16940 16996 16996 17388
rect 17052 17378 17108 17388
rect 16604 16770 16660 16782
rect 16604 16718 16606 16770
rect 16658 16718 16660 16770
rect 16604 15428 16660 16718
rect 16604 15362 16660 15372
rect 16380 15092 16660 15148
rect 16268 14662 16324 14700
rect 16492 14644 16548 14654
rect 16492 14550 16548 14588
rect 16604 13748 16660 15092
rect 16716 14756 16772 14766
rect 16716 13970 16772 14700
rect 16716 13918 16718 13970
rect 16770 13918 16772 13970
rect 16716 13906 16772 13918
rect 16940 13972 16996 16940
rect 17052 14644 17108 14654
rect 17164 14644 17220 22428
rect 17724 22372 17780 22382
rect 17836 22372 17892 22878
rect 18508 22484 18564 22990
rect 18620 22932 18676 23102
rect 18620 22866 18676 22876
rect 18508 22418 18564 22428
rect 17724 22370 18004 22372
rect 17724 22318 17726 22370
rect 17778 22318 18004 22370
rect 17724 22316 18004 22318
rect 17724 22306 17780 22316
rect 17388 20804 17444 20814
rect 17388 20710 17444 20748
rect 17948 20690 18004 22316
rect 17948 20638 17950 20690
rect 18002 20638 18004 20690
rect 17948 20626 18004 20638
rect 18732 20188 18788 23772
rect 19516 23154 19572 24220
rect 19628 23938 19684 23950
rect 19628 23886 19630 23938
rect 19682 23886 19684 23938
rect 19628 23716 19684 23886
rect 19964 23716 20020 23726
rect 19628 23714 20020 23716
rect 19628 23662 19966 23714
rect 20018 23662 20020 23714
rect 19628 23660 20020 23662
rect 19628 23268 19684 23660
rect 19964 23650 20020 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23268 20244 23278
rect 19628 23266 20244 23268
rect 19628 23214 20190 23266
rect 20242 23214 20244 23266
rect 19628 23212 20244 23214
rect 19516 23102 19518 23154
rect 19570 23102 19572 23154
rect 19516 23090 19572 23102
rect 20188 23044 20244 23212
rect 20188 22978 20244 22988
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20076 21474 20132 21486
rect 20076 21422 20078 21474
rect 20130 21422 20132 21474
rect 20076 20580 20132 21422
rect 20076 20514 20132 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 18620 20132 18788 20188
rect 17276 19124 17332 19134
rect 17276 19030 17332 19068
rect 17276 18452 17332 18462
rect 17276 16212 17332 18396
rect 17724 17556 17780 17566
rect 17388 16996 17444 17006
rect 17612 16996 17668 17006
rect 17388 16902 17444 16940
rect 17500 16940 17612 16996
rect 17276 16098 17332 16156
rect 17276 16046 17278 16098
rect 17330 16046 17332 16098
rect 17276 16034 17332 16046
rect 17388 15428 17444 15438
rect 17388 15334 17444 15372
rect 17052 14642 17220 14644
rect 17052 14590 17054 14642
rect 17106 14590 17220 14642
rect 17052 14588 17220 14590
rect 17052 14578 17108 14588
rect 17164 14532 17220 14588
rect 17164 14466 17220 14476
rect 17388 14308 17444 14318
rect 16940 13906 16996 13916
rect 17164 14306 17444 14308
rect 17164 14254 17390 14306
rect 17442 14254 17444 14306
rect 17164 14252 17444 14254
rect 16604 13692 16772 13748
rect 16156 11732 16324 11788
rect 16268 10836 16324 11732
rect 16268 10742 16324 10780
rect 16604 9828 16660 9838
rect 15820 9772 15988 9828
rect 15708 9762 15764 9772
rect 15596 9650 15652 9660
rect 15708 9602 15764 9614
rect 15708 9550 15710 9602
rect 15762 9550 15764 9602
rect 15708 9380 15764 9550
rect 15820 9602 15876 9614
rect 15820 9550 15822 9602
rect 15874 9550 15876 9602
rect 15820 9492 15876 9550
rect 15820 9426 15876 9436
rect 15708 9314 15764 9324
rect 15596 9268 15652 9278
rect 15372 9212 15596 9268
rect 15596 9154 15652 9212
rect 15596 9102 15598 9154
rect 15650 9102 15652 9154
rect 15596 9090 15652 9102
rect 15708 9154 15764 9166
rect 15708 9102 15710 9154
rect 15762 9102 15764 9154
rect 15148 8990 15150 9042
rect 15202 8990 15204 9042
rect 15148 8978 15204 8990
rect 15708 9044 15764 9102
rect 15932 9156 15988 9772
rect 16380 9826 16660 9828
rect 16380 9774 16606 9826
rect 16658 9774 16660 9826
rect 16380 9772 16660 9774
rect 16044 9716 16100 9726
rect 16380 9716 16436 9772
rect 16604 9762 16660 9772
rect 16044 9714 16436 9716
rect 16044 9662 16046 9714
rect 16098 9662 16436 9714
rect 16044 9660 16436 9662
rect 16044 9650 16100 9660
rect 15932 9100 16212 9156
rect 15708 8978 15764 8988
rect 14924 8930 14980 8942
rect 14924 8878 14926 8930
rect 14978 8878 14980 8930
rect 14924 8428 14980 8878
rect 15708 8820 15764 8830
rect 15708 8726 15764 8764
rect 12572 7522 12628 7532
rect 14252 8372 14980 8428
rect 11788 6638 11790 6690
rect 11842 6638 11844 6690
rect 11788 6626 11844 6638
rect 12572 6690 12628 6702
rect 12572 6638 12574 6690
rect 12626 6638 12628 6690
rect 12572 6468 12628 6638
rect 12572 6402 12628 6412
rect 13580 6468 13636 6478
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 13580 5124 13636 6412
rect 13580 4338 13636 5068
rect 14252 4450 14308 8372
rect 15372 5124 15428 5134
rect 15820 5124 15876 5134
rect 16156 5124 16212 9100
rect 16268 8820 16324 9660
rect 16492 9604 16548 9614
rect 16492 9210 16548 9548
rect 16716 9492 16772 13692
rect 17164 12740 17220 14252
rect 17388 14242 17444 14252
rect 17164 11394 17220 12684
rect 17164 11342 17166 11394
rect 17218 11342 17220 11394
rect 17164 11330 17220 11342
rect 17500 11396 17556 16940
rect 17612 16930 17668 16940
rect 17724 15538 17780 17500
rect 17948 16996 18004 17006
rect 17724 15486 17726 15538
rect 17778 15486 17780 15538
rect 17724 15474 17780 15486
rect 17836 16884 17892 16894
rect 17836 15538 17892 16828
rect 17948 16882 18004 16940
rect 17948 16830 17950 16882
rect 18002 16830 18004 16882
rect 17948 16818 18004 16830
rect 17836 15486 17838 15538
rect 17890 15486 17892 15538
rect 17836 15474 17892 15486
rect 18060 15540 18116 15550
rect 17612 15314 17668 15326
rect 17612 15262 17614 15314
rect 17666 15262 17668 15314
rect 17612 15204 17668 15262
rect 17612 15138 17668 15148
rect 17724 15316 17780 15326
rect 17612 14644 17668 14654
rect 17612 12404 17668 14588
rect 17724 14530 17780 15260
rect 18060 15314 18116 15484
rect 18060 15262 18062 15314
rect 18114 15262 18116 15314
rect 18060 15204 18116 15262
rect 18620 15316 18676 20132
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 18732 18340 18788 18350
rect 18732 18246 18788 18284
rect 19516 18340 19572 18350
rect 19516 17778 19572 18284
rect 20188 17780 20244 17790
rect 20300 17780 20356 28700
rect 21308 28756 21364 28766
rect 21308 28642 21364 28700
rect 21980 28756 22036 28766
rect 21308 28590 21310 28642
rect 21362 28590 21364 28642
rect 21308 28578 21364 28590
rect 21532 28644 21588 28654
rect 21532 28550 21588 28588
rect 21980 28642 22036 28700
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21980 28578 22036 28590
rect 22316 28644 22372 28654
rect 22316 28550 22372 28588
rect 21756 28418 21812 28430
rect 21756 28366 21758 28418
rect 21810 28366 21812 28418
rect 21756 27972 21812 28366
rect 21868 27972 21924 27982
rect 21756 27970 21924 27972
rect 21756 27918 21870 27970
rect 21922 27918 21924 27970
rect 21756 27916 21924 27918
rect 21868 27906 21924 27916
rect 21644 26516 21700 26526
rect 21644 25506 21700 26460
rect 21644 25454 21646 25506
rect 21698 25454 21700 25506
rect 21644 25442 21700 25454
rect 21308 25396 21364 25406
rect 21196 25394 21364 25396
rect 21196 25342 21310 25394
rect 21362 25342 21364 25394
rect 21196 25340 21364 25342
rect 20860 24948 20916 24958
rect 20860 24388 20916 24892
rect 20860 24050 20916 24332
rect 20860 23998 20862 24050
rect 20914 23998 20916 24050
rect 20860 23986 20916 23998
rect 21196 24052 21252 25340
rect 21308 25330 21364 25340
rect 21420 25396 21476 25406
rect 22540 25396 22596 30268
rect 23436 29764 23492 31388
rect 22988 29708 23492 29764
rect 22988 29650 23044 29708
rect 22988 29598 22990 29650
rect 23042 29598 23044 29650
rect 22988 29586 23044 29598
rect 23212 29540 23268 29550
rect 23100 29538 23268 29540
rect 23100 29486 23214 29538
rect 23266 29486 23268 29538
rect 23100 29484 23268 29486
rect 22988 28756 23044 28766
rect 22876 28700 22988 28756
rect 22652 28084 22708 28094
rect 22652 27858 22708 28028
rect 22876 28082 22932 28700
rect 22988 28690 23044 28700
rect 23100 28644 23156 29484
rect 23212 29474 23268 29484
rect 23436 29426 23492 29708
rect 24108 29650 24164 31500
rect 25564 31556 25620 31566
rect 25564 31462 25620 31500
rect 24108 29598 24110 29650
rect 24162 29598 24164 29650
rect 24108 29586 24164 29598
rect 23436 29374 23438 29426
rect 23490 29374 23492 29426
rect 23436 29362 23492 29374
rect 23996 29314 24052 29326
rect 23996 29262 23998 29314
rect 24050 29262 24052 29314
rect 23100 28578 23156 28588
rect 23212 28980 23268 28990
rect 22876 28030 22878 28082
rect 22930 28030 22932 28082
rect 22876 28018 22932 28030
rect 22652 27806 22654 27858
rect 22706 27806 22708 27858
rect 22652 27794 22708 27806
rect 23100 27970 23156 27982
rect 23100 27918 23102 27970
rect 23154 27918 23156 27970
rect 22652 26852 22708 26862
rect 22652 25620 22708 26796
rect 23100 26516 23156 27918
rect 23212 27970 23268 28924
rect 23996 28756 24052 29262
rect 23996 28690 24052 28700
rect 26012 28868 26068 28878
rect 23660 28084 23716 28094
rect 23660 27990 23716 28028
rect 25340 28084 25396 28094
rect 23212 27918 23214 27970
rect 23266 27918 23268 27970
rect 23212 27906 23268 27918
rect 25340 27858 25396 28028
rect 26012 27970 26068 28812
rect 26012 27918 26014 27970
rect 26066 27918 26068 27970
rect 26012 27906 26068 27918
rect 25340 27806 25342 27858
rect 25394 27806 25396 27858
rect 25340 27794 25396 27806
rect 23100 26450 23156 26460
rect 23884 26852 23940 26862
rect 23100 25620 23156 25630
rect 22652 25618 23156 25620
rect 22652 25566 22654 25618
rect 22706 25566 23102 25618
rect 23154 25566 23156 25618
rect 22652 25564 23156 25566
rect 22652 25554 22708 25564
rect 23100 25508 23156 25564
rect 23100 25442 23156 25452
rect 23772 25508 23828 25518
rect 23772 25414 23828 25452
rect 23884 25396 23940 26796
rect 26124 26852 26180 31614
rect 26460 31668 26516 31678
rect 26460 31574 26516 31612
rect 26236 28980 26292 28990
rect 26236 28530 26292 28924
rect 27020 28756 27076 32060
rect 27132 31890 27188 32956
rect 27132 31838 27134 31890
rect 27186 31838 27188 31890
rect 27132 31668 27188 31838
rect 27132 31602 27188 31612
rect 26572 28754 27076 28756
rect 26572 28702 27022 28754
rect 27074 28702 27076 28754
rect 26572 28700 27076 28702
rect 26572 28642 26628 28700
rect 27020 28690 27076 28700
rect 26572 28590 26574 28642
rect 26626 28590 26628 28642
rect 26572 28578 26628 28590
rect 26236 28478 26238 28530
rect 26290 28478 26292 28530
rect 26236 28466 26292 28478
rect 26124 26786 26180 26796
rect 26012 25844 26068 25854
rect 25228 25620 25284 25630
rect 25228 25526 25284 25564
rect 24220 25508 24276 25518
rect 24220 25414 24276 25452
rect 24892 25506 24948 25518
rect 24892 25454 24894 25506
rect 24946 25454 24948 25506
rect 22540 25340 22820 25396
rect 21420 25302 21476 25340
rect 22316 24724 22372 24734
rect 22092 24612 22148 24622
rect 21532 24388 21588 24398
rect 21532 24162 21588 24332
rect 21532 24110 21534 24162
rect 21586 24110 21588 24162
rect 21532 24098 21588 24110
rect 21196 23986 21252 23996
rect 21532 23940 21588 23950
rect 21532 23846 21588 23884
rect 22092 23938 22148 24556
rect 22092 23886 22094 23938
rect 22146 23886 22148 23938
rect 22092 23874 22148 23886
rect 21868 23828 21924 23838
rect 21196 23044 21252 23054
rect 21196 22950 21252 22988
rect 21532 22372 21588 22382
rect 21756 22372 21812 22382
rect 21532 22370 21812 22372
rect 21532 22318 21534 22370
rect 21586 22318 21758 22370
rect 21810 22318 21812 22370
rect 21532 22316 21812 22318
rect 21532 22148 21588 22316
rect 21756 22306 21812 22316
rect 21532 22082 21588 22092
rect 21644 18452 21700 18462
rect 21644 18358 21700 18396
rect 20860 18340 20916 18350
rect 20860 18246 20916 18284
rect 21868 18228 21924 23772
rect 21980 23714 22036 23726
rect 21980 23662 21982 23714
rect 22034 23662 22036 23714
rect 21980 21700 22036 23662
rect 22204 21700 22260 21710
rect 21980 21698 22260 21700
rect 21980 21646 22206 21698
rect 22258 21646 22260 21698
rect 21980 21644 22260 21646
rect 22204 21634 22260 21644
rect 22316 20188 22372 24668
rect 22428 24612 22484 24622
rect 22428 23938 22484 24556
rect 22428 23886 22430 23938
rect 22482 23886 22484 23938
rect 22428 23874 22484 23886
rect 22540 23940 22596 23950
rect 22540 23846 22596 23884
rect 22652 23828 22708 23838
rect 22652 23734 22708 23772
rect 22764 20188 22820 25340
rect 23436 25284 23492 25294
rect 23100 25228 23436 25284
rect 23100 23938 23156 25228
rect 23436 25190 23492 25228
rect 23884 24834 23940 25340
rect 24444 25282 24500 25294
rect 24444 25230 24446 25282
rect 24498 25230 24500 25282
rect 24444 24948 24500 25230
rect 24892 25284 24948 25454
rect 26012 25394 26068 25788
rect 26012 25342 26014 25394
rect 26066 25342 26068 25394
rect 26012 25330 26068 25342
rect 24892 25218 24948 25228
rect 25564 25284 25620 25294
rect 25676 25284 25732 25294
rect 25620 25282 25732 25284
rect 25620 25230 25678 25282
rect 25730 25230 25732 25282
rect 25620 25228 25732 25230
rect 24444 24882 24500 24892
rect 25340 24948 25396 24958
rect 25340 24854 25396 24892
rect 23884 24782 23886 24834
rect 23938 24782 23940 24834
rect 23884 24770 23940 24782
rect 24220 24722 24276 24734
rect 24220 24670 24222 24722
rect 24274 24670 24276 24722
rect 23996 24612 24052 24622
rect 24220 24612 24276 24670
rect 24668 24612 24724 24622
rect 24220 24610 24724 24612
rect 24220 24558 24670 24610
rect 24722 24558 24724 24610
rect 24220 24556 24724 24558
rect 23996 24518 24052 24556
rect 24668 24500 24724 24556
rect 24668 24434 24724 24444
rect 23100 23886 23102 23938
rect 23154 23886 23156 23938
rect 23100 23874 23156 23886
rect 25452 23940 25508 23950
rect 25452 23846 25508 23884
rect 22988 21586 23044 21598
rect 22988 21534 22990 21586
rect 23042 21534 23044 21586
rect 22988 20244 23044 21534
rect 23548 21474 23604 21486
rect 23548 21422 23550 21474
rect 23602 21422 23604 21474
rect 23100 20244 23156 20254
rect 22988 20188 23100 20244
rect 21868 18162 21924 18172
rect 21980 20132 22372 20188
rect 22652 20132 22932 20188
rect 19516 17726 19518 17778
rect 19570 17726 19572 17778
rect 19516 17714 19572 17726
rect 19740 17778 20356 17780
rect 19740 17726 20190 17778
rect 20242 17726 20356 17778
rect 19740 17724 20356 17726
rect 19740 17666 19796 17724
rect 20188 17686 20244 17724
rect 19740 17614 19742 17666
rect 19794 17614 19796 17666
rect 19740 17602 19796 17614
rect 19404 17556 19460 17566
rect 19404 17462 19460 17500
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20300 16884 20356 17724
rect 20300 16818 20356 16828
rect 19292 16212 19348 16222
rect 19292 15876 19348 16156
rect 19292 15810 19348 15820
rect 20860 15988 20916 15998
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19516 15540 19572 15550
rect 19516 15446 19572 15484
rect 20860 15538 20916 15932
rect 20860 15486 20862 15538
rect 20914 15486 20916 15538
rect 18844 15428 18900 15438
rect 18844 15334 18900 15372
rect 19964 15428 20020 15438
rect 19964 15334 20020 15372
rect 18620 15222 18676 15260
rect 19180 15314 19236 15326
rect 19180 15262 19182 15314
rect 19234 15262 19236 15314
rect 19180 15148 19236 15262
rect 18060 15138 18116 15148
rect 18844 15092 19236 15148
rect 20412 15204 20468 15214
rect 20412 15110 20468 15148
rect 19292 15092 19348 15102
rect 18060 14644 18116 14654
rect 18060 14550 18116 14588
rect 18844 14642 18900 15092
rect 18844 14590 18846 14642
rect 18898 14590 18900 14642
rect 17724 14478 17726 14530
rect 17778 14478 17780 14530
rect 17724 14466 17780 14478
rect 18172 14532 18228 14542
rect 18172 14438 18228 14476
rect 18844 14532 18900 14590
rect 19292 14642 19348 15036
rect 19292 14590 19294 14642
rect 19346 14590 19348 14642
rect 19292 14578 19348 14590
rect 18844 14466 18900 14476
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 17612 12348 17780 12404
rect 17500 11340 17668 11396
rect 17276 11170 17332 11182
rect 17276 11118 17278 11170
rect 17330 11118 17332 11170
rect 17276 10386 17332 11118
rect 17276 10334 17278 10386
rect 17330 10334 17332 10386
rect 17276 10322 17332 10334
rect 17388 11170 17444 11182
rect 17388 11118 17390 11170
rect 17442 11118 17444 11170
rect 17164 10052 17220 10062
rect 17388 10052 17444 11118
rect 17500 11170 17556 11182
rect 17500 11118 17502 11170
rect 17554 11118 17556 11170
rect 17500 10276 17556 11118
rect 17612 10834 17668 11340
rect 17612 10782 17614 10834
rect 17666 10782 17668 10834
rect 17612 10500 17668 10782
rect 17724 11394 17780 12348
rect 17724 11342 17726 11394
rect 17778 11342 17780 11394
rect 17724 10836 17780 11342
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20860 10948 20916 15486
rect 21084 15428 21140 15438
rect 21084 15314 21140 15372
rect 21084 15262 21086 15314
rect 21138 15262 21140 15314
rect 21084 15250 21140 15262
rect 21532 15428 21588 15438
rect 21532 13858 21588 15372
rect 21868 15428 21924 15438
rect 21868 15334 21924 15372
rect 21868 15204 21924 15214
rect 21532 13806 21534 13858
rect 21586 13806 21588 13858
rect 21532 13794 21588 13806
rect 21644 13860 21700 13870
rect 21644 13858 21812 13860
rect 21644 13806 21646 13858
rect 21698 13806 21812 13858
rect 21644 13804 21812 13806
rect 21644 13794 21700 13804
rect 21644 13522 21700 13534
rect 21644 13470 21646 13522
rect 21698 13470 21700 13522
rect 21420 12964 21476 12974
rect 21308 12908 21420 12964
rect 21308 12290 21364 12908
rect 21420 12898 21476 12908
rect 21644 12850 21700 13470
rect 21644 12798 21646 12850
rect 21698 12798 21700 12850
rect 21644 12786 21700 12798
rect 21756 12852 21812 13804
rect 21756 12786 21812 12796
rect 21868 12962 21924 15148
rect 21868 12910 21870 12962
rect 21922 12910 21924 12962
rect 21868 12628 21924 12910
rect 21980 12964 22036 20132
rect 22652 20130 22708 20132
rect 22652 20078 22654 20130
rect 22706 20078 22708 20130
rect 22652 20066 22708 20078
rect 22876 20018 22932 20132
rect 22876 19966 22878 20018
rect 22930 19966 22932 20018
rect 22876 19954 22932 19966
rect 22876 19796 22932 19806
rect 22876 19702 22932 19740
rect 22988 19236 23044 19246
rect 23100 19236 23156 20188
rect 23548 20244 23604 21422
rect 23548 20178 23604 20188
rect 22988 19234 23156 19236
rect 22988 19182 22990 19234
rect 23042 19182 23156 19234
rect 22988 19180 23156 19182
rect 23212 19794 23268 19806
rect 23212 19742 23214 19794
rect 23266 19742 23268 19794
rect 22092 18452 22148 18462
rect 22092 18358 22148 18396
rect 22988 18452 23044 19180
rect 22988 18386 23044 18396
rect 23212 16210 23268 19742
rect 23660 19796 23716 19806
rect 23660 19346 23716 19740
rect 23660 19294 23662 19346
rect 23714 19294 23716 19346
rect 23660 19282 23716 19294
rect 23212 16158 23214 16210
rect 23266 16158 23268 16210
rect 23212 16146 23268 16158
rect 24220 16772 24276 16782
rect 24220 16210 24276 16716
rect 25564 16212 25620 25228
rect 25676 25218 25732 25228
rect 26236 24948 26292 24958
rect 26012 24892 26236 24948
rect 25900 24724 25956 24734
rect 25900 24630 25956 24668
rect 26012 23938 26068 24892
rect 26236 24854 26292 24892
rect 27132 24948 27188 24958
rect 27132 24854 27188 24892
rect 26684 24836 26740 24846
rect 26684 24610 26740 24780
rect 26684 24558 26686 24610
rect 26738 24558 26740 24610
rect 26684 24546 26740 24558
rect 27468 24612 27524 33068
rect 27580 31892 27636 31902
rect 27580 31798 27636 31836
rect 28252 31892 28308 36428
rect 29484 36390 29540 36428
rect 29148 36372 29204 36382
rect 29148 36278 29204 36316
rect 28364 36260 28420 36270
rect 28364 33012 28420 36204
rect 30268 34916 30324 37324
rect 30828 37380 30884 37390
rect 30828 37286 30884 37324
rect 31724 37380 31780 40348
rect 31836 40338 31892 40348
rect 33404 40404 33460 40414
rect 33404 40310 33460 40348
rect 34972 40292 35028 40302
rect 34412 39732 34468 39742
rect 34972 39732 35028 40236
rect 36316 40290 36372 41918
rect 37324 41860 37380 41870
rect 37324 41766 37380 41804
rect 39900 41860 39956 45200
rect 39900 41794 39956 41804
rect 40124 41970 40180 41982
rect 40124 41918 40126 41970
rect 40178 41918 40180 41970
rect 39788 40964 39844 40974
rect 40124 40964 40180 41918
rect 41132 41860 41188 41870
rect 41132 41766 41188 41804
rect 43596 41300 43652 41310
rect 43708 41300 43764 45200
rect 43596 41298 43764 41300
rect 43596 41246 43598 41298
rect 43650 41246 43764 41298
rect 43596 41244 43764 41246
rect 43596 41234 43652 41244
rect 39788 40962 40180 40964
rect 39788 40910 39790 40962
rect 39842 40910 40180 40962
rect 39788 40908 40180 40910
rect 41580 41186 41636 41198
rect 41580 41134 41582 41186
rect 41634 41134 41636 41186
rect 36316 40238 36318 40290
rect 36370 40238 36372 40290
rect 36316 40226 36372 40238
rect 36876 40402 36932 40414
rect 36876 40350 36878 40402
rect 36930 40350 36932 40402
rect 36876 40292 36932 40350
rect 36876 40226 36932 40236
rect 37996 40292 38052 40302
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 32172 39508 32228 39518
rect 31724 37314 31780 37324
rect 31836 39506 32228 39508
rect 31836 39454 32174 39506
rect 32226 39454 32228 39506
rect 31836 39452 32228 39454
rect 30380 37154 30436 37166
rect 30380 37102 30382 37154
rect 30434 37102 30436 37154
rect 30380 36596 30436 37102
rect 30380 36530 30436 36540
rect 30828 36484 30884 36494
rect 30828 36390 30884 36428
rect 31276 36482 31332 36494
rect 31276 36430 31278 36482
rect 31330 36430 31332 36482
rect 30380 36370 30436 36382
rect 30380 36318 30382 36370
rect 30434 36318 30436 36370
rect 30380 35812 30436 36318
rect 30380 35746 30436 35756
rect 30268 34822 30324 34860
rect 30940 34804 30996 34814
rect 30828 34802 30996 34804
rect 30828 34750 30942 34802
rect 30994 34750 30996 34802
rect 30828 34748 30996 34750
rect 30828 33570 30884 34748
rect 30940 34738 30996 34748
rect 31276 34356 31332 36430
rect 31836 35476 31892 39452
rect 32172 39442 32228 39452
rect 31276 34290 31332 34300
rect 31724 35420 31892 35476
rect 30828 33518 30830 33570
rect 30882 33518 30884 33570
rect 30828 33506 30884 33518
rect 31612 34244 31668 34254
rect 30940 33348 30996 33358
rect 31388 33348 31444 33358
rect 30940 33346 31444 33348
rect 30940 33294 30942 33346
rect 30994 33294 31390 33346
rect 31442 33294 31444 33346
rect 30940 33292 31444 33294
rect 30940 33282 30996 33292
rect 31388 33282 31444 33292
rect 28364 32946 28420 32956
rect 30716 33234 30772 33246
rect 30716 33182 30718 33234
rect 30770 33182 30772 33234
rect 30716 32788 30772 33182
rect 31612 33236 31668 34188
rect 31724 34020 31780 35420
rect 33068 35026 33124 35038
rect 33068 34974 33070 35026
rect 33122 34974 33124 35026
rect 32060 34356 32116 34366
rect 31836 34244 31892 34254
rect 31836 34150 31892 34188
rect 32060 34130 32116 34300
rect 33068 34356 33124 34974
rect 33068 34290 33124 34300
rect 33516 34916 33572 34926
rect 32060 34078 32062 34130
rect 32114 34078 32116 34130
rect 32060 34066 32116 34078
rect 31724 33964 31892 34020
rect 31612 33142 31668 33180
rect 31724 33234 31780 33246
rect 31724 33182 31726 33234
rect 31778 33182 31780 33234
rect 31164 33122 31220 33134
rect 31164 33070 31166 33122
rect 31218 33070 31220 33122
rect 31164 33012 31220 33070
rect 30940 32956 31556 33012
rect 30828 32788 30884 32798
rect 30716 32786 30884 32788
rect 30716 32734 30830 32786
rect 30882 32734 30884 32786
rect 30716 32732 30884 32734
rect 30828 32722 30884 32732
rect 30268 32564 30324 32574
rect 30940 32564 30996 32956
rect 31052 32788 31108 32798
rect 31052 32694 31108 32732
rect 31500 32786 31556 32956
rect 31724 32788 31780 33182
rect 31500 32734 31502 32786
rect 31554 32734 31556 32786
rect 31500 32722 31556 32734
rect 31612 32732 31780 32788
rect 28252 31826 28308 31836
rect 30044 32452 30100 32462
rect 30044 31778 30100 32396
rect 30044 31726 30046 31778
rect 30098 31726 30100 31778
rect 30044 31556 30100 31726
rect 30044 31490 30100 31500
rect 30268 31554 30324 32508
rect 30828 32508 30996 32564
rect 31164 32562 31220 32574
rect 31164 32510 31166 32562
rect 31218 32510 31220 32562
rect 30828 32004 30884 32508
rect 30268 31502 30270 31554
rect 30322 31502 30324 31554
rect 30156 30996 30212 31006
rect 30268 30996 30324 31502
rect 30716 31556 30772 31566
rect 30716 31462 30772 31500
rect 30716 31108 30772 31118
rect 30716 31014 30772 31052
rect 30604 30996 30660 31006
rect 30268 30994 30660 30996
rect 30268 30942 30606 30994
rect 30658 30942 30660 30994
rect 30268 30940 30660 30942
rect 28588 30884 28644 30894
rect 28588 30324 28644 30828
rect 28588 30210 28644 30268
rect 30156 30324 30212 30940
rect 28588 30158 28590 30210
rect 28642 30158 28644 30210
rect 28588 28644 28644 30158
rect 29708 30212 29764 30222
rect 28812 30100 28868 30110
rect 28812 29426 28868 30044
rect 28812 29374 28814 29426
rect 28866 29374 28868 29426
rect 28588 28588 28756 28644
rect 28588 28418 28644 28430
rect 28588 28366 28590 28418
rect 28642 28366 28644 28418
rect 28588 28308 28644 28366
rect 28476 28252 28644 28308
rect 28476 27860 28532 28252
rect 28588 28084 28644 28094
rect 28588 27990 28644 28028
rect 28588 27860 28644 27870
rect 28476 27804 28588 27860
rect 28588 27794 28644 27804
rect 28140 27748 28196 27758
rect 28140 27654 28196 27692
rect 28700 26908 28756 28588
rect 28812 28084 28868 29374
rect 29484 29316 29540 29326
rect 29484 29222 29540 29260
rect 29260 28868 29316 28878
rect 29260 28866 29652 28868
rect 29260 28814 29262 28866
rect 29314 28814 29652 28866
rect 29260 28812 29652 28814
rect 29260 28802 29316 28812
rect 29596 28642 29652 28812
rect 29596 28590 29598 28642
rect 29650 28590 29652 28642
rect 29596 28578 29652 28590
rect 29372 28532 29428 28542
rect 29372 28530 29540 28532
rect 29372 28478 29374 28530
rect 29426 28478 29540 28530
rect 29372 28476 29540 28478
rect 29372 28466 29428 28476
rect 29260 28418 29316 28430
rect 29260 28366 29262 28418
rect 29314 28366 29316 28418
rect 29260 28196 29316 28366
rect 29484 28420 29540 28476
rect 29708 28420 29764 30156
rect 30156 30210 30212 30268
rect 30156 30158 30158 30210
rect 30210 30158 30212 30210
rect 30156 30146 30212 30158
rect 30604 30212 30660 30940
rect 30604 30146 30660 30156
rect 30828 29988 30884 31948
rect 30604 29932 30884 29988
rect 30940 30994 30996 31006
rect 30940 30942 30942 30994
rect 30994 30942 30996 30994
rect 30380 29316 30436 29326
rect 29820 28868 29876 28878
rect 29820 28774 29876 28812
rect 30380 28866 30436 29260
rect 30380 28814 30382 28866
rect 30434 28814 30436 28866
rect 30380 28802 30436 28814
rect 29932 28644 29988 28654
rect 29932 28530 29988 28588
rect 29932 28478 29934 28530
rect 29986 28478 29988 28530
rect 29932 28466 29988 28478
rect 29484 28364 29764 28420
rect 30156 28420 30212 28430
rect 30492 28420 30548 28430
rect 30156 28418 30548 28420
rect 30156 28366 30158 28418
rect 30210 28366 30494 28418
rect 30546 28366 30548 28418
rect 30156 28364 30548 28366
rect 29260 28140 29428 28196
rect 28868 28028 29316 28084
rect 28812 28018 28868 28028
rect 28588 26852 28756 26908
rect 28924 27860 28980 27870
rect 27580 24612 27636 24622
rect 27468 24556 27580 24612
rect 27580 24518 27636 24556
rect 26012 23886 26014 23938
rect 26066 23886 26068 23938
rect 26012 23874 26068 23886
rect 26796 22260 26852 22270
rect 26796 22166 26852 22204
rect 28588 22260 28644 26852
rect 28924 25620 28980 27804
rect 28924 25554 28980 25564
rect 29260 23938 29316 28028
rect 29372 27748 29428 28140
rect 30156 27860 30212 28364
rect 30492 28354 30548 28364
rect 30604 28196 30660 29932
rect 30940 28642 30996 30942
rect 31164 30996 31220 32510
rect 31612 32564 31668 32732
rect 31612 32498 31668 32508
rect 31724 32562 31780 32574
rect 31724 32510 31726 32562
rect 31778 32510 31780 32562
rect 31724 31218 31780 32510
rect 31836 32450 31892 33964
rect 32956 33348 33012 33358
rect 32956 33254 33012 33292
rect 32620 33234 32676 33246
rect 32620 33182 32622 33234
rect 32674 33182 32676 33234
rect 32396 33124 32452 33134
rect 32396 32786 32452 33068
rect 32396 32734 32398 32786
rect 32450 32734 32452 32786
rect 32396 32722 32452 32734
rect 31836 32398 31838 32450
rect 31890 32398 31892 32450
rect 31836 32386 31892 32398
rect 32060 32562 32116 32574
rect 32060 32510 32062 32562
rect 32114 32510 32116 32562
rect 32060 32340 32116 32510
rect 32284 32564 32340 32574
rect 32284 32470 32340 32508
rect 32396 32340 32452 32350
rect 32060 32338 32452 32340
rect 32060 32286 32398 32338
rect 32450 32286 32452 32338
rect 32060 32284 32452 32286
rect 32396 32274 32452 32284
rect 31724 31166 31726 31218
rect 31778 31166 31780 31218
rect 31724 31154 31780 31166
rect 31500 31108 31556 31118
rect 31556 31052 31668 31108
rect 31500 31014 31556 31052
rect 31388 30996 31444 31006
rect 31164 30994 31444 30996
rect 31164 30942 31390 30994
rect 31442 30942 31444 30994
rect 31164 30940 31444 30942
rect 31388 29092 31444 30940
rect 31612 29314 31668 31052
rect 32508 30996 32564 31006
rect 32508 30902 32564 30940
rect 31612 29262 31614 29314
rect 31666 29262 31668 29314
rect 31612 29250 31668 29262
rect 32060 30100 32116 30110
rect 32060 29650 32116 30044
rect 32060 29598 32062 29650
rect 32114 29598 32116 29650
rect 31388 29036 31892 29092
rect 30940 28590 30942 28642
rect 30994 28590 30996 28642
rect 30940 28578 30996 28590
rect 30716 28420 30772 28430
rect 31836 28420 31892 29036
rect 31948 28980 32004 28990
rect 31948 28642 32004 28924
rect 31948 28590 31950 28642
rect 32002 28590 32004 28642
rect 31948 28578 32004 28590
rect 31948 28420 32004 28430
rect 30716 28418 31668 28420
rect 30716 28366 30718 28418
rect 30770 28366 31668 28418
rect 30716 28364 31668 28366
rect 31836 28364 31948 28420
rect 30716 28354 30772 28364
rect 30156 27766 30212 27804
rect 30380 28140 30660 28196
rect 29372 26964 29428 27692
rect 30380 26908 30436 28140
rect 30828 27076 30884 27086
rect 29372 26898 29428 26908
rect 30268 26852 30436 26908
rect 30716 26964 30772 27002
rect 30828 26982 30884 27020
rect 31612 27074 31668 28364
rect 31612 27022 31614 27074
rect 31666 27022 31668 27074
rect 31612 27010 31668 27022
rect 31948 27074 32004 28364
rect 31948 27022 31950 27074
rect 32002 27022 32004 27074
rect 31948 27010 32004 27022
rect 30716 26898 30772 26908
rect 32060 26908 32116 29598
rect 32620 29428 32676 33182
rect 32732 33236 32788 33246
rect 32732 33142 32788 33180
rect 33404 30996 33460 31006
rect 33404 30902 33460 30940
rect 33516 30100 33572 34860
rect 34412 33124 34468 39676
rect 34636 39730 35028 39732
rect 34636 39678 34974 39730
rect 35026 39678 35028 39730
rect 34636 39676 35028 39678
rect 34636 37266 34692 39676
rect 34972 39666 35028 39676
rect 37996 39730 38052 40236
rect 39788 40180 39844 40908
rect 39788 40114 39844 40124
rect 37996 39678 37998 39730
rect 38050 39678 38052 39730
rect 37996 39060 38052 39678
rect 37660 39004 37996 39060
rect 37660 38668 37716 39004
rect 37996 38994 38052 39004
rect 38332 39730 38388 39742
rect 38332 39678 38334 39730
rect 38386 39678 38388 39730
rect 37548 38612 37716 38668
rect 38332 38948 38388 39678
rect 41580 39732 41636 41134
rect 41580 39666 41636 39676
rect 40348 39620 40404 39630
rect 39228 39060 39284 39070
rect 39228 38966 39284 39004
rect 40348 39058 40404 39564
rect 41132 39618 41188 39630
rect 41132 39566 41134 39618
rect 41186 39566 41188 39618
rect 40460 39508 40516 39518
rect 40460 39414 40516 39452
rect 40348 39006 40350 39058
rect 40402 39006 40404 39058
rect 40348 38994 40404 39006
rect 41132 39060 41188 39566
rect 41468 39620 41524 39630
rect 41468 39526 41524 39564
rect 41804 39618 41860 39630
rect 41804 39566 41806 39618
rect 41858 39566 41860 39618
rect 41692 39508 41748 39518
rect 41692 39414 41748 39452
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34636 37214 34638 37266
rect 34690 37214 34692 37266
rect 34636 37202 34692 37214
rect 35308 37156 35364 37166
rect 35308 37154 35924 37156
rect 35308 37102 35310 37154
rect 35362 37102 35924 37154
rect 35308 37100 35924 37102
rect 35308 37090 35364 37100
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35532 34018 35588 34030
rect 35532 33966 35534 34018
rect 35586 33966 35588 34018
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34412 33058 34468 33068
rect 34748 33124 34804 33134
rect 35084 33124 35140 33134
rect 34748 33122 35140 33124
rect 34748 33070 34750 33122
rect 34802 33070 35086 33122
rect 35138 33070 35140 33122
rect 34748 33068 35140 33070
rect 34748 32116 34804 33068
rect 35084 33058 35140 33068
rect 35420 33122 35476 33134
rect 35420 33070 35422 33122
rect 35474 33070 35476 33122
rect 35420 33012 35476 33070
rect 35420 32946 35476 32956
rect 35532 32788 35588 33966
rect 35868 33458 35924 37100
rect 37436 37154 37492 37166
rect 37436 37102 37438 37154
rect 37490 37102 37492 37154
rect 37436 37044 37492 37102
rect 37436 36978 37492 36988
rect 37548 36596 37604 38612
rect 37884 38274 37940 38286
rect 37884 38222 37886 38274
rect 37938 38222 37940 38274
rect 37772 37266 37828 37278
rect 37772 37214 37774 37266
rect 37826 37214 37828 37266
rect 37772 37044 37828 37214
rect 37772 36978 37828 36988
rect 37660 36596 37716 36606
rect 37548 36594 37716 36596
rect 37548 36542 37662 36594
rect 37714 36542 37716 36594
rect 37548 36540 37716 36542
rect 35868 33406 35870 33458
rect 35922 33406 35924 33458
rect 35868 33394 35924 33406
rect 36652 35028 36708 35038
rect 36092 33348 36148 33358
rect 36092 33254 36148 33292
rect 35756 33236 35812 33246
rect 35756 33142 35812 33180
rect 36316 33234 36372 33246
rect 36316 33182 36318 33234
rect 36370 33182 36372 33234
rect 36316 32900 36372 33182
rect 36316 32834 36372 32844
rect 35532 32722 35588 32732
rect 35980 32564 36036 32574
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 33516 30006 33572 30044
rect 33628 31556 33684 31566
rect 33628 29876 33684 31500
rect 33628 29810 33684 29820
rect 32284 29372 32900 29428
rect 32284 28530 32340 29372
rect 32732 29204 32788 29214
rect 32508 28644 32564 28654
rect 32508 28550 32564 28588
rect 32284 28478 32286 28530
rect 32338 28478 32340 28530
rect 32284 28466 32340 28478
rect 32732 28530 32788 29148
rect 32732 28478 32734 28530
rect 32786 28478 32788 28530
rect 32732 28466 32788 28478
rect 32844 28642 32900 29372
rect 32844 28590 32846 28642
rect 32898 28590 32900 28642
rect 32844 27076 32900 28590
rect 34636 28980 34692 28990
rect 34636 28644 34692 28924
rect 34636 28550 34692 28588
rect 32844 26908 32900 27020
rect 30492 26852 30548 26862
rect 31836 26852 31892 26862
rect 32060 26852 32228 26908
rect 30268 25844 30324 26852
rect 30492 26850 30660 26852
rect 30492 26798 30494 26850
rect 30546 26798 30660 26850
rect 30492 26796 30660 26798
rect 30492 26786 30548 26796
rect 30604 26068 30660 26796
rect 31836 26758 31892 26796
rect 32060 26180 32116 26190
rect 31948 26124 32060 26180
rect 30604 26012 30884 26068
rect 30324 25788 30660 25844
rect 30268 25750 30324 25788
rect 30492 25620 30548 25630
rect 29932 25618 30548 25620
rect 29932 25566 30494 25618
rect 30546 25566 30548 25618
rect 29932 25564 30548 25566
rect 29932 24050 29988 25564
rect 30492 25554 30548 25564
rect 30604 25506 30660 25788
rect 30604 25454 30606 25506
rect 30658 25454 30660 25506
rect 30604 25442 30660 25454
rect 30828 25506 30884 26012
rect 30828 25454 30830 25506
rect 30882 25454 30884 25506
rect 30828 25442 30884 25454
rect 31052 25282 31108 25294
rect 31052 25230 31054 25282
rect 31106 25230 31108 25282
rect 31052 24276 31108 25230
rect 31276 25282 31332 25294
rect 31276 25230 31278 25282
rect 31330 25230 31332 25282
rect 31276 25060 31332 25230
rect 31276 24722 31332 25004
rect 31948 24834 32004 26124
rect 32060 26114 32116 26124
rect 31948 24782 31950 24834
rect 32002 24782 32004 24834
rect 31948 24770 32004 24782
rect 31276 24670 31278 24722
rect 31330 24670 31332 24722
rect 31276 24658 31332 24670
rect 31612 24722 31668 24734
rect 31612 24670 31614 24722
rect 31666 24670 31668 24722
rect 31500 24612 31556 24622
rect 31500 24518 31556 24556
rect 31612 24276 31668 24670
rect 31052 24220 31668 24276
rect 29932 23998 29934 24050
rect 29986 23998 29988 24050
rect 29932 23986 29988 23998
rect 29260 23886 29262 23938
rect 29314 23886 29316 23938
rect 29260 23874 29316 23886
rect 30156 23940 30212 23950
rect 25788 20244 25844 20254
rect 25788 20020 25844 20188
rect 25788 19926 25844 19964
rect 27132 20020 27188 20030
rect 26572 19906 26628 19918
rect 26572 19854 26574 19906
rect 26626 19854 26628 19906
rect 25788 19346 25844 19358
rect 25788 19294 25790 19346
rect 25842 19294 25844 19346
rect 25788 16436 25844 19294
rect 26572 19346 26628 19854
rect 26684 19796 26740 19806
rect 26684 19458 26740 19740
rect 26684 19406 26686 19458
rect 26738 19406 26740 19458
rect 26684 19394 26740 19406
rect 26572 19294 26574 19346
rect 26626 19294 26628 19346
rect 26572 19282 26628 19294
rect 27132 19348 27188 19964
rect 27132 19254 27188 19292
rect 26348 19234 26404 19246
rect 26348 19182 26350 19234
rect 26402 19182 26404 19234
rect 26012 18340 26068 18350
rect 26348 18340 26404 19182
rect 26012 18338 26404 18340
rect 26012 18286 26014 18338
rect 26066 18286 26404 18338
rect 26012 18284 26404 18286
rect 27244 19124 27300 19134
rect 26012 16884 26068 18284
rect 26012 16818 26068 16828
rect 25788 16380 26180 16436
rect 24220 16158 24222 16210
rect 24274 16158 24276 16210
rect 24220 16100 24276 16158
rect 24444 16156 24724 16212
rect 25564 16156 25844 16212
rect 24444 16100 24500 16156
rect 24220 16034 24276 16044
rect 24332 16044 24500 16100
rect 22428 15988 22484 15998
rect 22428 15538 22484 15932
rect 23324 15988 23380 15998
rect 23324 15894 23380 15932
rect 23548 15986 23604 15998
rect 23548 15934 23550 15986
rect 23602 15934 23604 15986
rect 22988 15874 23044 15886
rect 22988 15822 22990 15874
rect 23042 15822 23044 15874
rect 22988 15540 23044 15822
rect 23100 15876 23156 15886
rect 23100 15874 23268 15876
rect 23100 15822 23102 15874
rect 23154 15822 23268 15874
rect 23100 15820 23268 15822
rect 23100 15810 23156 15820
rect 23100 15540 23156 15550
rect 22428 15486 22430 15538
rect 22482 15486 22484 15538
rect 22428 15474 22484 15486
rect 22652 15538 23156 15540
rect 22652 15486 23102 15538
rect 23154 15486 23156 15538
rect 22652 15484 23156 15486
rect 22092 15316 22148 15326
rect 22652 15316 22708 15484
rect 23100 15474 23156 15484
rect 22092 15314 22708 15316
rect 22092 15262 22094 15314
rect 22146 15262 22708 15314
rect 22092 15260 22708 15262
rect 22764 15316 22820 15326
rect 22092 15250 22148 15260
rect 22764 15222 22820 15260
rect 23100 15316 23156 15326
rect 23100 15222 23156 15260
rect 23212 15316 23268 15820
rect 23548 15540 23604 15934
rect 23548 15474 23604 15484
rect 24108 15540 24164 15550
rect 23324 15316 23380 15326
rect 23212 15260 23324 15316
rect 21980 12898 22036 12908
rect 22092 12964 22148 12974
rect 23212 12964 23268 15260
rect 23324 15222 23380 15260
rect 23884 15314 23940 15326
rect 23884 15262 23886 15314
rect 23938 15262 23940 15314
rect 23436 15204 23492 15214
rect 23436 14756 23492 15148
rect 23548 14756 23604 14766
rect 23436 14754 23604 14756
rect 23436 14702 23550 14754
rect 23602 14702 23604 14754
rect 23436 14700 23604 14702
rect 23548 14690 23604 14700
rect 23884 14754 23940 15262
rect 23884 14702 23886 14754
rect 23938 14702 23940 14754
rect 23884 14690 23940 14702
rect 23996 15204 24052 15214
rect 23884 14532 23940 14542
rect 23996 14532 24052 15148
rect 23884 14530 24052 14532
rect 23884 14478 23886 14530
rect 23938 14478 24052 14530
rect 23884 14476 24052 14478
rect 23884 14466 23940 14476
rect 23996 13858 24052 14476
rect 23996 13806 23998 13858
rect 24050 13806 24052 13858
rect 23996 13794 24052 13806
rect 24108 13858 24164 15484
rect 24220 15316 24276 15326
rect 24220 15222 24276 15260
rect 24332 15204 24388 16044
rect 24556 15988 24612 15998
rect 24556 15894 24612 15932
rect 24668 15986 24724 16156
rect 25004 16098 25060 16110
rect 25004 16046 25006 16098
rect 25058 16046 25060 16098
rect 24668 15934 24670 15986
rect 24722 15934 24724 15986
rect 24668 15922 24724 15934
rect 24892 15988 24948 15998
rect 24892 15894 24948 15932
rect 25004 15652 25060 16046
rect 25452 15988 25508 15998
rect 25452 15894 25508 15932
rect 25676 15988 25732 15998
rect 25676 15894 25732 15932
rect 24556 15596 25060 15652
rect 25340 15874 25396 15886
rect 25340 15822 25342 15874
rect 25394 15822 25396 15874
rect 24444 15540 24500 15550
rect 24444 15446 24500 15484
rect 24556 15538 24612 15596
rect 24556 15486 24558 15538
rect 24610 15486 24612 15538
rect 24556 15474 24612 15486
rect 25340 15428 25396 15822
rect 25340 15362 25396 15372
rect 24444 15204 24500 15214
rect 24332 15148 24444 15204
rect 25788 15148 25844 16156
rect 26124 15988 26180 16380
rect 26348 15988 26404 15998
rect 26124 15986 26404 15988
rect 26124 15934 26350 15986
rect 26402 15934 26404 15986
rect 26124 15932 26404 15934
rect 26012 15874 26068 15886
rect 26012 15822 26014 15874
rect 26066 15822 26068 15874
rect 26012 15540 26068 15822
rect 26012 15474 26068 15484
rect 24444 15138 24500 15148
rect 24108 13806 24110 13858
rect 24162 13806 24164 13858
rect 24108 13794 24164 13806
rect 24780 15092 24836 15102
rect 22092 12962 23268 12964
rect 22092 12910 22094 12962
rect 22146 12910 23268 12962
rect 22092 12908 23268 12910
rect 22092 12898 22148 12908
rect 23212 12850 23268 12908
rect 23212 12798 23214 12850
rect 23266 12798 23268 12850
rect 23212 12786 23268 12798
rect 23324 13748 23380 13758
rect 21308 12238 21310 12290
rect 21362 12238 21364 12290
rect 21308 12226 21364 12238
rect 21420 12572 21924 12628
rect 21980 12738 22036 12750
rect 21980 12686 21982 12738
rect 22034 12686 22036 12738
rect 21308 11508 21364 11518
rect 21196 11506 21364 11508
rect 21196 11454 21310 11506
rect 21362 11454 21364 11506
rect 21196 11452 21364 11454
rect 20860 10892 21140 10948
rect 17724 10770 17780 10780
rect 18396 10722 18452 10734
rect 18396 10670 18398 10722
rect 18450 10670 18452 10722
rect 18284 10612 18340 10622
rect 18284 10518 18340 10556
rect 17612 10444 18004 10500
rect 17500 10220 17892 10276
rect 17164 10050 17444 10052
rect 17164 9998 17166 10050
rect 17218 9998 17444 10050
rect 17164 9996 17444 9998
rect 17836 10052 17892 10220
rect 17164 9986 17220 9996
rect 17836 9958 17892 9996
rect 16940 9826 16996 9838
rect 16940 9774 16942 9826
rect 16994 9774 16996 9826
rect 16716 9426 16772 9436
rect 16828 9602 16884 9614
rect 16828 9550 16830 9602
rect 16882 9550 16884 9602
rect 16828 9268 16884 9550
rect 16940 9380 16996 9774
rect 17388 9828 17444 9838
rect 17388 9734 17444 9772
rect 17612 9826 17668 9838
rect 17612 9774 17614 9826
rect 17666 9774 17668 9826
rect 16940 9324 17444 9380
rect 16828 9212 16996 9268
rect 16492 9158 16494 9210
rect 16546 9158 16548 9210
rect 16492 9146 16548 9158
rect 16716 9044 16772 9054
rect 16268 8754 16324 8764
rect 16380 8988 16716 9044
rect 15428 5122 16156 5124
rect 15428 5070 15822 5122
rect 15874 5070 16156 5122
rect 15428 5068 16156 5070
rect 15372 5030 15428 5068
rect 15820 5058 15876 5068
rect 16156 5030 16212 5068
rect 16380 5572 16436 8988
rect 16716 8950 16772 8988
rect 16940 7364 16996 9212
rect 17388 9266 17444 9324
rect 17388 9214 17390 9266
rect 17442 9214 17444 9266
rect 17388 9202 17444 9214
rect 17612 9268 17668 9774
rect 17948 9828 18004 10444
rect 17948 9762 18004 9772
rect 18060 10386 18116 10398
rect 18060 10334 18062 10386
rect 18114 10334 18116 10386
rect 17948 9604 18004 9614
rect 17948 9510 18004 9548
rect 18060 9604 18116 10334
rect 18172 9604 18228 9614
rect 18060 9602 18228 9604
rect 18060 9550 18174 9602
rect 18226 9550 18228 9602
rect 18060 9548 18228 9550
rect 17612 9202 17668 9212
rect 17948 9156 18004 9166
rect 18060 9156 18116 9548
rect 18172 9538 18228 9548
rect 18172 9268 18228 9278
rect 18396 9268 18452 10670
rect 20860 10722 20916 10734
rect 20860 10670 20862 10722
rect 20914 10670 20916 10722
rect 20300 10612 20356 10622
rect 20300 10518 20356 10556
rect 19292 10052 19348 10062
rect 19068 9828 19124 9838
rect 19068 9734 19124 9772
rect 19292 9826 19348 9996
rect 19292 9774 19294 9826
rect 19346 9774 19348 9826
rect 19292 9762 19348 9774
rect 19628 10052 19684 10062
rect 19628 9826 19684 9996
rect 19852 10052 19908 10062
rect 20412 10052 20468 10062
rect 19852 10050 20244 10052
rect 19852 9998 19854 10050
rect 19906 9998 20244 10050
rect 19852 9996 20244 9998
rect 19852 9986 19908 9996
rect 19628 9774 19630 9826
rect 19682 9774 19684 9826
rect 19628 9762 19684 9774
rect 19852 9828 19908 9838
rect 19852 9734 19908 9772
rect 19628 9602 19684 9614
rect 19628 9550 19630 9602
rect 19682 9550 19684 9602
rect 18172 9266 18452 9268
rect 18172 9214 18174 9266
rect 18226 9214 18452 9266
rect 18172 9212 18452 9214
rect 18620 9492 18676 9502
rect 18172 9202 18228 9212
rect 17948 9154 18116 9156
rect 17948 9102 17950 9154
rect 18002 9102 18116 9154
rect 17948 9100 18116 9102
rect 17948 9090 18004 9100
rect 17836 9044 17892 9054
rect 17836 8950 17892 8988
rect 17500 8930 17556 8942
rect 17500 8878 17502 8930
rect 17554 8878 17556 8930
rect 17500 8820 17556 8878
rect 18060 8820 18116 9100
rect 17500 8764 18116 8820
rect 14252 4398 14254 4450
rect 14306 4398 14308 4450
rect 14252 4386 14308 4398
rect 13580 4286 13582 4338
rect 13634 4286 13636 4338
rect 13580 4274 13636 4286
rect 16380 4226 16436 5516
rect 16492 7308 16996 7364
rect 16492 5234 16548 7308
rect 18060 6578 18116 8764
rect 18060 6526 18062 6578
rect 18114 6526 18116 6578
rect 18060 6514 18116 6526
rect 18396 6578 18452 6590
rect 18396 6526 18398 6578
rect 18450 6526 18452 6578
rect 18396 5908 18452 6526
rect 18620 6130 18676 9436
rect 18620 6078 18622 6130
rect 18674 6078 18676 6130
rect 18620 6066 18676 6078
rect 19068 6018 19124 6030
rect 19068 5966 19070 6018
rect 19122 5966 19124 6018
rect 18508 5908 18564 5918
rect 18396 5906 18676 5908
rect 18396 5854 18510 5906
rect 18562 5854 18676 5906
rect 18396 5852 18676 5854
rect 18508 5842 18564 5852
rect 16492 5182 16494 5234
rect 16546 5182 16548 5234
rect 16492 5170 16548 5182
rect 18620 5234 18676 5852
rect 18956 5572 19012 5582
rect 19068 5572 19124 5966
rect 19012 5516 19124 5572
rect 18956 5506 19012 5516
rect 18620 5182 18622 5234
rect 18674 5182 18676 5234
rect 18620 5170 18676 5182
rect 16828 5124 16884 5134
rect 16828 4564 16884 5068
rect 16828 4470 16884 4508
rect 18732 4564 18788 4574
rect 18732 4470 18788 4508
rect 19180 4564 19236 4574
rect 19628 4564 19684 9550
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20076 9268 20132 9278
rect 20076 9154 20132 9212
rect 20188 9266 20244 9996
rect 20412 9958 20468 9996
rect 20860 10052 20916 10670
rect 20860 9986 20916 9996
rect 20524 9716 20580 9726
rect 20188 9214 20190 9266
rect 20242 9214 20244 9266
rect 20188 9202 20244 9214
rect 20412 9714 20580 9716
rect 20412 9662 20526 9714
rect 20578 9662 20580 9714
rect 20412 9660 20580 9662
rect 20076 9102 20078 9154
rect 20130 9102 20132 9154
rect 20076 9090 20132 9102
rect 20412 9042 20468 9660
rect 20524 9650 20580 9660
rect 21084 9268 21140 10892
rect 21084 9174 21140 9212
rect 20412 8990 20414 9042
rect 20466 8990 20468 9042
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20412 5012 20468 8990
rect 20636 9044 20692 9054
rect 21196 9044 21252 11452
rect 21308 11442 21364 11452
rect 21420 11282 21476 12572
rect 21980 12516 22036 12686
rect 21532 12460 22036 12516
rect 22092 12740 22148 12750
rect 21532 12290 21588 12460
rect 21756 12348 22036 12404
rect 21532 12238 21534 12290
rect 21586 12238 21588 12290
rect 21532 12226 21588 12238
rect 21644 12290 21700 12302
rect 21644 12238 21646 12290
rect 21698 12238 21700 12290
rect 21644 12180 21700 12238
rect 21756 12290 21812 12348
rect 21756 12238 21758 12290
rect 21810 12238 21812 12290
rect 21756 12226 21812 12238
rect 21644 12068 21700 12124
rect 21420 11230 21422 11282
rect 21474 11230 21476 11282
rect 21420 11218 21476 11230
rect 21532 12012 21700 12068
rect 21868 12178 21924 12190
rect 21868 12126 21870 12178
rect 21922 12126 21924 12178
rect 20636 9042 21252 9044
rect 20636 8990 20638 9042
rect 20690 8990 21252 9042
rect 20636 8988 21252 8990
rect 20636 8978 20692 8988
rect 21084 6020 21140 6030
rect 21532 6020 21588 12012
rect 21868 11956 21924 12126
rect 21644 11900 21868 11956
rect 21644 11282 21700 11900
rect 21868 11890 21924 11900
rect 21980 11508 22036 12348
rect 21644 11230 21646 11282
rect 21698 11230 21700 11282
rect 21644 10498 21700 11230
rect 21644 10446 21646 10498
rect 21698 10446 21700 10498
rect 21644 10434 21700 10446
rect 21756 11452 22036 11508
rect 22092 11508 22148 12684
rect 22876 12738 22932 12750
rect 22876 12686 22878 12738
rect 22930 12686 22932 12738
rect 22876 12628 22932 12686
rect 23324 12628 23380 13692
rect 24220 13748 24276 13758
rect 24220 13654 24276 13692
rect 24668 13524 24724 13534
rect 22764 12572 23380 12628
rect 24220 13522 24724 13524
rect 24220 13470 24670 13522
rect 24722 13470 24724 13522
rect 24220 13468 24724 13470
rect 22764 12402 22820 12572
rect 22764 12350 22766 12402
rect 22818 12350 22820 12402
rect 22764 12338 22820 12350
rect 22204 12180 22260 12190
rect 22204 12086 22260 12124
rect 22428 11956 22484 11966
rect 22428 11862 22484 11900
rect 22204 11508 22260 11518
rect 22092 11506 22260 11508
rect 22092 11454 22206 11506
rect 22258 11454 22260 11506
rect 22092 11452 22260 11454
rect 21644 6692 21700 6702
rect 21756 6692 21812 11452
rect 22204 11442 22260 11452
rect 24220 10724 24276 13468
rect 24668 13458 24724 13468
rect 24780 12516 24836 15036
rect 24556 12460 24836 12516
rect 25676 15092 25844 15148
rect 25900 15204 25956 15214
rect 25956 15148 26292 15204
rect 25900 15110 25956 15148
rect 24556 11506 24612 12460
rect 25564 11620 25620 11630
rect 24556 11454 24558 11506
rect 24610 11454 24612 11506
rect 24556 11396 24612 11454
rect 24556 11330 24612 11340
rect 25228 11618 25620 11620
rect 25228 11566 25566 11618
rect 25618 11566 25620 11618
rect 25228 11564 25620 11566
rect 25116 11284 25172 11294
rect 25116 11190 25172 11228
rect 24780 11170 24836 11182
rect 24780 11118 24782 11170
rect 24834 11118 24836 11170
rect 24444 10836 24500 10846
rect 24444 10742 24500 10780
rect 24668 10836 24724 10846
rect 24668 10742 24724 10780
rect 24220 10630 24276 10668
rect 24668 10498 24724 10510
rect 24668 10446 24670 10498
rect 24722 10446 24724 10498
rect 24668 9604 24724 10446
rect 24668 9538 24724 9548
rect 24780 9826 24836 11118
rect 25004 11170 25060 11182
rect 25004 11118 25006 11170
rect 25058 11118 25060 11170
rect 25004 10948 25060 11118
rect 25004 10882 25060 10892
rect 25228 10388 25284 11564
rect 25564 11554 25620 11564
rect 25452 11396 25508 11406
rect 25452 11302 25508 11340
rect 25564 11170 25620 11182
rect 25564 11118 25566 11170
rect 25618 11118 25620 11170
rect 25564 10836 25620 11118
rect 25676 10836 25732 15092
rect 26236 13746 26292 15148
rect 26348 13858 26404 15932
rect 27244 13970 27300 19068
rect 28588 15876 28644 22204
rect 29932 20018 29988 20030
rect 29932 19966 29934 20018
rect 29986 19966 29988 20018
rect 28700 19908 28756 19918
rect 28700 19814 28756 19852
rect 29932 19908 29988 19966
rect 29260 19796 29316 19806
rect 29260 19702 29316 19740
rect 29260 19348 29316 19358
rect 29260 16212 29316 19292
rect 29932 19236 29988 19852
rect 30044 20020 30100 20030
rect 30044 19906 30100 19964
rect 30044 19854 30046 19906
rect 30098 19854 30100 19906
rect 30044 19842 30100 19854
rect 30044 19348 30100 19358
rect 30156 19348 30212 23884
rect 31164 23378 31220 24220
rect 31164 23326 31166 23378
rect 31218 23326 31220 23378
rect 31164 23314 31220 23326
rect 31276 24052 31332 24062
rect 31276 23266 31332 23996
rect 32060 24052 32116 24062
rect 32060 23958 32116 23996
rect 32172 23380 32228 26852
rect 32396 26852 32452 26862
rect 32844 26852 33124 26908
rect 32396 24050 32452 26796
rect 33068 26514 33124 26852
rect 33068 26462 33070 26514
rect 33122 26462 33124 26514
rect 33068 26450 33124 26462
rect 33292 26852 33348 26862
rect 33292 26514 33348 26796
rect 33292 26462 33294 26514
rect 33346 26462 33348 26514
rect 33292 26450 33348 26462
rect 33516 26402 33572 26414
rect 33516 26350 33518 26402
rect 33570 26350 33572 26402
rect 32508 26292 32564 26302
rect 32508 26178 32564 26236
rect 33516 26292 33572 26350
rect 33516 26226 33572 26236
rect 32508 26126 32510 26178
rect 32562 26126 32564 26178
rect 32508 25172 32564 26126
rect 33180 26180 33236 26190
rect 33180 26086 33236 26124
rect 34748 25620 34804 32060
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35308 30212 35364 30222
rect 35980 30212 36036 32508
rect 36428 31554 36484 31566
rect 36428 31502 36430 31554
rect 36482 31502 36484 31554
rect 36428 31444 36484 31502
rect 36428 31378 36484 31388
rect 35308 30210 36036 30212
rect 35308 30158 35310 30210
rect 35362 30158 36036 30210
rect 35308 30156 36036 30158
rect 35308 30146 35364 30156
rect 34972 30100 35028 30110
rect 34972 30006 35028 30044
rect 35980 30098 36036 30156
rect 35980 30046 35982 30098
rect 36034 30046 36036 30098
rect 35980 30034 36036 30046
rect 36652 31106 36708 34972
rect 37660 35028 37716 36540
rect 37660 34962 37716 34972
rect 37660 34020 37716 34030
rect 37100 34018 37716 34020
rect 37100 33966 37662 34018
rect 37714 33966 37716 34018
rect 37100 33964 37716 33966
rect 37100 33458 37156 33964
rect 37660 33954 37716 33964
rect 37100 33406 37102 33458
rect 37154 33406 37156 33458
rect 37100 33394 37156 33406
rect 37324 33404 37828 33460
rect 37324 33346 37380 33404
rect 37324 33294 37326 33346
rect 37378 33294 37380 33346
rect 37324 33282 37380 33294
rect 37772 33346 37828 33404
rect 37772 33294 37774 33346
rect 37826 33294 37828 33346
rect 37772 33282 37828 33294
rect 36988 33234 37044 33246
rect 36988 33182 36990 33234
rect 37042 33182 37044 33234
rect 36876 32788 36932 32798
rect 36988 32788 37044 33182
rect 37212 33236 37268 33246
rect 37100 32788 37156 32798
rect 36988 32786 37156 32788
rect 36988 32734 37102 32786
rect 37154 32734 37156 32786
rect 36988 32732 37156 32734
rect 36876 32694 36932 32732
rect 37100 32722 37156 32732
rect 37212 32786 37268 33180
rect 37548 33234 37604 33246
rect 37548 33182 37550 33234
rect 37602 33182 37604 33234
rect 37212 32734 37214 32786
rect 37266 32734 37268 32786
rect 37212 32722 37268 32734
rect 37324 32900 37380 32910
rect 37548 32900 37604 33182
rect 37380 32844 37604 32900
rect 36764 32564 36820 32574
rect 36764 32470 36820 32508
rect 36988 31554 37044 31566
rect 36988 31502 36990 31554
rect 37042 31502 37044 31554
rect 36988 31444 37044 31502
rect 37324 31556 37380 32844
rect 37436 32674 37492 32686
rect 37436 32622 37438 32674
rect 37490 32622 37492 32674
rect 37436 31780 37492 32622
rect 37548 32564 37604 32574
rect 37548 32004 37604 32508
rect 37548 31938 37604 31948
rect 37436 31714 37492 31724
rect 37324 31554 37492 31556
rect 37324 31502 37326 31554
rect 37378 31502 37492 31554
rect 37324 31500 37492 31502
rect 37324 31490 37380 31500
rect 36988 31378 37044 31388
rect 36652 31054 36654 31106
rect 36706 31054 36708 31106
rect 35196 29986 35252 29998
rect 35196 29934 35198 29986
rect 35250 29934 35252 29986
rect 34860 29316 34916 29326
rect 35196 29316 35252 29934
rect 34860 29314 35252 29316
rect 34860 29262 34862 29314
rect 34914 29262 35252 29314
rect 34860 29260 35252 29262
rect 35644 29986 35700 29998
rect 35644 29934 35646 29986
rect 35698 29934 35700 29986
rect 35644 29876 35700 29934
rect 34860 29204 34916 29260
rect 35644 29204 35700 29820
rect 34860 29138 34916 29148
rect 35084 29148 35700 29204
rect 36316 29988 36372 29998
rect 34972 28420 35028 28430
rect 34972 28326 35028 28364
rect 34636 25564 34748 25620
rect 32620 25172 32676 25182
rect 32508 25116 32620 25172
rect 32396 23998 32398 24050
rect 32450 23998 32452 24050
rect 32396 23986 32452 23998
rect 32396 23380 32452 23390
rect 32172 23378 32452 23380
rect 32172 23326 32398 23378
rect 32450 23326 32452 23378
rect 32172 23324 32452 23326
rect 32396 23314 32452 23324
rect 31276 23214 31278 23266
rect 31330 23214 31332 23266
rect 31276 23202 31332 23214
rect 30044 19346 30212 19348
rect 30044 19294 30046 19346
rect 30098 19294 30212 19346
rect 30044 19292 30212 19294
rect 30044 19282 30100 19292
rect 29932 19170 29988 19180
rect 30156 19012 30212 19292
rect 30380 20020 30436 20030
rect 30380 19234 30436 19964
rect 31388 20020 31444 20030
rect 31388 19926 31444 19964
rect 31948 19908 32004 19918
rect 31948 19906 32228 19908
rect 31948 19854 31950 19906
rect 32002 19854 32228 19906
rect 31948 19852 32228 19854
rect 31948 19842 32004 19852
rect 31724 19794 31780 19806
rect 31724 19742 31726 19794
rect 31778 19742 31780 19794
rect 30380 19182 30382 19234
rect 30434 19182 30436 19234
rect 30380 19170 30436 19182
rect 30716 19236 30772 19246
rect 31500 19236 31556 19246
rect 30716 19234 31556 19236
rect 30716 19182 30718 19234
rect 30770 19182 31502 19234
rect 31554 19182 31556 19234
rect 30716 19180 31556 19182
rect 30716 19170 30772 19180
rect 31500 19170 31556 19180
rect 30156 18946 30212 18956
rect 30604 19012 30660 19022
rect 31164 19012 31220 19022
rect 30604 19010 31108 19012
rect 30604 18958 30606 19010
rect 30658 18958 31108 19010
rect 30604 18956 31108 18958
rect 30604 18946 30660 18956
rect 29484 18900 29540 18910
rect 29484 18338 29540 18844
rect 31052 18676 31108 18956
rect 31164 18918 31220 18956
rect 31388 19010 31444 19022
rect 31388 18958 31390 19010
rect 31442 18958 31444 19010
rect 31388 18900 31444 18958
rect 31612 19012 31668 19022
rect 31724 19012 31780 19742
rect 32060 19236 32116 19246
rect 32060 19142 32116 19180
rect 32172 19124 32228 19852
rect 32172 19030 32228 19068
rect 31612 19010 31780 19012
rect 31612 18958 31614 19010
rect 31666 18958 31780 19010
rect 31612 18956 31780 18958
rect 31612 18946 31668 18956
rect 31388 18834 31444 18844
rect 31052 18620 31668 18676
rect 31612 18562 31668 18620
rect 31612 18510 31614 18562
rect 31666 18510 31668 18562
rect 31612 18498 31668 18510
rect 29484 18286 29486 18338
rect 29538 18286 29540 18338
rect 29484 18274 29540 18286
rect 31724 18228 31780 18956
rect 32396 18450 32452 18462
rect 32396 18398 32398 18450
rect 32450 18398 32452 18450
rect 32396 18340 32452 18398
rect 32396 18274 32452 18284
rect 31612 18172 31780 18228
rect 28700 15876 28756 15886
rect 28588 15820 28700 15876
rect 28700 15782 28756 15820
rect 29260 15540 29316 16156
rect 29372 17108 29428 17118
rect 29372 16098 29428 17052
rect 29372 16046 29374 16098
rect 29426 16046 29428 16098
rect 29372 15876 29428 16046
rect 29372 15810 29428 15820
rect 28812 15538 29652 15540
rect 28812 15486 29262 15538
rect 29314 15486 29652 15538
rect 28812 15484 29652 15486
rect 28028 15428 28084 15438
rect 28028 15334 28084 15372
rect 28812 15314 28868 15484
rect 29260 15474 29316 15484
rect 28812 15262 28814 15314
rect 28866 15262 28868 15314
rect 28812 15250 28868 15262
rect 29596 15314 29652 15484
rect 29596 15262 29598 15314
rect 29650 15262 29652 15314
rect 29596 15250 29652 15262
rect 30380 15204 30436 15214
rect 30380 15202 31556 15204
rect 30380 15150 30382 15202
rect 30434 15150 31556 15202
rect 30380 15148 31556 15150
rect 30380 15138 30436 15148
rect 31500 14642 31556 15148
rect 31500 14590 31502 14642
rect 31554 14590 31556 14642
rect 31500 14578 31556 14590
rect 27244 13918 27246 13970
rect 27298 13918 27300 13970
rect 27244 13906 27300 13918
rect 31388 14418 31444 14430
rect 31612 14420 31668 18172
rect 31948 16212 32004 16222
rect 31948 16118 32004 16156
rect 32508 15204 32564 15214
rect 32508 15110 32564 15148
rect 32620 14980 32676 25116
rect 34524 24612 34580 24622
rect 34524 24050 34580 24556
rect 34524 23998 34526 24050
rect 34578 23998 34580 24050
rect 34524 23986 34580 23998
rect 34636 23378 34692 25564
rect 34748 25554 34804 25564
rect 34636 23326 34638 23378
rect 34690 23326 34692 23378
rect 34636 23314 34692 23326
rect 34972 24500 35028 24510
rect 35084 24500 35140 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35980 28644 36036 28654
rect 35980 28550 36036 28588
rect 36316 28530 36372 29932
rect 36428 29986 36484 29998
rect 36428 29934 36430 29986
rect 36482 29934 36484 29986
rect 36428 29876 36484 29934
rect 36428 29810 36484 29820
rect 36652 29652 36708 31054
rect 37436 30210 37492 31500
rect 37436 30158 37438 30210
rect 37490 30158 37492 30210
rect 36988 30100 37044 30110
rect 36988 30006 37044 30044
rect 37324 30100 37380 30110
rect 37324 30006 37380 30044
rect 36652 29586 36708 29596
rect 37100 29986 37156 29998
rect 37100 29934 37102 29986
rect 37154 29934 37156 29986
rect 36988 29540 37044 29550
rect 37100 29540 37156 29934
rect 36988 29538 37156 29540
rect 36988 29486 36990 29538
rect 37042 29486 37156 29538
rect 36988 29484 37156 29486
rect 36988 29474 37044 29484
rect 36316 28478 36318 28530
rect 36370 28478 36372 28530
rect 36316 28466 36372 28478
rect 36988 28420 37044 28430
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 36652 26964 36708 26974
rect 36652 26402 36708 26908
rect 36988 26514 37044 28364
rect 36988 26462 36990 26514
rect 37042 26462 37044 26514
rect 36988 26450 37044 26462
rect 37324 26852 37380 26862
rect 36652 26350 36654 26402
rect 36706 26350 36708 26402
rect 36652 26338 36708 26350
rect 36764 26404 36820 26414
rect 36764 26310 36820 26348
rect 36204 26290 36260 26302
rect 36204 26238 36206 26290
rect 36258 26238 36260 26290
rect 35868 26180 35924 26190
rect 36204 26180 36260 26238
rect 36652 26180 36708 26190
rect 35868 26178 36260 26180
rect 35868 26126 35870 26178
rect 35922 26126 36260 26178
rect 35868 26124 36260 26126
rect 36428 26178 36708 26180
rect 36428 26126 36654 26178
rect 36706 26126 36708 26178
rect 36428 26124 36708 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35868 24948 35924 26124
rect 35980 25620 36036 25630
rect 35980 25526 36036 25564
rect 36428 25618 36484 26124
rect 36652 26114 36708 26124
rect 36428 25566 36430 25618
rect 36482 25566 36484 25618
rect 36428 25554 36484 25566
rect 36988 25620 37044 25630
rect 36988 25506 37044 25564
rect 36988 25454 36990 25506
rect 37042 25454 37044 25506
rect 36988 25442 37044 25454
rect 37324 25394 37380 26796
rect 37324 25342 37326 25394
rect 37378 25342 37380 25394
rect 37324 25330 37380 25342
rect 36316 25284 36372 25294
rect 35868 24882 35924 24892
rect 36204 25282 36372 25284
rect 36204 25230 36318 25282
rect 36370 25230 36372 25282
rect 36204 25228 36372 25230
rect 36204 24834 36260 25228
rect 36316 25218 36372 25228
rect 36204 24782 36206 24834
rect 36258 24782 36260 24834
rect 36204 24770 36260 24782
rect 35028 24444 35140 24500
rect 35532 24724 35588 24734
rect 34860 23154 34916 23166
rect 34860 23102 34862 23154
rect 34914 23102 34916 23154
rect 34860 23044 34916 23102
rect 34636 22988 34860 23044
rect 34636 21026 34692 22988
rect 34860 22978 34916 22988
rect 34972 22820 35028 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35308 23940 35364 23950
rect 35532 23940 35588 24668
rect 35868 23940 35924 23950
rect 35308 23938 35924 23940
rect 35308 23886 35310 23938
rect 35362 23886 35870 23938
rect 35922 23886 35924 23938
rect 35308 23884 35924 23886
rect 35308 23874 35364 23884
rect 35868 23874 35924 23884
rect 35420 23044 35476 23054
rect 35420 22950 35476 22988
rect 34636 20974 34638 21026
rect 34690 20974 34692 21026
rect 34636 20962 34692 20974
rect 34860 22764 35028 22820
rect 35196 22764 35460 22774
rect 34860 20244 34916 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 36092 21586 36148 21598
rect 36092 21534 36094 21586
rect 36146 21534 36148 21586
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34972 20692 35028 20702
rect 34972 20690 35140 20692
rect 34972 20638 34974 20690
rect 35026 20638 35140 20690
rect 34972 20636 35140 20638
rect 34972 20626 35028 20636
rect 34972 20244 35028 20254
rect 34860 20242 35028 20244
rect 34860 20190 34974 20242
rect 35026 20190 35028 20242
rect 34860 20188 35028 20190
rect 34972 20178 35028 20188
rect 35084 20020 35140 20636
rect 35196 20690 35252 20702
rect 35196 20638 35198 20690
rect 35250 20638 35252 20690
rect 35196 20132 35252 20638
rect 35196 20066 35252 20076
rect 35420 20690 35476 20702
rect 35420 20638 35422 20690
rect 35474 20638 35476 20690
rect 35420 20130 35476 20638
rect 36092 20356 36148 21534
rect 36876 21476 36932 21486
rect 36876 21474 37380 21476
rect 36876 21422 36878 21474
rect 36930 21422 37380 21474
rect 36876 21420 37380 21422
rect 36876 21410 36932 21420
rect 37324 20914 37380 21420
rect 37324 20862 37326 20914
rect 37378 20862 37380 20914
rect 37324 20850 37380 20862
rect 37212 20692 37268 20702
rect 37436 20692 37492 30158
rect 37772 29652 37828 29662
rect 37772 29426 37828 29596
rect 37772 29374 37774 29426
rect 37826 29374 37828 29426
rect 37772 29362 37828 29374
rect 37884 27074 37940 38222
rect 38332 38162 38388 38892
rect 40124 38948 40180 38958
rect 40124 38854 40180 38892
rect 40012 38834 40068 38846
rect 40012 38782 40014 38834
rect 40066 38782 40068 38834
rect 38332 38110 38334 38162
rect 38386 38110 38388 38162
rect 38332 38098 38388 38110
rect 39676 38724 39732 38734
rect 40012 38724 40068 38782
rect 41132 38834 41188 39004
rect 41132 38782 41134 38834
rect 41186 38782 41188 38834
rect 41132 38770 41188 38782
rect 39676 38722 40068 38724
rect 39676 38670 39678 38722
rect 39730 38670 40068 38722
rect 39676 38668 40068 38670
rect 38108 38050 38164 38062
rect 38108 37998 38110 38050
rect 38162 37998 38164 38050
rect 38108 37044 38164 37998
rect 39676 37828 39732 38668
rect 41804 38276 41860 39566
rect 42140 39506 42196 39518
rect 42140 39454 42142 39506
rect 42194 39454 42196 39506
rect 40796 38220 41860 38276
rect 41916 38722 41972 38734
rect 41916 38670 41918 38722
rect 41970 38670 41972 38722
rect 41916 38276 41972 38670
rect 42140 38276 42196 39454
rect 41916 38220 42084 38276
rect 40460 38052 40516 38062
rect 40460 37938 40516 37996
rect 40796 38050 40852 38220
rect 41356 38108 41860 38164
rect 40796 37998 40798 38050
rect 40850 37998 40852 38050
rect 40796 37986 40852 37998
rect 41020 38052 41076 38062
rect 41020 37958 41076 37996
rect 41356 38050 41412 38108
rect 41356 37998 41358 38050
rect 41410 37998 41412 38050
rect 41356 37986 41412 37998
rect 41804 38050 41860 38108
rect 42028 38162 42084 38220
rect 42140 38210 42196 38220
rect 44044 38722 44100 38734
rect 44044 38670 44046 38722
rect 44098 38670 44100 38722
rect 42028 38110 42030 38162
rect 42082 38110 42084 38162
rect 42028 38098 42084 38110
rect 41804 37998 41806 38050
rect 41858 37998 41860 38050
rect 41804 37986 41860 37998
rect 41916 38052 41972 38062
rect 40460 37886 40462 37938
rect 40514 37886 40516 37938
rect 39676 37762 39732 37772
rect 39788 37828 39844 37838
rect 40236 37828 40292 37838
rect 40460 37828 40516 37886
rect 41244 37940 41300 37950
rect 39788 37826 40516 37828
rect 39788 37774 39790 37826
rect 39842 37774 40238 37826
rect 40290 37774 40516 37826
rect 39788 37772 40516 37774
rect 40572 37828 40628 37838
rect 38108 36978 38164 36988
rect 38220 37156 38276 37166
rect 38108 33234 38164 33246
rect 38108 33182 38110 33234
rect 38162 33182 38164 33234
rect 37996 33124 38052 33134
rect 37996 33030 38052 33068
rect 38108 29988 38164 33182
rect 38220 31780 38276 37100
rect 38332 35028 38388 35038
rect 38332 34130 38388 34972
rect 38892 35028 38948 35038
rect 38892 34354 38948 34972
rect 38892 34302 38894 34354
rect 38946 34302 38948 34354
rect 38892 34290 38948 34302
rect 38332 34078 38334 34130
rect 38386 34078 38388 34130
rect 38332 34066 38388 34078
rect 39788 33012 39844 37772
rect 40236 37762 40292 37772
rect 40572 37734 40628 37772
rect 41132 37826 41188 37838
rect 41132 37774 41134 37826
rect 41186 37774 41188 37826
rect 41132 37268 41188 37774
rect 41132 37202 41188 37212
rect 41244 35924 41300 37884
rect 41580 37938 41636 37950
rect 41580 37886 41582 37938
rect 41634 37886 41636 37938
rect 41580 37828 41636 37886
rect 41916 37828 41972 37996
rect 42140 37940 42196 37950
rect 42364 37940 42420 37950
rect 42140 37938 42420 37940
rect 42140 37886 42142 37938
rect 42194 37886 42366 37938
rect 42418 37886 42420 37938
rect 42140 37884 42420 37886
rect 42140 37874 42196 37884
rect 42364 37874 42420 37884
rect 42700 37940 42756 37950
rect 42700 37846 42756 37884
rect 43148 37940 43204 37950
rect 43148 37846 43204 37884
rect 44044 37940 44100 38670
rect 44044 37874 44100 37884
rect 42588 37828 42644 37838
rect 41580 37772 42084 37828
rect 41692 35980 41972 36036
rect 41356 35924 41412 35934
rect 41692 35924 41748 35980
rect 41244 35922 41748 35924
rect 41244 35870 41358 35922
rect 41410 35870 41748 35922
rect 41244 35868 41748 35870
rect 41356 35858 41412 35868
rect 41804 35810 41860 35822
rect 41804 35758 41806 35810
rect 41858 35758 41860 35810
rect 41580 35698 41636 35710
rect 41580 35646 41582 35698
rect 41634 35646 41636 35698
rect 40572 35028 40628 35038
rect 40572 34934 40628 34972
rect 41020 35028 41076 35038
rect 41020 34914 41076 34972
rect 41020 34862 41022 34914
rect 41074 34862 41076 34914
rect 41020 34850 41076 34862
rect 41580 34356 41636 35646
rect 41804 35028 41860 35758
rect 41916 35810 41972 35980
rect 41916 35758 41918 35810
rect 41970 35758 41972 35810
rect 41916 35746 41972 35758
rect 41804 34916 41860 34972
rect 41804 34860 41972 34916
rect 41692 34804 41748 34814
rect 41692 34802 41860 34804
rect 41692 34750 41694 34802
rect 41746 34750 41860 34802
rect 41692 34748 41860 34750
rect 41692 34738 41748 34748
rect 41580 34300 41748 34356
rect 39788 32946 39844 32956
rect 41468 33906 41524 33918
rect 41468 33854 41470 33906
rect 41522 33854 41524 33906
rect 40348 32340 40404 32350
rect 40012 31892 40068 31902
rect 40068 31836 40180 31892
rect 40012 31826 40068 31836
rect 38220 31714 38276 31724
rect 39004 31780 39060 31790
rect 38108 29922 38164 29932
rect 38220 29652 38276 29662
rect 38220 29558 38276 29596
rect 37884 27022 37886 27074
rect 37938 27022 37940 27074
rect 37884 27010 37940 27022
rect 37548 26964 37604 27002
rect 37548 26898 37604 26908
rect 37772 26852 37828 26862
rect 37772 26758 37828 26796
rect 38332 26404 38388 26414
rect 38332 24610 38388 26348
rect 39004 25506 39060 31724
rect 39676 31556 39732 31566
rect 40012 31556 40068 31566
rect 39676 31554 40068 31556
rect 39676 31502 39678 31554
rect 39730 31502 40014 31554
rect 40066 31502 40068 31554
rect 39676 31500 40068 31502
rect 39676 31444 39732 31500
rect 40012 31490 40068 31500
rect 39676 31378 39732 31388
rect 40124 31332 40180 31836
rect 40348 31666 40404 32284
rect 41468 31948 41524 33854
rect 41692 33346 41748 34300
rect 41804 33458 41860 34748
rect 41916 34018 41972 34860
rect 41916 33966 41918 34018
rect 41970 33966 41972 34018
rect 41916 33954 41972 33966
rect 42028 34020 42084 37772
rect 42588 37734 42644 37772
rect 42140 37268 42196 37278
rect 42196 37212 42308 37268
rect 42140 37202 42196 37212
rect 42252 34130 42308 37212
rect 43820 35028 43876 35038
rect 43820 34934 43876 34972
rect 42252 34078 42254 34130
rect 42306 34078 42308 34130
rect 42252 34066 42308 34078
rect 42028 33964 42196 34020
rect 41804 33406 41806 33458
rect 41858 33406 41860 33458
rect 41804 33394 41860 33406
rect 41692 33294 41694 33346
rect 41746 33294 41748 33346
rect 41692 33282 41748 33294
rect 42140 33348 42196 33964
rect 42252 33348 42308 33358
rect 42140 33346 42308 33348
rect 42140 33294 42254 33346
rect 42306 33294 42308 33346
rect 42140 33292 42308 33294
rect 42028 33236 42084 33246
rect 42028 33234 42196 33236
rect 42028 33182 42030 33234
rect 42082 33182 42196 33234
rect 42028 33180 42196 33182
rect 42028 33170 42084 33180
rect 42140 32786 42196 33180
rect 42140 32734 42142 32786
rect 42194 32734 42196 32786
rect 42140 32722 42196 32734
rect 41916 32674 41972 32686
rect 41916 32622 41918 32674
rect 41970 32622 41972 32674
rect 41804 32564 41860 32574
rect 40348 31614 40350 31666
rect 40402 31614 40404 31666
rect 40348 31602 40404 31614
rect 41356 31892 41524 31948
rect 41692 32562 41860 32564
rect 41692 32510 41806 32562
rect 41858 32510 41860 32562
rect 41692 32508 41860 32510
rect 41916 32564 41972 32622
rect 41916 32508 42084 32564
rect 40012 31276 40180 31332
rect 40012 31106 40068 31276
rect 40012 31054 40014 31106
rect 40066 31054 40068 31106
rect 40012 31042 40068 31054
rect 40124 31106 40180 31118
rect 40124 31054 40126 31106
rect 40178 31054 40180 31106
rect 39340 30324 39396 30334
rect 39116 30100 39172 30110
rect 39116 30006 39172 30044
rect 39340 30098 39396 30268
rect 40124 30324 40180 31054
rect 40348 30996 40404 31006
rect 40348 30902 40404 30940
rect 41132 30996 41188 31006
rect 41132 30902 41188 30940
rect 40124 30258 40180 30268
rect 40684 30210 40740 30222
rect 40684 30158 40686 30210
rect 40738 30158 40740 30210
rect 39340 30046 39342 30098
rect 39394 30046 39396 30098
rect 39340 30034 39396 30046
rect 39452 30098 39508 30110
rect 39452 30046 39454 30098
rect 39506 30046 39508 30098
rect 39452 29988 39508 30046
rect 39452 29922 39508 29932
rect 40348 29988 40404 29998
rect 40684 29988 40740 30158
rect 40348 29986 40740 29988
rect 40348 29934 40350 29986
rect 40402 29934 40740 29986
rect 40348 29932 40740 29934
rect 40348 29316 40404 29932
rect 41356 29428 41412 31892
rect 41468 31218 41524 31230
rect 41468 31166 41470 31218
rect 41522 31166 41524 31218
rect 41468 30322 41524 31166
rect 41468 30270 41470 30322
rect 41522 30270 41524 30322
rect 41468 30258 41524 30270
rect 41580 30994 41636 31006
rect 41580 30942 41582 30994
rect 41634 30942 41636 30994
rect 41468 29652 41524 29662
rect 41580 29652 41636 30942
rect 41692 29988 41748 32508
rect 41804 32498 41860 32508
rect 41804 32340 41860 32350
rect 41804 31106 41860 32284
rect 42028 32116 42084 32508
rect 42252 32340 42308 33292
rect 42252 32274 42308 32284
rect 41804 31054 41806 31106
rect 41858 31054 41860 31106
rect 41804 31042 41860 31054
rect 41916 32060 42084 32116
rect 41748 29932 41860 29988
rect 41692 29922 41748 29932
rect 41468 29650 41636 29652
rect 41468 29598 41470 29650
rect 41522 29598 41636 29650
rect 41468 29596 41636 29598
rect 41468 29586 41524 29596
rect 41692 29538 41748 29550
rect 41692 29486 41694 29538
rect 41746 29486 41748 29538
rect 41356 29372 41636 29428
rect 40348 26964 40404 29260
rect 41244 27972 41300 27982
rect 41020 27074 41076 27086
rect 41020 27022 41022 27074
rect 41074 27022 41076 27074
rect 40684 26964 40740 26974
rect 41020 26964 41076 27022
rect 40236 26962 41076 26964
rect 40236 26910 40686 26962
rect 40738 26910 41076 26962
rect 40236 26908 41076 26910
rect 39228 26404 39284 26414
rect 39228 25618 39284 26348
rect 39228 25566 39230 25618
rect 39282 25566 39284 25618
rect 39228 25554 39284 25566
rect 39004 25454 39006 25506
rect 39058 25454 39060 25506
rect 39004 25442 39060 25454
rect 39900 25394 39956 25406
rect 39900 25342 39902 25394
rect 39954 25342 39956 25394
rect 39900 25060 39956 25342
rect 39900 24994 39956 25004
rect 38780 24724 38836 24734
rect 38780 24630 38836 24668
rect 40236 24724 40292 26908
rect 40684 26898 40740 26908
rect 41244 26852 41300 27916
rect 41580 27858 41636 29372
rect 41692 28196 41748 29486
rect 41804 29538 41860 29932
rect 41804 29486 41806 29538
rect 41858 29486 41860 29538
rect 41804 29474 41860 29486
rect 41692 28140 41860 28196
rect 41692 27972 41748 28010
rect 41692 27906 41748 27916
rect 41580 27806 41582 27858
rect 41634 27806 41636 27858
rect 41580 27794 41636 27806
rect 41804 27860 41860 28140
rect 41804 27794 41860 27804
rect 41132 26180 41188 26190
rect 41132 26068 41188 26124
rect 40236 24658 40292 24668
rect 40796 26012 41188 26068
rect 38332 24558 38334 24610
rect 38386 24558 38388 24610
rect 38332 24546 38388 24558
rect 40348 24612 40404 24622
rect 40796 24612 40852 26012
rect 41244 25956 41300 26796
rect 41580 27636 41636 27646
rect 41580 27188 41636 27580
rect 41580 26516 41636 27132
rect 41692 27634 41748 27646
rect 41692 27582 41694 27634
rect 41746 27582 41748 27634
rect 41692 26964 41748 27582
rect 41804 27300 41860 27310
rect 41804 27186 41860 27244
rect 41804 27134 41806 27186
rect 41858 27134 41860 27186
rect 41804 27122 41860 27134
rect 41692 26908 41860 26964
rect 41692 26516 41748 26526
rect 41580 26514 41748 26516
rect 41580 26462 41694 26514
rect 41746 26462 41748 26514
rect 41580 26460 41748 26462
rect 41692 26450 41748 26460
rect 41804 26402 41860 26908
rect 41804 26350 41806 26402
rect 41858 26350 41860 26402
rect 41804 26338 41860 26350
rect 40908 25900 41300 25956
rect 41468 26290 41524 26302
rect 41468 26238 41470 26290
rect 41522 26238 41524 26290
rect 40908 25508 40964 25900
rect 40908 25506 41076 25508
rect 40908 25454 40910 25506
rect 40962 25454 41076 25506
rect 40908 25452 41076 25454
rect 40908 25442 40964 25452
rect 40908 25060 40964 25070
rect 40908 24834 40964 25004
rect 41020 24946 41076 25452
rect 41020 24894 41022 24946
rect 41074 24894 41076 24946
rect 41020 24882 41076 24894
rect 41132 25284 41188 25294
rect 41468 25284 41524 26238
rect 41132 25282 41524 25284
rect 41132 25230 41134 25282
rect 41186 25230 41524 25282
rect 41132 25228 41524 25230
rect 41132 25172 41188 25228
rect 40908 24782 40910 24834
rect 40962 24782 40964 24834
rect 40908 24770 40964 24782
rect 40908 24612 40964 24622
rect 40796 24556 40908 24612
rect 39452 22148 39508 22158
rect 39004 21476 39060 21486
rect 38780 21474 39060 21476
rect 38780 21422 39006 21474
rect 39058 21422 39060 21474
rect 38780 21420 39060 21422
rect 37548 20804 37604 20814
rect 37548 20710 37604 20748
rect 38780 20804 38836 21420
rect 39004 21410 39060 21420
rect 39452 21474 39508 22092
rect 39452 21422 39454 21474
rect 39506 21422 39508 21474
rect 37212 20690 37492 20692
rect 37212 20638 37214 20690
rect 37266 20638 37492 20690
rect 37212 20636 37492 20638
rect 37212 20626 37268 20636
rect 36092 20188 36148 20300
rect 35420 20078 35422 20130
rect 35474 20078 35476 20130
rect 35084 19954 35140 19964
rect 35420 19796 35476 20078
rect 35644 20132 35700 20142
rect 35644 20038 35700 20076
rect 35756 20132 36148 20188
rect 37548 20132 37604 20142
rect 35420 19740 35588 19796
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35420 19348 35476 19358
rect 35532 19348 35588 19740
rect 35420 19346 35588 19348
rect 35420 19294 35422 19346
rect 35474 19294 35588 19346
rect 35420 19292 35588 19294
rect 35420 19282 35476 19292
rect 34076 19236 34132 19246
rect 33628 19234 34132 19236
rect 33628 19182 34078 19234
rect 34130 19182 34132 19234
rect 33628 19180 34132 19182
rect 33180 18340 33236 18350
rect 33180 18246 33236 18284
rect 32956 17220 33012 17230
rect 32956 16996 33012 17164
rect 32956 16930 33012 16940
rect 33180 17108 33236 17118
rect 33180 16884 33236 17052
rect 33516 16884 33572 16894
rect 33180 16882 33572 16884
rect 33180 16830 33182 16882
rect 33234 16830 33518 16882
rect 33570 16830 33572 16882
rect 33180 16828 33572 16830
rect 33180 16818 33236 16828
rect 33516 16818 33572 16828
rect 33628 16660 33684 19180
rect 34076 19170 34132 19180
rect 33404 16604 33684 16660
rect 34636 19122 34692 19134
rect 34636 19070 34638 19122
rect 34690 19070 34692 19122
rect 32396 14924 32676 14980
rect 32732 16212 32788 16222
rect 31836 14868 31892 14878
rect 31836 14644 31892 14812
rect 31724 14588 32116 14644
rect 31724 14530 31780 14588
rect 31724 14478 31726 14530
rect 31778 14478 31780 14530
rect 31724 14466 31780 14478
rect 31388 14366 31390 14418
rect 31442 14366 31444 14418
rect 28812 13860 28868 13870
rect 26348 13806 26350 13858
rect 26402 13806 26404 13858
rect 26348 13794 26404 13806
rect 28700 13858 28868 13860
rect 28700 13806 28814 13858
rect 28866 13806 28868 13858
rect 28700 13804 28868 13806
rect 26236 13694 26238 13746
rect 26290 13694 26292 13746
rect 26236 13682 26292 13694
rect 28364 13748 28420 13758
rect 28364 13746 28532 13748
rect 28364 13694 28366 13746
rect 28418 13694 28532 13746
rect 28364 13692 28532 13694
rect 28364 13682 28420 13692
rect 28476 13412 28532 13692
rect 28476 13356 28644 13412
rect 26012 11282 26068 11294
rect 26012 11230 26014 11282
rect 26066 11230 26068 11282
rect 25788 10836 25844 10846
rect 25676 10834 25844 10836
rect 25676 10782 25790 10834
rect 25842 10782 25844 10834
rect 25676 10780 25844 10782
rect 25564 10742 25620 10780
rect 25788 10770 25844 10780
rect 25340 10724 25396 10734
rect 25340 10630 25396 10668
rect 26012 10724 26068 11230
rect 26348 11284 26404 11294
rect 26348 11190 26404 11228
rect 26124 11170 26180 11182
rect 26124 11118 26126 11170
rect 26178 11118 26180 11170
rect 26124 10836 26180 11118
rect 26124 10770 26180 10780
rect 26684 10836 26740 10846
rect 26684 10742 26740 10780
rect 26012 10658 26068 10668
rect 27020 10724 27076 10734
rect 27020 10630 27076 10668
rect 28588 10724 28644 13356
rect 25116 10332 25284 10388
rect 25452 10498 25508 10510
rect 25452 10446 25454 10498
rect 25506 10446 25508 10498
rect 24892 9940 24948 9950
rect 24892 9846 24948 9884
rect 24780 9774 24782 9826
rect 24834 9774 24836 9826
rect 23996 9268 24052 9278
rect 24780 9268 24836 9774
rect 25116 9826 25172 10332
rect 25116 9774 25118 9826
rect 25170 9774 25172 9826
rect 25116 9762 25172 9774
rect 25340 9828 25396 9838
rect 25452 9828 25508 10446
rect 26460 9940 26516 9950
rect 26460 9846 26516 9884
rect 28588 9938 28644 10668
rect 28588 9886 28590 9938
rect 28642 9886 28644 9938
rect 28588 9874 28644 9886
rect 25788 9828 25844 9838
rect 25340 9826 25508 9828
rect 25340 9774 25342 9826
rect 25394 9774 25508 9826
rect 25340 9772 25508 9774
rect 25564 9772 25788 9828
rect 25340 9762 25396 9772
rect 24052 9212 24388 9268
rect 24780 9212 25172 9268
rect 23996 9174 24052 9212
rect 24332 9154 24388 9212
rect 24332 9102 24334 9154
rect 24386 9102 24388 9154
rect 24332 9090 24388 9102
rect 24556 9156 24612 9166
rect 24556 9062 24612 9100
rect 25004 9044 25060 9054
rect 24668 8932 24724 8942
rect 24668 8838 24724 8876
rect 25004 8370 25060 8988
rect 25116 9042 25172 9212
rect 25116 8990 25118 9042
rect 25170 8990 25172 9042
rect 25116 8978 25172 8990
rect 25452 9042 25508 9054
rect 25452 8990 25454 9042
rect 25506 8990 25508 9042
rect 25452 8932 25508 8990
rect 25452 8866 25508 8876
rect 25004 8318 25006 8370
rect 25058 8318 25060 8370
rect 25004 8306 25060 8318
rect 21644 6690 21812 6692
rect 21644 6638 21646 6690
rect 21698 6638 21812 6690
rect 21644 6636 21812 6638
rect 21644 6626 21700 6636
rect 21756 6468 21812 6478
rect 21756 6374 21812 6412
rect 23436 6468 23492 6478
rect 21084 6018 21588 6020
rect 21084 5966 21086 6018
rect 21138 5966 21588 6018
rect 21084 5964 21588 5966
rect 21084 5236 21140 5964
rect 22204 5906 22260 5918
rect 22204 5854 22206 5906
rect 22258 5854 22260 5906
rect 21308 5236 21364 5246
rect 21084 5234 21364 5236
rect 21084 5182 21310 5234
rect 21362 5182 21364 5234
rect 21084 5180 21364 5182
rect 21308 5170 21364 5180
rect 20412 4946 20468 4956
rect 22204 5012 22260 5854
rect 23436 5234 23492 6412
rect 25340 5908 25396 5918
rect 25564 5908 25620 9772
rect 25788 9734 25844 9772
rect 28700 9716 28756 13804
rect 28812 13794 28868 13804
rect 31388 13522 31444 14366
rect 31388 13470 31390 13522
rect 31442 13470 31444 13522
rect 31388 13458 31444 13470
rect 31500 14364 31668 14420
rect 31948 14418 32004 14430
rect 31948 14366 31950 14418
rect 32002 14366 32004 14418
rect 31500 11620 31556 14364
rect 31948 13970 32004 14366
rect 31948 13918 31950 13970
rect 32002 13918 32004 13970
rect 31948 13906 32004 13918
rect 31612 13748 31668 13758
rect 31836 13748 31892 13758
rect 31612 13654 31668 13692
rect 31724 13746 31892 13748
rect 31724 13694 31838 13746
rect 31890 13694 31892 13746
rect 31724 13692 31892 13694
rect 31612 13524 31668 13534
rect 31724 13524 31780 13692
rect 31836 13682 31892 13692
rect 32060 13746 32116 14588
rect 32060 13694 32062 13746
rect 32114 13694 32116 13746
rect 31612 13522 31780 13524
rect 31612 13470 31614 13522
rect 31666 13470 31780 13522
rect 31612 13468 31780 13470
rect 31612 13458 31668 13468
rect 31612 11620 31668 11630
rect 31500 11564 31612 11620
rect 31612 11554 31668 11564
rect 31612 11396 31668 11406
rect 31612 11302 31668 11340
rect 31276 11282 31332 11294
rect 31276 11230 31278 11282
rect 31330 11230 31332 11282
rect 31276 11060 31332 11230
rect 31500 11172 31556 11182
rect 31500 11170 31668 11172
rect 31500 11118 31502 11170
rect 31554 11118 31668 11170
rect 31500 11116 31668 11118
rect 31500 11106 31556 11116
rect 31276 10994 31332 11004
rect 29708 10836 29764 10846
rect 29708 10612 29764 10780
rect 28140 9660 28756 9716
rect 29260 10610 29764 10612
rect 29260 10558 29710 10610
rect 29762 10558 29764 10610
rect 29260 10556 29764 10558
rect 29260 9938 29316 10556
rect 29708 10546 29764 10556
rect 30380 10498 30436 10510
rect 30380 10446 30382 10498
rect 30434 10446 30436 10498
rect 30380 10052 30436 10446
rect 31276 10052 31332 10062
rect 30380 10050 31332 10052
rect 30380 9998 31278 10050
rect 31330 9998 31332 10050
rect 30380 9996 31332 9998
rect 31276 9986 31332 9996
rect 31612 10050 31668 11116
rect 31724 11060 31780 13468
rect 31948 11620 32004 11630
rect 31836 11508 31892 11518
rect 31836 11394 31892 11452
rect 31836 11342 31838 11394
rect 31890 11342 31892 11394
rect 31836 11330 31892 11342
rect 31724 10994 31780 11004
rect 31948 11172 32004 11564
rect 32060 11396 32116 13694
rect 32396 13748 32452 14924
rect 32732 14644 32788 16156
rect 33404 15538 33460 16604
rect 33404 15486 33406 15538
rect 33458 15486 33460 15538
rect 33068 15426 33124 15438
rect 33068 15374 33070 15426
rect 33122 15374 33124 15426
rect 33068 14868 33124 15374
rect 33404 15204 33460 15486
rect 33404 15138 33460 15148
rect 33068 14802 33124 14812
rect 32396 13654 32452 13692
rect 32508 14642 32788 14644
rect 32508 14590 32734 14642
rect 32786 14590 32788 14642
rect 32508 14588 32788 14590
rect 32060 11330 32116 11340
rect 32396 11508 32452 11518
rect 32172 11172 32228 11182
rect 31948 11170 32228 11172
rect 31948 11118 32174 11170
rect 32226 11118 32228 11170
rect 31948 11116 32228 11118
rect 31948 10948 32004 11116
rect 32172 11106 32228 11116
rect 31612 9998 31614 10050
rect 31666 9998 31668 10050
rect 31612 9986 31668 9998
rect 31836 10892 32004 10948
rect 29260 9886 29262 9938
rect 29314 9886 29316 9938
rect 29260 9828 29316 9886
rect 25900 9604 25956 9614
rect 25676 9044 25732 9054
rect 25676 8950 25732 8988
rect 25900 9042 25956 9548
rect 26124 9156 26180 9166
rect 26460 9156 26516 9166
rect 26180 9154 26516 9156
rect 26180 9102 26462 9154
rect 26514 9102 26516 9154
rect 26180 9100 26516 9102
rect 26124 9062 26180 9100
rect 26460 9090 26516 9100
rect 26572 9156 26628 9166
rect 26572 9062 26628 9100
rect 28140 9156 28196 9660
rect 25900 8990 25902 9042
rect 25954 8990 25956 9042
rect 25900 8978 25956 8990
rect 26012 8930 26068 8942
rect 26012 8878 26014 8930
rect 26066 8878 26068 8930
rect 26012 6018 26068 8878
rect 26012 5966 26014 6018
rect 26066 5966 26068 6018
rect 26012 5954 26068 5966
rect 23436 5182 23438 5234
rect 23490 5182 23492 5234
rect 23436 5170 23492 5182
rect 24780 5906 25620 5908
rect 24780 5854 25342 5906
rect 25394 5854 25620 5906
rect 24780 5852 25620 5854
rect 24780 5234 24836 5852
rect 25340 5842 25396 5852
rect 28140 5794 28196 9100
rect 29260 8428 29316 9772
rect 31388 9826 31444 9838
rect 31388 9774 31390 9826
rect 31442 9774 31444 9826
rect 30940 9604 30996 9614
rect 31388 9604 31444 9774
rect 31836 9826 31892 10892
rect 32396 10500 32452 11452
rect 32508 10836 32564 14588
rect 32732 14578 32788 14588
rect 32732 11396 32788 11406
rect 32732 11302 32788 11340
rect 32956 11396 33012 11406
rect 32956 11302 33012 11340
rect 34636 11396 34692 19070
rect 35756 18450 35812 20132
rect 35980 20020 36036 20030
rect 35980 19926 36036 19964
rect 37548 19348 37604 20076
rect 38780 19460 38836 20748
rect 38892 20356 38948 20366
rect 39452 20356 39508 21422
rect 38948 20300 39508 20356
rect 38892 20290 38948 20300
rect 39004 20020 39060 20030
rect 38892 19460 38948 19470
rect 35756 18398 35758 18450
rect 35810 18398 35812 18450
rect 35756 18340 35812 18398
rect 37324 19346 37604 19348
rect 37324 19294 37550 19346
rect 37602 19294 37604 19346
rect 37324 19292 37604 19294
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 34860 16884 34916 16894
rect 34860 15314 34916 16828
rect 35756 16884 35812 18284
rect 36540 18338 36596 18350
rect 36540 18286 36542 18338
rect 36594 18286 36596 18338
rect 36540 17892 36596 18286
rect 36988 17892 37044 17902
rect 36540 17890 37044 17892
rect 36540 17838 36990 17890
rect 37042 17838 37044 17890
rect 36540 17836 37044 17838
rect 36988 17826 37044 17836
rect 37324 17890 37380 19292
rect 37548 19282 37604 19292
rect 38556 19458 38948 19460
rect 38556 19406 38894 19458
rect 38946 19406 38948 19458
rect 38556 19404 38948 19406
rect 37996 19236 38052 19246
rect 37996 19142 38052 19180
rect 38332 19236 38388 19246
rect 38556 19236 38612 19404
rect 38892 19394 38948 19404
rect 38332 19234 38612 19236
rect 38332 19182 38334 19234
rect 38386 19182 38612 19234
rect 38332 19180 38612 19182
rect 38668 19236 38724 19246
rect 38332 19170 38388 19180
rect 38668 18338 38724 19180
rect 38668 18286 38670 18338
rect 38722 18286 38724 18338
rect 38668 18274 38724 18286
rect 37324 17838 37326 17890
rect 37378 17838 37380 17890
rect 37324 17826 37380 17838
rect 37100 17666 37156 17678
rect 37100 17614 37102 17666
rect 37154 17614 37156 17666
rect 36428 17442 36484 17454
rect 36428 17390 36430 17442
rect 36482 17390 36484 17442
rect 36428 17220 36484 17390
rect 35756 16818 35812 16828
rect 36316 17164 36428 17220
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34860 15262 34862 15314
rect 34914 15262 34916 15314
rect 34860 15250 34916 15262
rect 35532 15204 35588 15214
rect 35532 15202 36036 15204
rect 35532 15150 35534 15202
rect 35586 15150 36036 15202
rect 35532 15148 36036 15150
rect 35532 15138 35588 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35756 13972 35812 13982
rect 35980 13972 36036 15148
rect 36092 14308 36148 14318
rect 36092 14306 36260 14308
rect 36092 14254 36094 14306
rect 36146 14254 36260 14306
rect 36092 14252 36260 14254
rect 36092 14242 36148 14252
rect 36092 13972 36148 13982
rect 35980 13970 36148 13972
rect 35980 13918 36094 13970
rect 36146 13918 36148 13970
rect 35980 13916 36148 13918
rect 35756 13748 35812 13916
rect 36092 13906 36148 13916
rect 35756 13654 35812 13692
rect 35868 13860 35924 13870
rect 35868 13746 35924 13804
rect 35868 13694 35870 13746
rect 35922 13694 35924 13746
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34636 11330 34692 11340
rect 35868 11394 35924 13694
rect 35868 11342 35870 11394
rect 35922 11342 35924 11394
rect 35868 11330 35924 11342
rect 36204 13746 36260 14252
rect 36204 13694 36206 13746
rect 36258 13694 36260 13746
rect 36204 13636 36260 13694
rect 36204 11396 36260 13580
rect 36204 11302 36260 11340
rect 32620 11282 32676 11294
rect 32620 11230 32622 11282
rect 32674 11230 32676 11282
rect 32620 11172 32676 11230
rect 32620 11106 32676 11116
rect 34188 11170 34244 11182
rect 34188 11118 34190 11170
rect 34242 11118 34244 11170
rect 34188 11060 34244 11118
rect 34524 11172 34580 11182
rect 34524 11078 34580 11116
rect 35980 11170 36036 11182
rect 35980 11118 35982 11170
rect 36034 11118 36036 11170
rect 34188 10994 34244 11004
rect 35756 11060 35812 11070
rect 32508 10770 32564 10780
rect 33180 10836 33236 10846
rect 33180 10742 33236 10780
rect 35084 10836 35140 10846
rect 35084 10742 35140 10780
rect 35532 10836 35588 10846
rect 35532 10610 35588 10780
rect 35532 10558 35534 10610
rect 35586 10558 35588 10610
rect 35532 10546 35588 10558
rect 35756 10610 35812 11004
rect 35756 10558 35758 10610
rect 35810 10558 35812 10610
rect 35756 10546 35812 10558
rect 35868 10834 35924 10846
rect 35868 10782 35870 10834
rect 35922 10782 35924 10834
rect 32508 10500 32564 10510
rect 32396 10498 32564 10500
rect 32396 10446 32510 10498
rect 32562 10446 32564 10498
rect 32396 10444 32564 10446
rect 32508 10434 32564 10444
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 31836 9774 31838 9826
rect 31890 9774 31892 9826
rect 31836 9762 31892 9774
rect 30940 9602 31388 9604
rect 30940 9550 30942 9602
rect 30994 9550 31388 9602
rect 30940 9548 31388 9550
rect 30940 9044 30996 9548
rect 31388 9510 31444 9548
rect 35756 9156 35812 9166
rect 35868 9156 35924 10782
rect 35980 10610 36036 11118
rect 36316 10836 36372 17164
rect 36428 17154 36484 17164
rect 37100 17220 37156 17614
rect 37548 17668 37604 17678
rect 37548 17574 37604 17612
rect 37100 17154 37156 17164
rect 38108 16884 38164 16894
rect 38108 16770 38164 16828
rect 38108 16718 38110 16770
rect 38162 16718 38164 16770
rect 37660 15202 37716 15214
rect 37660 15150 37662 15202
rect 37714 15150 37716 15202
rect 36428 14532 36484 14542
rect 36428 14438 36484 14476
rect 37548 14530 37604 14542
rect 37548 14478 37550 14530
rect 37602 14478 37604 14530
rect 36764 13972 36820 13982
rect 36540 13748 36596 13758
rect 36540 13654 36596 13692
rect 36764 13746 36820 13916
rect 37436 13860 37492 13870
rect 37436 13766 37492 13804
rect 36764 13694 36766 13746
rect 36818 13694 36820 13746
rect 36764 13682 36820 13694
rect 37212 13746 37268 13758
rect 37212 13694 37214 13746
rect 37266 13694 37268 13746
rect 37212 13636 37268 13694
rect 37324 13748 37380 13758
rect 37324 13654 37380 13692
rect 37212 13570 37268 13580
rect 37548 13188 37604 14478
rect 37660 14532 37716 15150
rect 38108 15204 38164 16718
rect 38108 15202 38276 15204
rect 38108 15150 38110 15202
rect 38162 15150 38276 15202
rect 38108 15148 38276 15150
rect 38108 15138 38164 15148
rect 37660 14418 37716 14476
rect 37660 14366 37662 14418
rect 37714 14366 37716 14418
rect 37660 14354 37716 14366
rect 37996 13860 38052 13870
rect 38052 13804 38164 13860
rect 37996 13794 38052 13804
rect 37548 13132 37828 13188
rect 37660 12964 37716 12974
rect 37660 12402 37716 12908
rect 37660 12350 37662 12402
rect 37714 12350 37716 12402
rect 37660 12338 37716 12350
rect 37436 12178 37492 12190
rect 37772 12180 37828 13132
rect 37436 12126 37438 12178
rect 37490 12126 37492 12178
rect 37100 12068 37156 12078
rect 37436 12068 37492 12126
rect 37660 12124 37828 12180
rect 38108 12290 38164 13804
rect 38108 12238 38110 12290
rect 38162 12238 38164 12290
rect 37100 12066 37492 12068
rect 37100 12014 37102 12066
rect 37154 12014 37492 12066
rect 37100 12012 37492 12014
rect 37548 12068 37604 12078
rect 36428 11508 36484 11518
rect 36428 11394 36484 11452
rect 36428 11342 36430 11394
rect 36482 11342 36484 11394
rect 36428 11330 36484 11342
rect 36988 11172 37044 11182
rect 36988 11078 37044 11116
rect 36316 10770 36372 10780
rect 35980 10558 35982 10610
rect 36034 10558 36036 10610
rect 35980 10546 36036 10558
rect 37100 9604 37156 12012
rect 37548 11732 37604 12012
rect 37436 11676 37604 11732
rect 37436 11394 37492 11676
rect 37660 11508 37716 12124
rect 37772 11956 37828 11966
rect 38108 11956 38164 12238
rect 37772 11954 38164 11956
rect 37772 11902 37774 11954
rect 37826 11902 38164 11954
rect 37772 11900 38164 11902
rect 37772 11890 37828 11900
rect 37436 11342 37438 11394
rect 37490 11342 37492 11394
rect 37436 11330 37492 11342
rect 37548 11396 37604 11406
rect 37548 11302 37604 11340
rect 37660 11396 37716 11452
rect 37660 11394 37940 11396
rect 37660 11342 37662 11394
rect 37714 11342 37940 11394
rect 37660 11340 37940 11342
rect 37660 11330 37716 11340
rect 37100 9538 37156 9548
rect 35756 9154 35924 9156
rect 35756 9102 35758 9154
rect 35810 9102 35924 9154
rect 35756 9100 35924 9102
rect 35756 9090 35812 9100
rect 30940 8978 30996 8988
rect 35084 9044 35140 9054
rect 35084 8950 35140 8988
rect 37884 8930 37940 11340
rect 38220 9044 38276 15148
rect 39004 14306 39060 19964
rect 39116 18452 39172 20300
rect 39228 19010 39284 19022
rect 39228 18958 39230 19010
rect 39282 18958 39284 19010
rect 39228 18564 39284 18958
rect 39228 18508 39732 18564
rect 39116 18450 39620 18452
rect 39116 18398 39118 18450
rect 39170 18398 39620 18450
rect 39116 18396 39620 18398
rect 39116 18386 39172 18396
rect 39564 17780 39620 18396
rect 39564 17686 39620 17724
rect 39676 17668 39732 18508
rect 40348 18340 40404 24556
rect 40908 24052 40964 24556
rect 40908 23958 40964 23996
rect 41132 23940 41188 25116
rect 41244 24724 41300 24734
rect 41244 24722 41636 24724
rect 41244 24670 41246 24722
rect 41298 24670 41636 24722
rect 41244 24668 41636 24670
rect 41244 24658 41300 24668
rect 41468 24500 41524 24510
rect 41244 23940 41300 23950
rect 41132 23938 41300 23940
rect 41132 23886 41246 23938
rect 41298 23886 41300 23938
rect 41132 23884 41300 23886
rect 41244 23874 41300 23884
rect 41468 23826 41524 24444
rect 41468 23774 41470 23826
rect 41522 23774 41524 23826
rect 41468 23762 41524 23774
rect 41580 23826 41636 24668
rect 41916 24500 41972 32060
rect 43596 30324 43652 30334
rect 43596 30230 43652 30268
rect 42252 27746 42308 27758
rect 42252 27694 42254 27746
rect 42306 27694 42308 27746
rect 42140 27634 42196 27646
rect 42140 27582 42142 27634
rect 42194 27582 42196 27634
rect 42140 27300 42196 27582
rect 42140 27234 42196 27244
rect 42028 26402 42084 26414
rect 42028 26350 42030 26402
rect 42082 26350 42084 26402
rect 42028 26180 42084 26350
rect 42028 26114 42084 26124
rect 42252 26178 42308 27694
rect 43932 27188 43988 27198
rect 43932 27094 43988 27132
rect 42252 26126 42254 26178
rect 42306 26126 42308 26178
rect 42252 26114 42308 26126
rect 41916 24434 41972 24444
rect 43708 24500 43764 24510
rect 41580 23774 41582 23826
rect 41634 23774 41636 23826
rect 41580 23762 41636 23774
rect 41692 24052 41748 24062
rect 41692 23826 41748 23996
rect 41692 23774 41694 23826
rect 41746 23774 41748 23826
rect 41692 23762 41748 23774
rect 41356 23714 41412 23726
rect 41356 23662 41358 23714
rect 41410 23662 41412 23714
rect 41356 23380 41412 23662
rect 41356 23324 41860 23380
rect 41804 23266 41860 23324
rect 41804 23214 41806 23266
rect 41858 23214 41860 23266
rect 41804 23202 41860 23214
rect 41692 22932 41748 22942
rect 41580 22930 41748 22932
rect 41580 22878 41694 22930
rect 41746 22878 41748 22930
rect 41580 22876 41748 22878
rect 41580 22482 41636 22876
rect 41692 22866 41748 22876
rect 41580 22430 41582 22482
rect 41634 22430 41636 22482
rect 41580 22418 41636 22430
rect 43708 22482 43764 24444
rect 43708 22430 43710 22482
rect 43762 22430 43764 22482
rect 43708 22418 43764 22430
rect 40908 22370 40964 22382
rect 40908 22318 40910 22370
rect 40962 22318 40964 22370
rect 40460 22148 40516 22158
rect 40460 22054 40516 22092
rect 40908 22148 40964 22318
rect 40908 22082 40964 22092
rect 41804 18450 41860 18462
rect 41804 18398 41806 18450
rect 41858 18398 41860 18450
rect 40012 18284 40516 18340
rect 39676 16996 39732 17612
rect 39676 16930 39732 16940
rect 39900 17780 39956 17790
rect 39004 14254 39006 14306
rect 39058 14254 39060 14306
rect 39004 14242 39060 14254
rect 39900 13972 39956 17724
rect 40012 17778 40068 18284
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 40012 17714 40068 17726
rect 40348 17554 40404 17566
rect 40348 17502 40350 17554
rect 40402 17502 40404 17554
rect 40236 17108 40292 17118
rect 40236 17014 40292 17052
rect 40124 16996 40180 17006
rect 40124 16902 40180 16940
rect 40348 16884 40404 17502
rect 40460 17554 40516 18284
rect 41692 18338 41748 18350
rect 41692 18286 41694 18338
rect 41746 18286 41748 18338
rect 41468 18228 41524 18238
rect 40684 18226 41524 18228
rect 40684 18174 41470 18226
rect 41522 18174 41524 18226
rect 40684 18172 41524 18174
rect 40684 17666 40740 18172
rect 41468 18162 41524 18172
rect 40684 17614 40686 17666
rect 40738 17614 40740 17666
rect 40684 17602 40740 17614
rect 40908 17780 40964 17790
rect 41580 17780 41636 17790
rect 40908 17666 40964 17724
rect 40908 17614 40910 17666
rect 40962 17614 40964 17666
rect 40908 17602 40964 17614
rect 41468 17724 41580 17780
rect 40460 17502 40462 17554
rect 40514 17502 40516 17554
rect 40460 17490 40516 17502
rect 41468 17108 41524 17724
rect 41580 17714 41636 17724
rect 41692 17778 41748 18286
rect 41692 17726 41694 17778
rect 41746 17726 41748 17778
rect 41692 17714 41748 17726
rect 41244 16996 41300 17006
rect 41244 16902 41300 16940
rect 40460 16884 40516 16894
rect 40348 16882 40516 16884
rect 40348 16830 40462 16882
rect 40514 16830 40516 16882
rect 40348 16828 40516 16830
rect 39900 13878 39956 13916
rect 40348 13636 40404 13646
rect 40348 13542 40404 13580
rect 40236 13522 40292 13534
rect 40236 13470 40238 13522
rect 40290 13470 40292 13522
rect 38444 13076 38500 13086
rect 38444 12402 38500 13020
rect 40124 13076 40180 13086
rect 40124 12982 40180 13020
rect 38444 12350 38446 12402
rect 38498 12350 38500 12402
rect 38444 12068 38500 12350
rect 40236 12850 40292 13470
rect 40236 12798 40238 12850
rect 40290 12798 40292 12850
rect 40236 12404 40292 12798
rect 40236 12338 40292 12348
rect 40460 12850 40516 16828
rect 41468 14644 41524 17052
rect 41804 16996 41860 18398
rect 43820 17780 43876 17790
rect 43820 17686 43876 17724
rect 41580 16940 41860 16996
rect 41580 16770 41636 16940
rect 41580 16718 41582 16770
rect 41634 16718 41636 16770
rect 41580 16706 41636 16718
rect 41244 14588 41524 14644
rect 41244 14530 41300 14588
rect 41244 14478 41246 14530
rect 41298 14478 41300 14530
rect 41244 14466 41300 14478
rect 41356 14418 41412 14430
rect 41356 14366 41358 14418
rect 41410 14366 41412 14418
rect 41020 13972 41076 13982
rect 41020 13746 41076 13916
rect 41020 13694 41022 13746
rect 41074 13694 41076 13746
rect 41020 13682 41076 13694
rect 41356 13636 41412 14366
rect 41356 13570 41412 13580
rect 41804 13636 41860 13646
rect 43932 13636 43988 13646
rect 41804 13634 41972 13636
rect 41804 13582 41806 13634
rect 41858 13582 41972 13634
rect 41804 13580 41972 13582
rect 41804 13570 41860 13580
rect 40460 12798 40462 12850
rect 40514 12798 40516 12850
rect 40460 12180 40516 12798
rect 40796 12962 40852 12974
rect 40796 12910 40798 12962
rect 40850 12910 40852 12962
rect 40796 12402 40852 12910
rect 41020 12964 41076 12974
rect 41020 12870 41076 12908
rect 41356 12852 41412 12862
rect 41692 12852 41748 12862
rect 41356 12850 41748 12852
rect 41356 12798 41358 12850
rect 41410 12798 41694 12850
rect 41746 12798 41748 12850
rect 41356 12796 41748 12798
rect 41916 12852 41972 13580
rect 43932 13542 43988 13580
rect 42028 12852 42084 12862
rect 41916 12850 42084 12852
rect 41916 12798 42030 12850
rect 42082 12798 42084 12850
rect 41916 12796 42084 12798
rect 41356 12786 41412 12796
rect 41692 12786 41748 12796
rect 42028 12786 42084 12796
rect 40796 12350 40798 12402
rect 40850 12350 40852 12402
rect 40796 12338 40852 12350
rect 41020 12404 41076 12414
rect 41020 12310 41076 12348
rect 41132 12180 41188 12190
rect 40460 12178 41188 12180
rect 40460 12126 41134 12178
rect 41186 12126 41188 12178
rect 40460 12124 41188 12126
rect 41132 12114 41188 12124
rect 38444 12002 38500 12012
rect 38332 9044 38388 9054
rect 38220 8988 38332 9044
rect 38332 8950 38388 8988
rect 37884 8878 37886 8930
rect 37938 8878 37940 8930
rect 37884 8866 37940 8878
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 28700 8372 29316 8428
rect 28588 6132 28644 6142
rect 28700 6132 28756 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 28588 6130 28756 6132
rect 28588 6078 28590 6130
rect 28642 6078 28756 6130
rect 28588 6076 28756 6078
rect 28588 6066 28644 6076
rect 28140 5742 28142 5794
rect 28194 5742 28196 5794
rect 28140 5730 28196 5742
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 24780 5182 24782 5234
rect 24834 5182 24836 5234
rect 24108 5124 24164 5134
rect 24108 5030 24164 5068
rect 24780 5124 24836 5182
rect 24780 5058 24836 5068
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4508 19908 4564
rect 19180 4338 19236 4508
rect 19852 4450 19908 4508
rect 19852 4398 19854 4450
rect 19906 4398 19908 4450
rect 19852 4386 19908 4398
rect 19180 4286 19182 4338
rect 19234 4286 19236 4338
rect 19180 4274 19236 4286
rect 16380 4174 16382 4226
rect 16434 4174 16436 4226
rect 16380 4162 16436 4174
rect 21980 4228 22036 4238
rect 22204 4228 22260 4956
rect 21980 4226 22260 4228
rect 21980 4174 21982 4226
rect 22034 4174 22260 4226
rect 21980 4172 22260 4174
rect 21980 4162 22036 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
<< via2 >>
rect 1932 33964 1988 34020
rect 2156 31500 2212 31556
rect 1932 22204 1988 22260
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5180 40908 5236 40964
rect 3276 40348 3332 40404
rect 5180 40348 5236 40404
rect 3724 40290 3780 40292
rect 3724 40238 3726 40290
rect 3726 40238 3778 40290
rect 3778 40238 3780 40290
rect 3724 40236 3780 40238
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 6300 40908 6356 40964
rect 6188 40348 6244 40404
rect 8092 40460 8148 40516
rect 5852 40124 5908 40180
rect 6412 40236 6468 40292
rect 6972 39452 7028 39508
rect 7644 39506 7700 39508
rect 7644 39454 7646 39506
rect 7646 39454 7698 39506
rect 7698 39454 7700 39506
rect 7644 39452 7700 39454
rect 6300 39394 6356 39396
rect 6300 39342 6302 39394
rect 6302 39342 6354 39394
rect 6354 39342 6356 39394
rect 6300 39340 6356 39342
rect 2604 38946 2660 38948
rect 2604 38894 2606 38946
rect 2606 38894 2658 38946
rect 2658 38894 2660 38946
rect 2604 38892 2660 38894
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 2604 35810 2660 35812
rect 2604 35758 2606 35810
rect 2606 35758 2658 35810
rect 2658 35758 2660 35810
rect 2604 35756 2660 35758
rect 4732 35420 4788 35476
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4844 34972 4900 35028
rect 4956 36204 5012 36260
rect 7532 39394 7588 39396
rect 7532 39342 7534 39394
rect 7534 39342 7586 39394
rect 7586 39342 7588 39394
rect 7532 39340 7588 39342
rect 7308 39004 7364 39060
rect 7868 39004 7924 39060
rect 4284 33964 4340 34020
rect 7196 36258 7252 36260
rect 7196 36206 7198 36258
rect 7198 36206 7250 36258
rect 7250 36206 7252 36258
rect 7196 36204 7252 36206
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 13244 41916 13300 41972
rect 10780 40908 10836 40964
rect 10444 40626 10500 40628
rect 10444 40574 10446 40626
rect 10446 40574 10498 40626
rect 10498 40574 10500 40626
rect 10444 40572 10500 40574
rect 10220 40514 10276 40516
rect 10220 40462 10222 40514
rect 10222 40462 10274 40514
rect 10274 40462 10276 40514
rect 10220 40460 10276 40462
rect 8764 40348 8820 40404
rect 8316 39394 8372 39396
rect 8316 39342 8318 39394
rect 8318 39342 8370 39394
rect 8370 39342 8372 39394
rect 8316 39340 8372 39342
rect 8652 39394 8708 39396
rect 8652 39342 8654 39394
rect 8654 39342 8706 39394
rect 8706 39342 8708 39394
rect 8652 39340 8708 39342
rect 8540 39004 8596 39060
rect 7644 35810 7700 35812
rect 7644 35758 7646 35810
rect 7646 35758 7698 35810
rect 7698 35758 7700 35810
rect 7644 35756 7700 35758
rect 7980 35084 8036 35140
rect 9100 39676 9156 39732
rect 9212 39618 9268 39620
rect 9212 39566 9214 39618
rect 9214 39566 9266 39618
rect 9266 39566 9268 39618
rect 9212 39564 9268 39566
rect 9100 39116 9156 39172
rect 8876 38946 8932 38948
rect 8876 38894 8878 38946
rect 8878 38894 8930 38946
rect 8930 38894 8932 38946
rect 8876 38892 8932 38894
rect 8988 38834 9044 38836
rect 8988 38782 8990 38834
rect 8990 38782 9042 38834
rect 9042 38782 9044 38834
rect 8988 38780 9044 38782
rect 9324 35420 9380 35476
rect 7084 34748 7140 34804
rect 9100 34524 9156 34580
rect 10108 39788 10164 39844
rect 11228 39788 11284 39844
rect 9548 39116 9604 39172
rect 10220 39618 10276 39620
rect 10220 39566 10222 39618
rect 10222 39566 10274 39618
rect 10274 39566 10276 39618
rect 10220 39564 10276 39566
rect 9660 38892 9716 38948
rect 9884 39394 9940 39396
rect 9884 39342 9886 39394
rect 9886 39342 9938 39394
rect 9938 39342 9940 39394
rect 9884 39340 9940 39342
rect 9884 38834 9940 38836
rect 9884 38782 9886 38834
rect 9886 38782 9938 38834
rect 9938 38782 9940 38834
rect 9884 38780 9940 38782
rect 10108 38556 10164 38612
rect 10780 39452 10836 39508
rect 14476 41916 14532 41972
rect 13916 40962 13972 40964
rect 13916 40910 13918 40962
rect 13918 40910 13970 40962
rect 13970 40910 13972 40962
rect 13916 40908 13972 40910
rect 14028 40402 14084 40404
rect 14028 40350 14030 40402
rect 14030 40350 14082 40402
rect 14082 40350 14084 40402
rect 14028 40348 14084 40350
rect 13580 40290 13636 40292
rect 13580 40238 13582 40290
rect 13582 40238 13634 40290
rect 13634 40238 13636 40290
rect 13580 40236 13636 40238
rect 13468 40124 13524 40180
rect 11900 39788 11956 39844
rect 11788 39676 11844 39732
rect 10780 38946 10836 38948
rect 10780 38894 10782 38946
rect 10782 38894 10834 38946
rect 10834 38894 10836 38946
rect 10780 38892 10836 38894
rect 10556 38780 10612 38836
rect 12124 39394 12180 39396
rect 12124 39342 12126 39394
rect 12126 39342 12178 39394
rect 12178 39342 12180 39394
rect 12124 39340 12180 39342
rect 12124 39058 12180 39060
rect 12124 39006 12126 39058
rect 12126 39006 12178 39058
rect 12178 39006 12180 39058
rect 12124 39004 12180 39006
rect 20860 41804 20916 41860
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 17052 40348 17108 40404
rect 17612 40402 17668 40404
rect 17612 40350 17614 40402
rect 17614 40350 17666 40402
rect 17666 40350 17668 40402
rect 17612 40348 17668 40350
rect 19740 40348 19796 40404
rect 18172 39228 18228 39284
rect 13916 39004 13972 39060
rect 11676 38892 11732 38948
rect 11228 38780 11284 38836
rect 9660 36204 9716 36260
rect 10332 35420 10388 35476
rect 11452 37772 11508 37828
rect 10444 35196 10500 35252
rect 10108 34860 10164 34916
rect 10220 34972 10276 35028
rect 5180 33964 5236 34020
rect 7084 34076 7140 34132
rect 9548 34300 9604 34356
rect 7532 34018 7588 34020
rect 7532 33966 7534 34018
rect 7534 33966 7586 34018
rect 7586 33966 7588 34018
rect 7532 33964 7588 33966
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 2940 31666 2996 31668
rect 2940 31614 2942 31666
rect 2942 31614 2994 31666
rect 2994 31614 2996 31666
rect 2940 31612 2996 31614
rect 4172 31612 4228 31668
rect 2604 28812 2660 28868
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5740 31554 5796 31556
rect 5740 31502 5742 31554
rect 5742 31502 5794 31554
rect 5794 31502 5796 31554
rect 5740 31500 5796 31502
rect 7532 31500 7588 31556
rect 7532 30828 7588 30884
rect 6860 29596 6916 29652
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4508 28866 4564 28868
rect 4508 28814 4510 28866
rect 4510 28814 4562 28866
rect 4562 28814 4564 28866
rect 4508 28812 4564 28814
rect 4284 28700 4340 28756
rect 4060 28364 4116 28420
rect 4620 28252 4676 28308
rect 5068 28530 5124 28532
rect 5068 28478 5070 28530
rect 5070 28478 5122 28530
rect 5122 28478 5124 28530
rect 5068 28476 5124 28478
rect 5740 28754 5796 28756
rect 5740 28702 5742 28754
rect 5742 28702 5794 28754
rect 5794 28702 5796 28754
rect 5740 28700 5796 28702
rect 5628 28418 5684 28420
rect 5628 28366 5630 28418
rect 5630 28366 5682 28418
rect 5682 28366 5684 28418
rect 5628 28364 5684 28366
rect 5516 28252 5572 28308
rect 4956 28140 5012 28196
rect 5404 28140 5460 28196
rect 4844 28028 4900 28084
rect 5628 28082 5684 28084
rect 5628 28030 5630 28082
rect 5630 28030 5682 28082
rect 5682 28030 5684 28082
rect 5628 28028 5684 28030
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 6412 28700 6468 28756
rect 6972 28754 7028 28756
rect 6972 28702 6974 28754
rect 6974 28702 7026 28754
rect 7026 28702 7028 28754
rect 6972 28700 7028 28702
rect 7756 28476 7812 28532
rect 5292 26460 5348 26516
rect 5852 26348 5908 26404
rect 4284 26012 4340 26068
rect 4620 26290 4676 26292
rect 4620 26238 4622 26290
rect 4622 26238 4674 26290
rect 4674 26238 4676 26290
rect 4620 26236 4676 26238
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4844 25506 4900 25508
rect 4844 25454 4846 25506
rect 4846 25454 4898 25506
rect 4898 25454 4900 25506
rect 4844 25452 4900 25454
rect 2604 23660 2660 23716
rect 4060 24892 4116 24948
rect 4844 25228 4900 25284
rect 4620 24668 4676 24724
rect 5516 25452 5572 25508
rect 6076 26348 6132 26404
rect 6412 26460 6468 26516
rect 6300 26236 6356 26292
rect 5740 25394 5796 25396
rect 5740 25342 5742 25394
rect 5742 25342 5794 25394
rect 5794 25342 5796 25394
rect 5740 25340 5796 25342
rect 6188 25506 6244 25508
rect 6188 25454 6190 25506
rect 6190 25454 6242 25506
rect 6242 25454 6244 25506
rect 6188 25452 6244 25454
rect 5852 25228 5908 25284
rect 5292 25004 5348 25060
rect 5068 24946 5124 24948
rect 5068 24894 5070 24946
rect 5070 24894 5122 24946
rect 5122 24894 5124 24946
rect 5068 24892 5124 24894
rect 5852 24946 5908 24948
rect 5852 24894 5854 24946
rect 5854 24894 5906 24946
rect 5906 24894 5908 24946
rect 5852 24892 5908 24894
rect 4956 24668 5012 24724
rect 5404 24722 5460 24724
rect 5404 24670 5406 24722
rect 5406 24670 5458 24722
rect 5458 24670 5460 24722
rect 5404 24668 5460 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 3724 23660 3780 23716
rect 3164 23548 3220 23604
rect 2268 22092 2324 22148
rect 6076 24668 6132 24724
rect 6188 25228 6244 25284
rect 6412 25340 6468 25396
rect 6300 24780 6356 24836
rect 6076 23772 6132 23828
rect 6300 23714 6356 23716
rect 6300 23662 6302 23714
rect 6302 23662 6354 23714
rect 6354 23662 6356 23714
rect 6300 23660 6356 23662
rect 6524 23436 6580 23492
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4732 22316 4788 22372
rect 5292 22316 5348 22372
rect 5516 22204 5572 22260
rect 5404 21420 5460 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 6412 21420 6468 21476
rect 7196 25506 7252 25508
rect 7196 25454 7198 25506
rect 7198 25454 7250 25506
rect 7250 25454 7252 25506
rect 7196 25452 7252 25454
rect 7644 24834 7700 24836
rect 7644 24782 7646 24834
rect 7646 24782 7698 24834
rect 7698 24782 7700 24834
rect 7644 24780 7700 24782
rect 8764 27132 8820 27188
rect 8316 25618 8372 25620
rect 8316 25566 8318 25618
rect 8318 25566 8370 25618
rect 8370 25566 8372 25618
rect 8316 25564 8372 25566
rect 7868 24946 7924 24948
rect 7868 24894 7870 24946
rect 7870 24894 7922 24946
rect 7922 24894 7924 24946
rect 7868 24892 7924 24894
rect 7756 24108 7812 24164
rect 7084 23826 7140 23828
rect 7084 23774 7086 23826
rect 7086 23774 7138 23826
rect 7138 23774 7140 23826
rect 7084 23772 7140 23774
rect 7084 22370 7140 22372
rect 7084 22318 7086 22370
rect 7086 22318 7138 22370
rect 7138 22318 7140 22370
rect 7084 22316 7140 22318
rect 6748 21532 6804 21588
rect 7644 22316 7700 22372
rect 8204 25506 8260 25508
rect 8204 25454 8206 25506
rect 8206 25454 8258 25506
rect 8258 25454 8260 25506
rect 8204 25452 8260 25454
rect 9660 30882 9716 30884
rect 9660 30830 9662 30882
rect 9662 30830 9714 30882
rect 9714 30830 9716 30882
rect 9660 30828 9716 30830
rect 9548 28588 9604 28644
rect 10108 34636 10164 34692
rect 11228 35810 11284 35812
rect 11228 35758 11230 35810
rect 11230 35758 11282 35810
rect 11282 35758 11284 35810
rect 11228 35756 11284 35758
rect 12124 37826 12180 37828
rect 12124 37774 12126 37826
rect 12126 37774 12178 37826
rect 12178 37774 12180 37826
rect 12124 37772 12180 37774
rect 20076 40402 20132 40404
rect 20076 40350 20078 40402
rect 20078 40350 20130 40402
rect 20130 40350 20132 40402
rect 20076 40348 20132 40350
rect 23212 41916 23268 41972
rect 22092 41858 22148 41860
rect 22092 41806 22094 41858
rect 22094 41806 22146 41858
rect 22146 41806 22148 41858
rect 22092 41804 22148 41806
rect 24668 41804 24724 41860
rect 25900 41858 25956 41860
rect 25900 41806 25902 41858
rect 25902 41806 25954 41858
rect 25954 41806 25956 41858
rect 25900 41804 25956 41806
rect 28700 41970 28756 41972
rect 28700 41918 28702 41970
rect 28702 41918 28754 41970
rect 28754 41918 28756 41970
rect 28700 41916 28756 41918
rect 31388 41916 31444 41972
rect 28476 41804 28532 41860
rect 29708 41858 29764 41860
rect 29708 41806 29710 41858
rect 29710 41806 29762 41858
rect 29762 41806 29764 41858
rect 29708 41804 29764 41806
rect 25340 40402 25396 40404
rect 25340 40350 25342 40402
rect 25342 40350 25394 40402
rect 25394 40350 25396 40402
rect 25340 40348 25396 40350
rect 28476 40402 28532 40404
rect 28476 40350 28478 40402
rect 28478 40350 28530 40402
rect 28530 40350 28532 40402
rect 28476 40348 28532 40350
rect 24892 40236 24948 40292
rect 21084 39452 21140 39508
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 21868 37884 21924 37940
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 17276 36482 17332 36484
rect 17276 36430 17278 36482
rect 17278 36430 17330 36482
rect 17330 36430 17332 36482
rect 17276 36428 17332 36430
rect 15596 36370 15652 36372
rect 15596 36318 15598 36370
rect 15598 36318 15650 36370
rect 15650 36318 15652 36370
rect 15596 36316 15652 36318
rect 11116 35196 11172 35252
rect 11564 35420 11620 35476
rect 11116 34914 11172 34916
rect 11116 34862 11118 34914
rect 11118 34862 11170 34914
rect 11170 34862 11172 34914
rect 11116 34860 11172 34862
rect 10444 34524 10500 34580
rect 10556 34300 10612 34356
rect 10220 33516 10276 33572
rect 10892 34690 10948 34692
rect 10892 34638 10894 34690
rect 10894 34638 10946 34690
rect 10946 34638 10948 34690
rect 10892 34636 10948 34638
rect 11340 35026 11396 35028
rect 11340 34974 11342 35026
rect 11342 34974 11394 35026
rect 11394 34974 11396 35026
rect 11340 34972 11396 34974
rect 14588 35474 14644 35476
rect 14588 35422 14590 35474
rect 14590 35422 14642 35474
rect 14642 35422 14644 35474
rect 14588 35420 14644 35422
rect 14924 35420 14980 35476
rect 14140 35196 14196 35252
rect 10668 33516 10724 33572
rect 11340 34300 11396 34356
rect 10332 28588 10388 28644
rect 8988 27020 9044 27076
rect 9996 28028 10052 28084
rect 8764 24946 8820 24948
rect 8764 24894 8766 24946
rect 8766 24894 8818 24946
rect 8818 24894 8820 24946
rect 8764 24892 8820 24894
rect 9212 25676 9268 25732
rect 8316 24444 8372 24500
rect 8092 24220 8148 24276
rect 7980 23436 8036 23492
rect 8764 23548 8820 23604
rect 8652 22370 8708 22372
rect 8652 22318 8654 22370
rect 8654 22318 8706 22370
rect 8706 22318 8708 22370
rect 8652 22316 8708 22318
rect 9100 23212 9156 23268
rect 7420 21586 7476 21588
rect 7420 21534 7422 21586
rect 7422 21534 7474 21586
rect 7474 21534 7476 21586
rect 7420 21532 7476 21534
rect 7420 20636 7476 20692
rect 7756 20130 7812 20132
rect 7756 20078 7758 20130
rect 7758 20078 7810 20130
rect 7810 20078 7812 20130
rect 7756 20076 7812 20078
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 6972 18284 7028 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4396 16994 4452 16996
rect 4396 16942 4398 16994
rect 4398 16942 4450 16994
rect 4450 16942 4452 16994
rect 4396 16940 4452 16942
rect 1932 16828 1988 16884
rect 3612 16882 3668 16884
rect 3612 16830 3614 16882
rect 3614 16830 3666 16882
rect 3666 16830 3668 16882
rect 3612 16828 3668 16830
rect 4844 16828 4900 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 2604 16210 2660 16212
rect 2604 16158 2606 16210
rect 2606 16158 2658 16210
rect 2658 16158 2660 16210
rect 2604 16156 2660 16158
rect 6524 16770 6580 16772
rect 6524 16718 6526 16770
rect 6526 16718 6578 16770
rect 6578 16718 6580 16770
rect 6524 16716 6580 16718
rect 5740 16210 5796 16212
rect 5740 16158 5742 16210
rect 5742 16158 5794 16210
rect 5794 16158 5796 16210
rect 5740 16156 5796 16158
rect 6972 16156 7028 16212
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4172 13580 4228 13636
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 6412 12402 6468 12404
rect 6412 12350 6414 12402
rect 6414 12350 6466 12402
rect 6466 12350 6468 12402
rect 6412 12348 6468 12350
rect 4844 12236 4900 12292
rect 1932 11900 1988 11956
rect 3500 11900 3556 11956
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5740 11900 5796 11956
rect 5740 11506 5796 11508
rect 5740 11454 5742 11506
rect 5742 11454 5794 11506
rect 5794 11454 5796 11506
rect 5740 11452 5796 11454
rect 6972 11452 7028 11508
rect 2604 11394 2660 11396
rect 2604 11342 2606 11394
rect 2606 11342 2658 11394
rect 2658 11342 2660 11394
rect 2604 11340 2660 11342
rect 6972 10332 7028 10388
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 8316 21644 8372 21700
rect 8204 18508 8260 18564
rect 9548 25452 9604 25508
rect 9884 27074 9940 27076
rect 9884 27022 9886 27074
rect 9886 27022 9938 27074
rect 9938 27022 9940 27074
rect 9884 27020 9940 27022
rect 9660 25004 9716 25060
rect 9548 23212 9604 23268
rect 9996 23548 10052 23604
rect 10220 24498 10276 24500
rect 10220 24446 10222 24498
rect 10222 24446 10274 24498
rect 10274 24446 10276 24498
rect 10220 24444 10276 24446
rect 12348 34690 12404 34692
rect 12348 34638 12350 34690
rect 12350 34638 12402 34690
rect 12402 34638 12404 34690
rect 12348 34636 12404 34638
rect 14700 34972 14756 35028
rect 16940 36370 16996 36372
rect 16940 36318 16942 36370
rect 16942 36318 16994 36370
rect 16994 36318 16996 36370
rect 16940 36316 16996 36318
rect 16156 36204 16212 36260
rect 15708 35420 15764 35476
rect 15596 35026 15652 35028
rect 15596 34974 15598 35026
rect 15598 34974 15650 35026
rect 15650 34974 15652 35026
rect 15596 34972 15652 34974
rect 15372 34914 15428 34916
rect 15372 34862 15374 34914
rect 15374 34862 15426 34914
rect 15426 34862 15428 34914
rect 15372 34860 15428 34862
rect 14364 34802 14420 34804
rect 14364 34750 14366 34802
rect 14366 34750 14418 34802
rect 14418 34750 14420 34802
rect 14364 34748 14420 34750
rect 11676 34300 11732 34356
rect 14140 34130 14196 34132
rect 14140 34078 14142 34130
rect 14142 34078 14194 34130
rect 14194 34078 14196 34130
rect 14140 34076 14196 34078
rect 14364 33906 14420 33908
rect 14364 33854 14366 33906
rect 14366 33854 14418 33906
rect 14418 33854 14420 33906
rect 14364 33852 14420 33854
rect 11452 33516 11508 33572
rect 11676 33122 11732 33124
rect 11676 33070 11678 33122
rect 11678 33070 11730 33122
rect 11730 33070 11732 33122
rect 11676 33068 11732 33070
rect 12908 33068 12964 33124
rect 12908 31778 12964 31780
rect 12908 31726 12910 31778
rect 12910 31726 12962 31778
rect 12962 31726 12964 31778
rect 12908 31724 12964 31726
rect 13580 31778 13636 31780
rect 13580 31726 13582 31778
rect 13582 31726 13634 31778
rect 13634 31726 13636 31778
rect 13580 31724 13636 31726
rect 13020 31612 13076 31668
rect 10892 30882 10948 30884
rect 10892 30830 10894 30882
rect 10894 30830 10946 30882
rect 10946 30830 10948 30882
rect 10892 30828 10948 30830
rect 14028 31500 14084 31556
rect 11228 29650 11284 29652
rect 11228 29598 11230 29650
rect 11230 29598 11282 29650
rect 11282 29598 11284 29650
rect 11228 29596 11284 29598
rect 11452 29596 11508 29652
rect 10892 27132 10948 27188
rect 11900 29650 11956 29652
rect 11900 29598 11902 29650
rect 11902 29598 11954 29650
rect 11954 29598 11956 29650
rect 11900 29596 11956 29598
rect 14028 29596 14084 29652
rect 14364 30268 14420 30324
rect 11676 28700 11732 28756
rect 12572 28700 12628 28756
rect 11452 28588 11508 28644
rect 11900 28364 11956 28420
rect 12796 28700 12852 28756
rect 12460 28364 12516 28420
rect 11900 27970 11956 27972
rect 11900 27918 11902 27970
rect 11902 27918 11954 27970
rect 11954 27918 11956 27970
rect 11900 27916 11956 27918
rect 11676 27858 11732 27860
rect 11676 27806 11678 27858
rect 11678 27806 11730 27858
rect 11730 27806 11732 27858
rect 11676 27804 11732 27806
rect 10780 26348 10836 26404
rect 10444 25676 10500 25732
rect 10556 26290 10612 26292
rect 10556 26238 10558 26290
rect 10558 26238 10610 26290
rect 10610 26238 10612 26290
rect 10556 26236 10612 26238
rect 10556 25564 10612 25620
rect 10780 25676 10836 25732
rect 10668 25282 10724 25284
rect 10668 25230 10670 25282
rect 10670 25230 10722 25282
rect 10722 25230 10724 25282
rect 10668 25228 10724 25230
rect 10556 25004 10612 25060
rect 10668 24220 10724 24276
rect 9996 22482 10052 22484
rect 9996 22430 9998 22482
rect 9998 22430 10050 22482
rect 10050 22430 10052 22482
rect 9996 22428 10052 22430
rect 9436 20076 9492 20132
rect 9996 20076 10052 20132
rect 10556 19964 10612 20020
rect 8988 17554 9044 17556
rect 8988 17502 8990 17554
rect 8990 17502 9042 17554
rect 9042 17502 9044 17554
rect 8988 17500 9044 17502
rect 9436 18844 9492 18900
rect 8988 16716 9044 16772
rect 9100 16940 9156 16996
rect 8988 16156 9044 16212
rect 9660 18732 9716 18788
rect 10108 19794 10164 19796
rect 10108 19742 10110 19794
rect 10110 19742 10162 19794
rect 10162 19742 10164 19794
rect 10108 19740 10164 19742
rect 11564 26908 11620 26964
rect 11452 26236 11508 26292
rect 11004 25676 11060 25732
rect 11340 25676 11396 25732
rect 11004 25394 11060 25396
rect 11004 25342 11006 25394
rect 11006 25342 11058 25394
rect 11058 25342 11060 25394
rect 11004 25340 11060 25342
rect 11116 25004 11172 25060
rect 12124 27186 12180 27188
rect 12124 27134 12126 27186
rect 12126 27134 12178 27186
rect 12178 27134 12180 27186
rect 12124 27132 12180 27134
rect 12908 28642 12964 28644
rect 12908 28590 12910 28642
rect 12910 28590 12962 28642
rect 12962 28590 12964 28642
rect 12908 28588 12964 28590
rect 12572 27020 12628 27076
rect 12684 26908 12740 26964
rect 12236 26514 12292 26516
rect 12236 26462 12238 26514
rect 12238 26462 12290 26514
rect 12290 26462 12292 26514
rect 12236 26460 12292 26462
rect 13132 26514 13188 26516
rect 13132 26462 13134 26514
rect 13134 26462 13186 26514
rect 13186 26462 13188 26514
rect 13132 26460 13188 26462
rect 11900 26402 11956 26404
rect 11900 26350 11902 26402
rect 11902 26350 11954 26402
rect 11954 26350 11956 26402
rect 11900 26348 11956 26350
rect 12908 25676 12964 25732
rect 14140 27020 14196 27076
rect 13580 26290 13636 26292
rect 13580 26238 13582 26290
rect 13582 26238 13634 26290
rect 13634 26238 13636 26290
rect 13580 26236 13636 26238
rect 13580 25730 13636 25732
rect 13580 25678 13582 25730
rect 13582 25678 13634 25730
rect 13634 25678 13636 25730
rect 13580 25676 13636 25678
rect 14028 25564 14084 25620
rect 13244 24556 13300 24612
rect 15372 34636 15428 34692
rect 15260 33852 15316 33908
rect 15260 32562 15316 32564
rect 15260 32510 15262 32562
rect 15262 32510 15314 32562
rect 15314 32510 15316 32562
rect 15260 32508 15316 32510
rect 15148 31666 15204 31668
rect 15148 31614 15150 31666
rect 15150 31614 15202 31666
rect 15202 31614 15204 31666
rect 15148 31612 15204 31614
rect 14924 30268 14980 30324
rect 15148 28588 15204 28644
rect 15932 35084 15988 35140
rect 19068 36428 19124 36484
rect 17724 36258 17780 36260
rect 17724 36206 17726 36258
rect 17726 36206 17778 36258
rect 17778 36206 17780 36258
rect 17724 36204 17780 36206
rect 17500 36092 17556 36148
rect 18060 36092 18116 36148
rect 16268 35756 16324 35812
rect 16380 35698 16436 35700
rect 16380 35646 16382 35698
rect 16382 35646 16434 35698
rect 16434 35646 16436 35698
rect 16380 35644 16436 35646
rect 17388 35698 17444 35700
rect 17388 35646 17390 35698
rect 17390 35646 17442 35698
rect 17442 35646 17444 35698
rect 17388 35644 17444 35646
rect 16492 35474 16548 35476
rect 16492 35422 16494 35474
rect 16494 35422 16546 35474
rect 16546 35422 16548 35474
rect 16492 35420 16548 35422
rect 17164 35420 17220 35476
rect 16828 34860 16884 34916
rect 18172 35756 18228 35812
rect 17836 35698 17892 35700
rect 17836 35646 17838 35698
rect 17838 35646 17890 35698
rect 17890 35646 17892 35698
rect 17836 35644 17892 35646
rect 18620 35810 18676 35812
rect 18620 35758 18622 35810
rect 18622 35758 18674 35810
rect 18674 35758 18676 35810
rect 18620 35756 18676 35758
rect 18732 35698 18788 35700
rect 18732 35646 18734 35698
rect 18734 35646 18786 35698
rect 18786 35646 18788 35698
rect 18732 35644 18788 35646
rect 19180 35698 19236 35700
rect 19180 35646 19182 35698
rect 19182 35646 19234 35698
rect 19234 35646 19236 35698
rect 19180 35644 19236 35646
rect 17724 35138 17780 35140
rect 17724 35086 17726 35138
rect 17726 35086 17778 35138
rect 17778 35086 17780 35138
rect 17724 35084 17780 35086
rect 18620 35474 18676 35476
rect 18620 35422 18622 35474
rect 18622 35422 18674 35474
rect 18674 35422 18676 35474
rect 18620 35420 18676 35422
rect 17052 33516 17108 33572
rect 16940 32508 16996 32564
rect 15932 30994 15988 30996
rect 15932 30942 15934 30994
rect 15934 30942 15986 30994
rect 15986 30942 15988 30994
rect 15932 30940 15988 30942
rect 16156 30322 16212 30324
rect 16156 30270 16158 30322
rect 16158 30270 16210 30322
rect 16210 30270 16212 30322
rect 16156 30268 16212 30270
rect 15708 30098 15764 30100
rect 15708 30046 15710 30098
rect 15710 30046 15762 30098
rect 15762 30046 15764 30098
rect 15708 30044 15764 30046
rect 15372 27916 15428 27972
rect 15148 27804 15204 27860
rect 14476 26796 14532 26852
rect 15372 27020 15428 27076
rect 14588 25564 14644 25620
rect 14364 25506 14420 25508
rect 14364 25454 14366 25506
rect 14366 25454 14418 25506
rect 14418 25454 14420 25506
rect 14364 25452 14420 25454
rect 14364 23266 14420 23268
rect 14364 23214 14366 23266
rect 14366 23214 14418 23266
rect 14418 23214 14420 23266
rect 14364 23212 14420 23214
rect 11452 21532 11508 21588
rect 11340 20690 11396 20692
rect 11340 20638 11342 20690
rect 11342 20638 11394 20690
rect 11394 20638 11396 20690
rect 11340 20636 11396 20638
rect 10780 20188 10836 20244
rect 10892 19740 10948 19796
rect 9884 18396 9940 18452
rect 10108 18338 10164 18340
rect 10108 18286 10110 18338
rect 10110 18286 10162 18338
rect 10162 18286 10164 18338
rect 10108 18284 10164 18286
rect 10108 17500 10164 17556
rect 9548 16882 9604 16884
rect 9548 16830 9550 16882
rect 9550 16830 9602 16882
rect 9602 16830 9604 16882
rect 9548 16828 9604 16830
rect 9884 16716 9940 16772
rect 8092 13132 8148 13188
rect 7980 12684 8036 12740
rect 8652 13244 8708 13300
rect 9772 16098 9828 16100
rect 9772 16046 9774 16098
rect 9774 16046 9826 16098
rect 9826 16046 9828 16098
rect 9772 16044 9828 16046
rect 9772 15820 9828 15876
rect 10444 18508 10500 18564
rect 10332 17106 10388 17108
rect 10332 17054 10334 17106
rect 10334 17054 10386 17106
rect 10386 17054 10388 17106
rect 10332 17052 10388 17054
rect 10668 17554 10724 17556
rect 10668 17502 10670 17554
rect 10670 17502 10722 17554
rect 10722 17502 10724 17554
rect 10668 17500 10724 17502
rect 10220 16882 10276 16884
rect 10220 16830 10222 16882
rect 10222 16830 10274 16882
rect 10274 16830 10276 16882
rect 10220 16828 10276 16830
rect 10220 16044 10276 16100
rect 8316 12684 8372 12740
rect 7980 12348 8036 12404
rect 9660 13634 9716 13636
rect 9660 13582 9662 13634
rect 9662 13582 9714 13634
rect 9714 13582 9716 13634
rect 9660 13580 9716 13582
rect 9212 13468 9268 13524
rect 9660 13132 9716 13188
rect 10108 13916 10164 13972
rect 9996 13522 10052 13524
rect 9996 13470 9998 13522
rect 9998 13470 10050 13522
rect 10050 13470 10052 13522
rect 9996 13468 10052 13470
rect 9772 13020 9828 13076
rect 9996 13244 10052 13300
rect 8876 12850 8932 12852
rect 8876 12798 8878 12850
rect 8878 12798 8930 12850
rect 8930 12798 8932 12850
rect 8876 12796 8932 12798
rect 9100 12738 9156 12740
rect 9100 12686 9102 12738
rect 9102 12686 9154 12738
rect 9154 12686 9156 12738
rect 9100 12684 9156 12686
rect 9212 12572 9268 12628
rect 9100 12124 9156 12180
rect 10108 12908 10164 12964
rect 10556 13916 10612 13972
rect 10444 13186 10500 13188
rect 10444 13134 10446 13186
rect 10446 13134 10498 13186
rect 10498 13134 10500 13186
rect 10444 13132 10500 13134
rect 10444 12962 10500 12964
rect 10444 12910 10446 12962
rect 10446 12910 10498 12962
rect 10498 12910 10500 12962
rect 10444 12908 10500 12910
rect 9548 12178 9604 12180
rect 9548 12126 9550 12178
rect 9550 12126 9602 12178
rect 9602 12126 9604 12178
rect 9548 12124 9604 12126
rect 9996 11676 10052 11732
rect 8876 11170 8932 11172
rect 8876 11118 8878 11170
rect 8878 11118 8930 11170
rect 8930 11118 8932 11170
rect 8876 11116 8932 11118
rect 10556 12572 10612 12628
rect 11004 16380 11060 16436
rect 11116 16044 11172 16100
rect 12124 21586 12180 21588
rect 12124 21534 12126 21586
rect 12126 21534 12178 21586
rect 12178 21534 12180 21586
rect 12124 21532 12180 21534
rect 11788 21420 11844 21476
rect 13692 21698 13748 21700
rect 13692 21646 13694 21698
rect 13694 21646 13746 21698
rect 13746 21646 13748 21698
rect 13692 21644 13748 21646
rect 12572 20578 12628 20580
rect 12572 20526 12574 20578
rect 12574 20526 12626 20578
rect 12626 20526 12628 20578
rect 12572 20524 12628 20526
rect 12684 20412 12740 20468
rect 12236 20188 12292 20244
rect 11900 19010 11956 19012
rect 11900 18958 11902 19010
rect 11902 18958 11954 19010
rect 11954 18958 11956 19010
rect 11900 18956 11956 18958
rect 12124 18844 12180 18900
rect 12348 20076 12404 20132
rect 12908 20018 12964 20020
rect 12908 19966 12910 20018
rect 12910 19966 12962 20018
rect 12962 19966 12964 20018
rect 12908 19964 12964 19966
rect 14588 23212 14644 23268
rect 14252 20412 14308 20468
rect 15148 25452 15204 25508
rect 15932 28476 15988 28532
rect 16828 30828 16884 30884
rect 16716 28642 16772 28644
rect 16716 28590 16718 28642
rect 16718 28590 16770 28642
rect 16770 28590 16772 28642
rect 16716 28588 16772 28590
rect 16492 27916 16548 27972
rect 16604 27804 16660 27860
rect 15708 26236 15764 26292
rect 16604 26236 16660 26292
rect 15708 25394 15764 25396
rect 15708 25342 15710 25394
rect 15710 25342 15762 25394
rect 15762 25342 15764 25394
rect 15708 25340 15764 25342
rect 15260 23266 15316 23268
rect 15260 23214 15262 23266
rect 15262 23214 15314 23266
rect 15314 23214 15316 23266
rect 15260 23212 15316 23214
rect 16604 24722 16660 24724
rect 16604 24670 16606 24722
rect 16606 24670 16658 24722
rect 16658 24670 16660 24722
rect 16604 24668 16660 24670
rect 16828 23772 16884 23828
rect 16828 23548 16884 23604
rect 16268 22876 16324 22932
rect 16492 22482 16548 22484
rect 16492 22430 16494 22482
rect 16494 22430 16546 22482
rect 16546 22430 16548 22482
rect 16492 22428 16548 22430
rect 17836 33404 17892 33460
rect 24892 37938 24948 37940
rect 24892 37886 24894 37938
rect 24894 37886 24946 37938
rect 24946 37886 24948 37938
rect 24892 37884 24948 37886
rect 24332 37324 24388 37380
rect 22988 37212 23044 37268
rect 24220 37212 24276 37268
rect 20524 36428 20580 36484
rect 19628 36092 19684 36148
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20076 35756 20132 35812
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 18956 31612 19012 31668
rect 17948 30994 18004 30996
rect 17948 30942 17950 30994
rect 17950 30942 18002 30994
rect 18002 30942 18004 30994
rect 17948 30940 18004 30942
rect 17500 30882 17556 30884
rect 17500 30830 17502 30882
rect 17502 30830 17554 30882
rect 17554 30830 17556 30882
rect 17500 30828 17556 30830
rect 17276 28642 17332 28644
rect 17276 28590 17278 28642
rect 17278 28590 17330 28642
rect 17330 28590 17332 28642
rect 17276 28588 17332 28590
rect 17388 28530 17444 28532
rect 17388 28478 17390 28530
rect 17390 28478 17442 28530
rect 17442 28478 17444 28530
rect 17388 28476 17444 28478
rect 17164 27916 17220 27972
rect 17164 27692 17220 27748
rect 17164 27074 17220 27076
rect 17164 27022 17166 27074
rect 17166 27022 17218 27074
rect 17218 27022 17220 27074
rect 17164 27020 17220 27022
rect 17388 26290 17444 26292
rect 17388 26238 17390 26290
rect 17390 26238 17442 26290
rect 17442 26238 17444 26290
rect 17388 26236 17444 26238
rect 18956 30268 19012 30324
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20748 31554 20804 31556
rect 20748 31502 20750 31554
rect 20750 31502 20802 31554
rect 20802 31502 20804 31554
rect 20748 31500 20804 31502
rect 25788 37772 25844 37828
rect 25564 37378 25620 37380
rect 25564 37326 25566 37378
rect 25566 37326 25618 37378
rect 25618 37326 25620 37378
rect 25564 37324 25620 37326
rect 25228 37266 25284 37268
rect 25228 37214 25230 37266
rect 25230 37214 25282 37266
rect 25282 37214 25284 37266
rect 25228 37212 25284 37214
rect 24556 36988 24612 37044
rect 24220 36428 24276 36484
rect 25564 36428 25620 36484
rect 23660 35644 23716 35700
rect 25676 36204 25732 36260
rect 25788 34802 25844 34804
rect 25788 34750 25790 34802
rect 25790 34750 25842 34802
rect 25842 34750 25844 34802
rect 25788 34748 25844 34750
rect 23772 34636 23828 34692
rect 23100 33458 23156 33460
rect 23100 33406 23102 33458
rect 23102 33406 23154 33458
rect 23154 33406 23156 33458
rect 23100 33404 23156 33406
rect 25676 34690 25732 34692
rect 25676 34638 25678 34690
rect 25678 34638 25730 34690
rect 25730 34638 25732 34690
rect 25676 34636 25732 34638
rect 28364 40124 28420 40180
rect 28252 39394 28308 39396
rect 28252 39342 28254 39394
rect 28254 39342 28306 39394
rect 28306 39342 28308 39394
rect 28252 39340 28308 39342
rect 26348 37826 26404 37828
rect 26348 37774 26350 37826
rect 26350 37774 26402 37826
rect 26402 37774 26404 37826
rect 26348 37772 26404 37774
rect 26012 34690 26068 34692
rect 26012 34638 26014 34690
rect 26014 34638 26066 34690
rect 26066 34638 26068 34690
rect 26012 34636 26068 34638
rect 23884 33180 23940 33236
rect 22876 32508 22932 32564
rect 24668 33234 24724 33236
rect 24668 33182 24670 33234
rect 24670 33182 24722 33234
rect 24722 33182 24724 33234
rect 24668 33180 24724 33182
rect 25116 32732 25172 32788
rect 23884 32562 23940 32564
rect 23884 32510 23886 32562
rect 23886 32510 23938 32562
rect 23938 32510 23940 32562
rect 23884 32508 23940 32510
rect 24108 32562 24164 32564
rect 24108 32510 24110 32562
rect 24110 32510 24162 32562
rect 24162 32510 24164 32562
rect 24108 32508 24164 32510
rect 25564 31836 25620 31892
rect 27580 37324 27636 37380
rect 26796 36316 26852 36372
rect 26572 36204 26628 36260
rect 26908 36204 26964 36260
rect 27468 36204 27524 36260
rect 27356 34748 27412 34804
rect 27132 34188 27188 34244
rect 26348 34130 26404 34132
rect 26348 34078 26350 34130
rect 26350 34078 26402 34130
rect 26402 34078 26404 34130
rect 26348 34076 26404 34078
rect 26908 34076 26964 34132
rect 26796 33122 26852 33124
rect 26796 33070 26798 33122
rect 26798 33070 26850 33122
rect 26850 33070 26852 33122
rect 26796 33068 26852 33070
rect 26684 32508 26740 32564
rect 26572 32396 26628 32452
rect 27244 34076 27300 34132
rect 27468 34130 27524 34132
rect 27468 34078 27470 34130
rect 27470 34078 27522 34130
rect 27522 34078 27524 34130
rect 27468 34076 27524 34078
rect 32508 41970 32564 41972
rect 32508 41918 32510 41970
rect 32510 41918 32562 41970
rect 32562 41918 32564 41970
rect 32508 41916 32564 41918
rect 36092 41804 36148 41860
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 32620 40626 32676 40628
rect 32620 40574 32622 40626
rect 32622 40574 32674 40626
rect 32674 40574 32676 40626
rect 32620 40572 32676 40574
rect 34188 40572 34244 40628
rect 31500 40236 31556 40292
rect 29260 39340 29316 39396
rect 28476 37324 28532 37380
rect 30268 37324 30324 37380
rect 29484 36482 29540 36484
rect 29484 36430 29486 36482
rect 29486 36430 29538 36482
rect 29538 36430 29540 36482
rect 29484 36428 29540 36430
rect 27692 34636 27748 34692
rect 27916 34242 27972 34244
rect 27916 34190 27918 34242
rect 27918 34190 27970 34242
rect 27970 34190 27972 34242
rect 27916 34188 27972 34190
rect 28028 34130 28084 34132
rect 28028 34078 28030 34130
rect 28030 34078 28082 34130
rect 28082 34078 28084 34130
rect 28028 34076 28084 34078
rect 27468 33122 27524 33124
rect 27468 33070 27470 33122
rect 27470 33070 27522 33122
rect 27522 33070 27524 33122
rect 27468 33068 27524 33070
rect 27132 32956 27188 33012
rect 27020 32450 27076 32452
rect 27020 32398 27022 32450
rect 27022 32398 27074 32450
rect 27074 32398 27076 32450
rect 27020 32396 27076 32398
rect 27020 32060 27076 32116
rect 26684 31778 26740 31780
rect 26684 31726 26686 31778
rect 26686 31726 26738 31778
rect 26738 31726 26740 31778
rect 26684 31724 26740 31726
rect 21644 31554 21700 31556
rect 21644 31502 21646 31554
rect 21646 31502 21698 31554
rect 21698 31502 21700 31554
rect 21644 31500 21700 31502
rect 20188 30882 20244 30884
rect 20188 30830 20190 30882
rect 20190 30830 20242 30882
rect 20242 30830 20244 30882
rect 20188 30828 20244 30830
rect 19628 30268 19684 30324
rect 24108 31500 24164 31556
rect 23436 31388 23492 31444
rect 21644 30268 21700 30324
rect 22540 30268 22596 30324
rect 18284 30098 18340 30100
rect 18284 30046 18286 30098
rect 18286 30046 18338 30098
rect 18338 30046 18340 30098
rect 18284 30044 18340 30046
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20300 28700 20356 28756
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19740 27746 19796 27748
rect 19740 27694 19742 27746
rect 19742 27694 19794 27746
rect 19794 27694 19796 27746
rect 19740 27692 19796 27694
rect 17724 27132 17780 27188
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 18732 26514 18788 26516
rect 18732 26462 18734 26514
rect 18734 26462 18786 26514
rect 18786 26462 18788 26514
rect 18732 26460 18788 26462
rect 17724 24892 17780 24948
rect 18060 25004 18116 25060
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 17500 24780 17556 24836
rect 17388 24722 17444 24724
rect 17388 24670 17390 24722
rect 17390 24670 17442 24722
rect 17442 24670 17444 24722
rect 17388 24668 17444 24670
rect 17948 24220 18004 24276
rect 19516 24220 19572 24276
rect 17724 23548 17780 23604
rect 18284 23938 18340 23940
rect 18284 23886 18286 23938
rect 18286 23886 18338 23938
rect 18338 23886 18340 23938
rect 18284 23884 18340 23886
rect 18284 23548 18340 23604
rect 18732 23826 18788 23828
rect 18732 23774 18734 23826
rect 18734 23774 18786 23826
rect 18786 23774 18788 23826
rect 18732 23772 18788 23774
rect 15372 21308 15428 21364
rect 15260 20636 15316 20692
rect 14588 20412 14644 20468
rect 13804 18732 13860 18788
rect 11452 17500 11508 17556
rect 11340 17052 11396 17108
rect 11900 16994 11956 16996
rect 11900 16942 11902 16994
rect 11902 16942 11954 16994
rect 11954 16942 11956 16994
rect 11900 16940 11956 16942
rect 11452 16658 11508 16660
rect 11452 16606 11454 16658
rect 11454 16606 11506 16658
rect 11506 16606 11508 16658
rect 11452 16604 11508 16606
rect 11676 16044 11732 16100
rect 12348 16604 12404 16660
rect 12124 16156 12180 16212
rect 12460 16098 12516 16100
rect 12460 16046 12462 16098
rect 12462 16046 12514 16098
rect 12514 16046 12516 16098
rect 12460 16044 12516 16046
rect 12236 15986 12292 15988
rect 12236 15934 12238 15986
rect 12238 15934 12290 15986
rect 12290 15934 12292 15986
rect 12236 15932 12292 15934
rect 12796 15932 12852 15988
rect 16268 21362 16324 21364
rect 16268 21310 16270 21362
rect 16270 21310 16322 21362
rect 16322 21310 16324 21362
rect 16268 21308 16324 21310
rect 16604 20748 16660 20804
rect 15708 18508 15764 18564
rect 14700 18396 14756 18452
rect 15372 18450 15428 18452
rect 15372 18398 15374 18450
rect 15374 18398 15426 18450
rect 15426 18398 15428 18450
rect 15372 18396 15428 18398
rect 14140 18172 14196 18228
rect 13356 16882 13412 16884
rect 13356 16830 13358 16882
rect 13358 16830 13410 16882
rect 13410 16830 13412 16882
rect 13356 16828 13412 16830
rect 13804 16994 13860 16996
rect 13804 16942 13806 16994
rect 13806 16942 13858 16994
rect 13858 16942 13860 16994
rect 13804 16940 13860 16942
rect 14028 16828 14084 16884
rect 16268 18956 16324 19012
rect 16156 18562 16212 18564
rect 16156 18510 16158 18562
rect 16158 18510 16210 18562
rect 16210 18510 16212 18562
rect 16156 18508 16212 18510
rect 16156 18284 16212 18340
rect 16156 16882 16212 16884
rect 16156 16830 16158 16882
rect 16158 16830 16210 16882
rect 16210 16830 16212 16882
rect 16156 16828 16212 16830
rect 13132 16716 13188 16772
rect 13020 16156 13076 16212
rect 13132 16044 13188 16100
rect 14588 15820 14644 15876
rect 11340 13916 11396 13972
rect 11116 13132 11172 13188
rect 11452 12850 11508 12852
rect 11452 12798 11454 12850
rect 11454 12798 11506 12850
rect 11506 12798 11508 12850
rect 11452 12796 11508 12798
rect 11116 12738 11172 12740
rect 11116 12686 11118 12738
rect 11118 12686 11170 12738
rect 11170 12686 11172 12738
rect 11116 12684 11172 12686
rect 10780 12236 10836 12292
rect 11116 12290 11172 12292
rect 11116 12238 11118 12290
rect 11118 12238 11170 12290
rect 11170 12238 11172 12290
rect 11116 12236 11172 12238
rect 11228 11676 11284 11732
rect 10220 11340 10276 11396
rect 9996 11116 10052 11172
rect 7868 10610 7924 10612
rect 7868 10558 7870 10610
rect 7870 10558 7922 10610
rect 7922 10558 7924 10610
rect 7868 10556 7924 10558
rect 8204 10610 8260 10612
rect 8204 10558 8206 10610
rect 8206 10558 8258 10610
rect 8258 10558 8260 10610
rect 8204 10556 8260 10558
rect 8876 10498 8932 10500
rect 8876 10446 8878 10498
rect 8878 10446 8930 10498
rect 8930 10446 8932 10498
rect 8876 10444 8932 10446
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 5628 8370 5684 8372
rect 5628 8318 5630 8370
rect 5630 8318 5682 8370
rect 5682 8318 5684 8370
rect 5628 8316 5684 8318
rect 8764 10332 8820 10388
rect 7532 8316 7588 8372
rect 7756 9548 7812 9604
rect 8540 9602 8596 9604
rect 8540 9550 8542 9602
rect 8542 9550 8594 9602
rect 8594 9550 8596 9602
rect 8540 9548 8596 9550
rect 11788 11170 11844 11172
rect 11788 11118 11790 11170
rect 11790 11118 11842 11170
rect 11842 11118 11844 11170
rect 11788 11116 11844 11118
rect 10220 10780 10276 10836
rect 10668 10834 10724 10836
rect 10668 10782 10670 10834
rect 10670 10782 10722 10834
rect 10722 10782 10724 10834
rect 10668 10780 10724 10782
rect 9772 9436 9828 9492
rect 12124 11282 12180 11284
rect 12124 11230 12126 11282
rect 12126 11230 12178 11282
rect 12178 11230 12180 11282
rect 12124 11228 12180 11230
rect 12684 11228 12740 11284
rect 12684 10668 12740 10724
rect 12460 9826 12516 9828
rect 12460 9774 12462 9826
rect 12462 9774 12514 9826
rect 12514 9774 12516 9826
rect 12460 9772 12516 9774
rect 12348 9266 12404 9268
rect 12348 9214 12350 9266
rect 12350 9214 12402 9266
rect 12402 9214 12404 9266
rect 12348 9212 12404 9214
rect 9660 7532 9716 7588
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 12908 11116 12964 11172
rect 15260 15148 15316 15204
rect 14924 14530 14980 14532
rect 14924 14478 14926 14530
rect 14926 14478 14978 14530
rect 14978 14478 14980 14530
rect 14924 14476 14980 14478
rect 15484 14530 15540 14532
rect 15484 14478 15486 14530
rect 15486 14478 15538 14530
rect 15538 14478 15540 14530
rect 15484 14476 15540 14478
rect 14812 13970 14868 13972
rect 14812 13918 14814 13970
rect 14814 13918 14866 13970
rect 14866 13918 14868 13970
rect 14812 13916 14868 13918
rect 13580 10722 13636 10724
rect 13580 10670 13582 10722
rect 13582 10670 13634 10722
rect 13634 10670 13636 10722
rect 13580 10668 13636 10670
rect 13916 10668 13972 10724
rect 12908 10556 12964 10612
rect 12908 10332 12964 10388
rect 14364 10444 14420 10500
rect 13692 10332 13748 10388
rect 12796 9436 12852 9492
rect 12908 9212 12964 9268
rect 13580 9772 13636 9828
rect 13916 9772 13972 9828
rect 15596 13970 15652 13972
rect 15596 13918 15598 13970
rect 15598 13918 15650 13970
rect 15650 13918 15652 13970
rect 15596 13916 15652 13918
rect 15260 10498 15316 10500
rect 15260 10446 15262 10498
rect 15262 10446 15314 10498
rect 15314 10446 15316 10498
rect 15260 10444 15316 10446
rect 13580 9100 13636 9156
rect 15036 9826 15092 9828
rect 15036 9774 15038 9826
rect 15038 9774 15090 9826
rect 15090 9774 15092 9826
rect 15036 9772 15092 9774
rect 15484 9826 15540 9828
rect 15484 9774 15486 9826
rect 15486 9774 15538 9826
rect 15538 9774 15540 9826
rect 15484 9772 15540 9774
rect 15372 9660 15428 9716
rect 14812 9602 14868 9604
rect 14812 9550 14814 9602
rect 14814 9550 14866 9602
rect 14866 9550 14868 9602
rect 14812 9548 14868 9550
rect 14700 9100 14756 9156
rect 15148 9324 15204 9380
rect 15708 9772 15764 9828
rect 16156 15484 16212 15540
rect 15932 14530 15988 14532
rect 15932 14478 15934 14530
rect 15934 14478 15986 14530
rect 15986 14478 15988 14530
rect 15932 14476 15988 14478
rect 16716 20636 16772 20692
rect 16716 20412 16772 20468
rect 16492 18172 16548 18228
rect 16940 16940 16996 16996
rect 16604 15372 16660 15428
rect 16268 14754 16324 14756
rect 16268 14702 16270 14754
rect 16270 14702 16322 14754
rect 16322 14702 16324 14754
rect 16268 14700 16324 14702
rect 16492 14642 16548 14644
rect 16492 14590 16494 14642
rect 16494 14590 16546 14642
rect 16546 14590 16548 14642
rect 16492 14588 16548 14590
rect 16716 14700 16772 14756
rect 18620 22876 18676 22932
rect 18508 22428 18564 22484
rect 17388 20802 17444 20804
rect 17388 20750 17390 20802
rect 17390 20750 17442 20802
rect 17442 20750 17444 20802
rect 17388 20748 17444 20750
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20188 22988 20244 23044
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 20524 20132 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 17276 19122 17332 19124
rect 17276 19070 17278 19122
rect 17278 19070 17330 19122
rect 17330 19070 17332 19122
rect 17276 19068 17332 19070
rect 17276 18396 17332 18452
rect 17724 17500 17780 17556
rect 17388 16994 17444 16996
rect 17388 16942 17390 16994
rect 17390 16942 17442 16994
rect 17442 16942 17444 16994
rect 17388 16940 17444 16942
rect 17612 16940 17668 16996
rect 17276 16156 17332 16212
rect 17388 15426 17444 15428
rect 17388 15374 17390 15426
rect 17390 15374 17442 15426
rect 17442 15374 17444 15426
rect 17388 15372 17444 15374
rect 17164 14476 17220 14532
rect 16940 13916 16996 13972
rect 16268 10834 16324 10836
rect 16268 10782 16270 10834
rect 16270 10782 16322 10834
rect 16322 10782 16324 10834
rect 16268 10780 16324 10782
rect 15596 9660 15652 9716
rect 15820 9436 15876 9492
rect 15708 9324 15764 9380
rect 15596 9212 15652 9268
rect 15708 8988 15764 9044
rect 15708 8818 15764 8820
rect 15708 8766 15710 8818
rect 15710 8766 15762 8818
rect 15762 8766 15764 8818
rect 15708 8764 15764 8766
rect 12572 7532 12628 7588
rect 12572 6412 12628 6468
rect 13580 6466 13636 6468
rect 13580 6414 13582 6466
rect 13582 6414 13634 6466
rect 13634 6414 13636 6466
rect 13580 6412 13636 6414
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 13580 5068 13636 5124
rect 16492 9548 16548 9604
rect 17164 12684 17220 12740
rect 17948 16940 18004 16996
rect 17836 16828 17892 16884
rect 18060 15484 18116 15540
rect 17612 15148 17668 15204
rect 17724 15260 17780 15316
rect 17612 14588 17668 14644
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 18732 18338 18788 18340
rect 18732 18286 18734 18338
rect 18734 18286 18786 18338
rect 18786 18286 18788 18338
rect 18732 18284 18788 18286
rect 19516 18284 19572 18340
rect 21308 28700 21364 28756
rect 21980 28700 22036 28756
rect 21532 28642 21588 28644
rect 21532 28590 21534 28642
rect 21534 28590 21586 28642
rect 21586 28590 21588 28642
rect 21532 28588 21588 28590
rect 22316 28642 22372 28644
rect 22316 28590 22318 28642
rect 22318 28590 22370 28642
rect 22370 28590 22372 28642
rect 22316 28588 22372 28590
rect 21644 26460 21700 26516
rect 20860 24892 20916 24948
rect 20860 24332 20916 24388
rect 21420 25394 21476 25396
rect 21420 25342 21422 25394
rect 21422 25342 21474 25394
rect 21474 25342 21476 25394
rect 21420 25340 21476 25342
rect 22988 28700 23044 28756
rect 22652 28028 22708 28084
rect 25564 31554 25620 31556
rect 25564 31502 25566 31554
rect 25566 31502 25618 31554
rect 25618 31502 25620 31554
rect 25564 31500 25620 31502
rect 23100 28588 23156 28644
rect 23212 28924 23268 28980
rect 22652 26796 22708 26852
rect 23996 28700 24052 28756
rect 26012 28812 26068 28868
rect 23660 28082 23716 28084
rect 23660 28030 23662 28082
rect 23662 28030 23714 28082
rect 23714 28030 23716 28082
rect 23660 28028 23716 28030
rect 25340 28028 25396 28084
rect 23100 26460 23156 26516
rect 23884 26796 23940 26852
rect 23100 25452 23156 25508
rect 23772 25506 23828 25508
rect 23772 25454 23774 25506
rect 23774 25454 23826 25506
rect 23826 25454 23828 25506
rect 23772 25452 23828 25454
rect 26460 31666 26516 31668
rect 26460 31614 26462 31666
rect 26462 31614 26514 31666
rect 26514 31614 26516 31666
rect 26460 31612 26516 31614
rect 26236 28924 26292 28980
rect 27132 31612 27188 31668
rect 26124 26796 26180 26852
rect 26012 25788 26068 25844
rect 25228 25618 25284 25620
rect 25228 25566 25230 25618
rect 25230 25566 25282 25618
rect 25282 25566 25284 25618
rect 25228 25564 25284 25566
rect 24220 25506 24276 25508
rect 24220 25454 24222 25506
rect 24222 25454 24274 25506
rect 24274 25454 24276 25506
rect 24220 25452 24276 25454
rect 22316 24668 22372 24724
rect 22092 24556 22148 24612
rect 21532 24332 21588 24388
rect 21196 23996 21252 24052
rect 21532 23938 21588 23940
rect 21532 23886 21534 23938
rect 21534 23886 21586 23938
rect 21586 23886 21588 23938
rect 21532 23884 21588 23886
rect 21868 23826 21924 23828
rect 21868 23774 21870 23826
rect 21870 23774 21922 23826
rect 21922 23774 21924 23826
rect 21868 23772 21924 23774
rect 21196 23042 21252 23044
rect 21196 22990 21198 23042
rect 21198 22990 21250 23042
rect 21250 22990 21252 23042
rect 21196 22988 21252 22990
rect 21532 22092 21588 22148
rect 21644 18450 21700 18452
rect 21644 18398 21646 18450
rect 21646 18398 21698 18450
rect 21698 18398 21700 18450
rect 21644 18396 21700 18398
rect 20860 18338 20916 18340
rect 20860 18286 20862 18338
rect 20862 18286 20914 18338
rect 20914 18286 20916 18338
rect 20860 18284 20916 18286
rect 22428 24556 22484 24612
rect 22540 23938 22596 23940
rect 22540 23886 22542 23938
rect 22542 23886 22594 23938
rect 22594 23886 22596 23938
rect 22540 23884 22596 23886
rect 22652 23826 22708 23828
rect 22652 23774 22654 23826
rect 22654 23774 22706 23826
rect 22706 23774 22708 23826
rect 22652 23772 22708 23774
rect 23884 25340 23940 25396
rect 23436 25282 23492 25284
rect 23436 25230 23438 25282
rect 23438 25230 23490 25282
rect 23490 25230 23492 25282
rect 23436 25228 23492 25230
rect 24892 25228 24948 25284
rect 25564 25228 25620 25284
rect 24444 24892 24500 24948
rect 25340 24946 25396 24948
rect 25340 24894 25342 24946
rect 25342 24894 25394 24946
rect 25394 24894 25396 24946
rect 25340 24892 25396 24894
rect 23996 24610 24052 24612
rect 23996 24558 23998 24610
rect 23998 24558 24050 24610
rect 24050 24558 24052 24610
rect 23996 24556 24052 24558
rect 24668 24444 24724 24500
rect 25452 23938 25508 23940
rect 25452 23886 25454 23938
rect 25454 23886 25506 23938
rect 25506 23886 25508 23938
rect 25452 23884 25508 23886
rect 23100 20188 23156 20244
rect 21868 18172 21924 18228
rect 19404 17554 19460 17556
rect 19404 17502 19406 17554
rect 19406 17502 19458 17554
rect 19458 17502 19460 17554
rect 19404 17500 19460 17502
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20300 16828 20356 16884
rect 19292 16210 19348 16212
rect 19292 16158 19294 16210
rect 19294 16158 19346 16210
rect 19346 16158 19348 16210
rect 19292 16156 19348 16158
rect 19292 15820 19348 15876
rect 20860 15932 20916 15988
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19516 15538 19572 15540
rect 19516 15486 19518 15538
rect 19518 15486 19570 15538
rect 19570 15486 19572 15538
rect 19516 15484 19572 15486
rect 18844 15426 18900 15428
rect 18844 15374 18846 15426
rect 18846 15374 18898 15426
rect 18898 15374 18900 15426
rect 18844 15372 18900 15374
rect 19964 15426 20020 15428
rect 19964 15374 19966 15426
rect 19966 15374 20018 15426
rect 20018 15374 20020 15426
rect 19964 15372 20020 15374
rect 18620 15314 18676 15316
rect 18620 15262 18622 15314
rect 18622 15262 18674 15314
rect 18674 15262 18676 15314
rect 18620 15260 18676 15262
rect 18060 15148 18116 15204
rect 20412 15202 20468 15204
rect 20412 15150 20414 15202
rect 20414 15150 20466 15202
rect 20466 15150 20468 15202
rect 20412 15148 20468 15150
rect 18060 14642 18116 14644
rect 18060 14590 18062 14642
rect 18062 14590 18114 14642
rect 18114 14590 18116 14642
rect 18060 14588 18116 14590
rect 18172 14530 18228 14532
rect 18172 14478 18174 14530
rect 18174 14478 18226 14530
rect 18226 14478 18228 14530
rect 18172 14476 18228 14478
rect 19292 15036 19348 15092
rect 18844 14476 18900 14532
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 21084 15372 21140 15428
rect 21532 15372 21588 15428
rect 21868 15426 21924 15428
rect 21868 15374 21870 15426
rect 21870 15374 21922 15426
rect 21922 15374 21924 15426
rect 21868 15372 21924 15374
rect 21868 15148 21924 15204
rect 21420 12908 21476 12964
rect 21756 12796 21812 12852
rect 22876 19794 22932 19796
rect 22876 19742 22878 19794
rect 22878 19742 22930 19794
rect 22930 19742 22932 19794
rect 22876 19740 22932 19742
rect 23548 20188 23604 20244
rect 22092 18450 22148 18452
rect 22092 18398 22094 18450
rect 22094 18398 22146 18450
rect 22146 18398 22148 18450
rect 22092 18396 22148 18398
rect 22988 18396 23044 18452
rect 23660 19740 23716 19796
rect 24220 16716 24276 16772
rect 26236 24946 26292 24948
rect 26236 24894 26238 24946
rect 26238 24894 26290 24946
rect 26290 24894 26292 24946
rect 26236 24892 26292 24894
rect 25900 24722 25956 24724
rect 25900 24670 25902 24722
rect 25902 24670 25954 24722
rect 25954 24670 25956 24722
rect 25900 24668 25956 24670
rect 27132 24946 27188 24948
rect 27132 24894 27134 24946
rect 27134 24894 27186 24946
rect 27186 24894 27188 24946
rect 27132 24892 27188 24894
rect 26684 24780 26740 24836
rect 27580 31890 27636 31892
rect 27580 31838 27582 31890
rect 27582 31838 27634 31890
rect 27634 31838 27636 31890
rect 27580 31836 27636 31838
rect 29148 36370 29204 36372
rect 29148 36318 29150 36370
rect 29150 36318 29202 36370
rect 29202 36318 29204 36370
rect 29148 36316 29204 36318
rect 28364 36258 28420 36260
rect 28364 36206 28366 36258
rect 28366 36206 28418 36258
rect 28418 36206 28420 36258
rect 28364 36204 28420 36206
rect 30828 37378 30884 37380
rect 30828 37326 30830 37378
rect 30830 37326 30882 37378
rect 30882 37326 30884 37378
rect 30828 37324 30884 37326
rect 33404 40402 33460 40404
rect 33404 40350 33406 40402
rect 33406 40350 33458 40402
rect 33458 40350 33460 40402
rect 33404 40348 33460 40350
rect 34972 40236 35028 40292
rect 37324 41858 37380 41860
rect 37324 41806 37326 41858
rect 37326 41806 37378 41858
rect 37378 41806 37380 41858
rect 37324 41804 37380 41806
rect 39900 41804 39956 41860
rect 41132 41858 41188 41860
rect 41132 41806 41134 41858
rect 41134 41806 41186 41858
rect 41186 41806 41188 41858
rect 41132 41804 41188 41806
rect 36876 40236 36932 40292
rect 37996 40236 38052 40292
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34412 39730 34468 39732
rect 34412 39678 34414 39730
rect 34414 39678 34466 39730
rect 34466 39678 34468 39730
rect 34412 39676 34468 39678
rect 31724 37324 31780 37380
rect 30380 36540 30436 36596
rect 30828 36482 30884 36484
rect 30828 36430 30830 36482
rect 30830 36430 30882 36482
rect 30882 36430 30884 36482
rect 30828 36428 30884 36430
rect 30380 35756 30436 35812
rect 30268 34914 30324 34916
rect 30268 34862 30270 34914
rect 30270 34862 30322 34914
rect 30322 34862 30324 34914
rect 30268 34860 30324 34862
rect 31276 34300 31332 34356
rect 31612 34188 31668 34244
rect 28364 32956 28420 33012
rect 32060 34300 32116 34356
rect 31836 34242 31892 34244
rect 31836 34190 31838 34242
rect 31838 34190 31890 34242
rect 31890 34190 31892 34242
rect 31836 34188 31892 34190
rect 33068 34300 33124 34356
rect 33516 34914 33572 34916
rect 33516 34862 33518 34914
rect 33518 34862 33570 34914
rect 33570 34862 33572 34914
rect 33516 34860 33572 34862
rect 31612 33234 31668 33236
rect 31612 33182 31614 33234
rect 31614 33182 31666 33234
rect 31666 33182 31668 33234
rect 31612 33180 31668 33182
rect 31052 32786 31108 32788
rect 31052 32734 31054 32786
rect 31054 32734 31106 32786
rect 31106 32734 31108 32786
rect 31052 32732 31108 32734
rect 30268 32508 30324 32564
rect 28252 31836 28308 31892
rect 30044 32396 30100 32452
rect 30044 31500 30100 31556
rect 30828 31948 30884 32004
rect 30156 30940 30212 30996
rect 30716 31554 30772 31556
rect 30716 31502 30718 31554
rect 30718 31502 30770 31554
rect 30770 31502 30772 31554
rect 30716 31500 30772 31502
rect 30716 31106 30772 31108
rect 30716 31054 30718 31106
rect 30718 31054 30770 31106
rect 30770 31054 30772 31106
rect 30716 31052 30772 31054
rect 28588 30828 28644 30884
rect 28588 30268 28644 30324
rect 30156 30268 30212 30324
rect 29708 30156 29764 30212
rect 28812 30044 28868 30100
rect 28588 28082 28644 28084
rect 28588 28030 28590 28082
rect 28590 28030 28642 28082
rect 28642 28030 28644 28082
rect 28588 28028 28644 28030
rect 28588 27804 28644 27860
rect 28140 27746 28196 27748
rect 28140 27694 28142 27746
rect 28142 27694 28194 27746
rect 28194 27694 28196 27746
rect 28140 27692 28196 27694
rect 29484 29314 29540 29316
rect 29484 29262 29486 29314
rect 29486 29262 29538 29314
rect 29538 29262 29540 29314
rect 29484 29260 29540 29262
rect 30604 30156 30660 30212
rect 30380 29260 30436 29316
rect 29820 28866 29876 28868
rect 29820 28814 29822 28866
rect 29822 28814 29874 28866
rect 29874 28814 29876 28866
rect 29820 28812 29876 28814
rect 29932 28588 29988 28644
rect 28812 28028 28868 28084
rect 28924 27804 28980 27860
rect 27580 24610 27636 24612
rect 27580 24558 27582 24610
rect 27582 24558 27634 24610
rect 27634 24558 27636 24610
rect 27580 24556 27636 24558
rect 26796 22258 26852 22260
rect 26796 22206 26798 22258
rect 26798 22206 26850 22258
rect 26850 22206 26852 22258
rect 26796 22204 26852 22206
rect 28924 25564 28980 25620
rect 31612 32508 31668 32564
rect 32956 33346 33012 33348
rect 32956 33294 32958 33346
rect 32958 33294 33010 33346
rect 33010 33294 33012 33346
rect 32956 33292 33012 33294
rect 32396 33068 32452 33124
rect 32284 32562 32340 32564
rect 32284 32510 32286 32562
rect 32286 32510 32338 32562
rect 32338 32510 32340 32562
rect 32284 32508 32340 32510
rect 31500 31106 31556 31108
rect 31500 31054 31502 31106
rect 31502 31054 31554 31106
rect 31554 31054 31556 31106
rect 31500 31052 31556 31054
rect 32508 30994 32564 30996
rect 32508 30942 32510 30994
rect 32510 30942 32562 30994
rect 32562 30942 32564 30994
rect 32508 30940 32564 30942
rect 32060 30044 32116 30100
rect 31948 28924 32004 28980
rect 31948 28364 32004 28420
rect 30156 27858 30212 27860
rect 30156 27806 30158 27858
rect 30158 27806 30210 27858
rect 30210 27806 30212 27858
rect 30156 27804 30212 27806
rect 29372 27692 29428 27748
rect 29372 26908 29428 26964
rect 30828 27074 30884 27076
rect 30828 27022 30830 27074
rect 30830 27022 30882 27074
rect 30882 27022 30884 27074
rect 30828 27020 30884 27022
rect 30716 26962 30772 26964
rect 30716 26910 30718 26962
rect 30718 26910 30770 26962
rect 30770 26910 30772 26962
rect 30716 26908 30772 26910
rect 32732 33234 32788 33236
rect 32732 33182 32734 33234
rect 32734 33182 32786 33234
rect 32786 33182 32788 33234
rect 32732 33180 32788 33182
rect 33404 30994 33460 30996
rect 33404 30942 33406 30994
rect 33406 30942 33458 30994
rect 33458 30942 33460 30994
rect 33404 30940 33460 30942
rect 39788 40124 39844 40180
rect 37996 39004 38052 39060
rect 41580 39676 41636 39732
rect 40348 39564 40404 39620
rect 39228 39058 39284 39060
rect 39228 39006 39230 39058
rect 39230 39006 39282 39058
rect 39282 39006 39284 39058
rect 39228 39004 39284 39006
rect 40460 39506 40516 39508
rect 40460 39454 40462 39506
rect 40462 39454 40514 39506
rect 40514 39454 40516 39506
rect 40460 39452 40516 39454
rect 41468 39618 41524 39620
rect 41468 39566 41470 39618
rect 41470 39566 41522 39618
rect 41522 39566 41524 39618
rect 41468 39564 41524 39566
rect 41692 39506 41748 39508
rect 41692 39454 41694 39506
rect 41694 39454 41746 39506
rect 41746 39454 41748 39506
rect 41692 39452 41748 39454
rect 41132 39004 41188 39060
rect 38332 38892 38388 38948
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34412 33068 34468 33124
rect 35420 32956 35476 33012
rect 37436 36988 37492 37044
rect 37772 36988 37828 37044
rect 36652 34972 36708 35028
rect 36092 33346 36148 33348
rect 36092 33294 36094 33346
rect 36094 33294 36146 33346
rect 36146 33294 36148 33346
rect 36092 33292 36148 33294
rect 35756 33234 35812 33236
rect 35756 33182 35758 33234
rect 35758 33182 35810 33234
rect 35810 33182 35812 33234
rect 35756 33180 35812 33182
rect 36316 32844 36372 32900
rect 35532 32732 35588 32788
rect 35980 32508 36036 32564
rect 34748 32060 34804 32116
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 33516 30098 33572 30100
rect 33516 30046 33518 30098
rect 33518 30046 33570 30098
rect 33570 30046 33572 30098
rect 33516 30044 33572 30046
rect 33628 31500 33684 31556
rect 33628 29820 33684 29876
rect 32732 29148 32788 29204
rect 32508 28642 32564 28644
rect 32508 28590 32510 28642
rect 32510 28590 32562 28642
rect 32562 28590 32564 28642
rect 32508 28588 32564 28590
rect 34636 28924 34692 28980
rect 34636 28642 34692 28644
rect 34636 28590 34638 28642
rect 34638 28590 34690 28642
rect 34690 28590 34692 28642
rect 34636 28588 34692 28590
rect 32844 27020 32900 27076
rect 31836 26850 31892 26852
rect 31836 26798 31838 26850
rect 31838 26798 31890 26850
rect 31890 26798 31892 26850
rect 31836 26796 31892 26798
rect 32060 26124 32116 26180
rect 30268 25788 30324 25844
rect 31276 25004 31332 25060
rect 31500 24610 31556 24612
rect 31500 24558 31502 24610
rect 31502 24558 31554 24610
rect 31554 24558 31556 24610
rect 31500 24556 31556 24558
rect 30156 23884 30212 23940
rect 28588 22204 28644 22260
rect 25788 20188 25844 20244
rect 25788 20018 25844 20020
rect 25788 19966 25790 20018
rect 25790 19966 25842 20018
rect 25842 19966 25844 20018
rect 25788 19964 25844 19966
rect 27132 19964 27188 20020
rect 26684 19740 26740 19796
rect 27132 19346 27188 19348
rect 27132 19294 27134 19346
rect 27134 19294 27186 19346
rect 27186 19294 27188 19346
rect 27132 19292 27188 19294
rect 27244 19068 27300 19124
rect 26012 16828 26068 16884
rect 24220 16044 24276 16100
rect 22428 15932 22484 15988
rect 23324 15986 23380 15988
rect 23324 15934 23326 15986
rect 23326 15934 23378 15986
rect 23378 15934 23380 15986
rect 23324 15932 23380 15934
rect 22764 15314 22820 15316
rect 22764 15262 22766 15314
rect 22766 15262 22818 15314
rect 22818 15262 22820 15314
rect 22764 15260 22820 15262
rect 23100 15314 23156 15316
rect 23100 15262 23102 15314
rect 23102 15262 23154 15314
rect 23154 15262 23156 15314
rect 23100 15260 23156 15262
rect 23548 15484 23604 15540
rect 24108 15484 24164 15540
rect 23324 15314 23380 15316
rect 23324 15262 23326 15314
rect 23326 15262 23378 15314
rect 23378 15262 23380 15314
rect 23324 15260 23380 15262
rect 21980 12908 22036 12964
rect 23436 15148 23492 15204
rect 23996 15148 24052 15204
rect 24220 15314 24276 15316
rect 24220 15262 24222 15314
rect 24222 15262 24274 15314
rect 24274 15262 24276 15314
rect 24220 15260 24276 15262
rect 24556 15986 24612 15988
rect 24556 15934 24558 15986
rect 24558 15934 24610 15986
rect 24610 15934 24612 15986
rect 24556 15932 24612 15934
rect 24892 15986 24948 15988
rect 24892 15934 24894 15986
rect 24894 15934 24946 15986
rect 24946 15934 24948 15986
rect 24892 15932 24948 15934
rect 25452 15986 25508 15988
rect 25452 15934 25454 15986
rect 25454 15934 25506 15986
rect 25506 15934 25508 15986
rect 25452 15932 25508 15934
rect 25676 15986 25732 15988
rect 25676 15934 25678 15986
rect 25678 15934 25730 15986
rect 25730 15934 25732 15986
rect 25676 15932 25732 15934
rect 24444 15538 24500 15540
rect 24444 15486 24446 15538
rect 24446 15486 24498 15538
rect 24498 15486 24500 15538
rect 24444 15484 24500 15486
rect 25340 15372 25396 15428
rect 24444 15148 24500 15204
rect 26012 15484 26068 15540
rect 24780 15036 24836 15092
rect 23324 13692 23380 13748
rect 17724 10780 17780 10836
rect 18284 10610 18340 10612
rect 18284 10558 18286 10610
rect 18286 10558 18338 10610
rect 18338 10558 18340 10610
rect 18284 10556 18340 10558
rect 17836 10050 17892 10052
rect 17836 9998 17838 10050
rect 17838 9998 17890 10050
rect 17890 9998 17892 10050
rect 17836 9996 17892 9998
rect 16716 9436 16772 9492
rect 17388 9826 17444 9828
rect 17388 9774 17390 9826
rect 17390 9774 17442 9826
rect 17442 9774 17444 9826
rect 17388 9772 17444 9774
rect 16268 8764 16324 8820
rect 16716 9042 16772 9044
rect 16716 8990 16718 9042
rect 16718 8990 16770 9042
rect 16770 8990 16772 9042
rect 16716 8988 16772 8990
rect 15372 5122 15428 5124
rect 15372 5070 15374 5122
rect 15374 5070 15426 5122
rect 15426 5070 15428 5122
rect 15372 5068 15428 5070
rect 16156 5068 16212 5124
rect 17948 9772 18004 9828
rect 17948 9602 18004 9604
rect 17948 9550 17950 9602
rect 17950 9550 18002 9602
rect 18002 9550 18004 9602
rect 17948 9548 18004 9550
rect 17612 9212 17668 9268
rect 20300 10610 20356 10612
rect 20300 10558 20302 10610
rect 20302 10558 20354 10610
rect 20354 10558 20356 10610
rect 20300 10556 20356 10558
rect 19292 9996 19348 10052
rect 19068 9826 19124 9828
rect 19068 9774 19070 9826
rect 19070 9774 19122 9826
rect 19122 9774 19124 9826
rect 19068 9772 19124 9774
rect 19628 9996 19684 10052
rect 19852 9826 19908 9828
rect 19852 9774 19854 9826
rect 19854 9774 19906 9826
rect 19906 9774 19908 9826
rect 19852 9772 19908 9774
rect 18620 9436 18676 9492
rect 17836 9042 17892 9044
rect 17836 8990 17838 9042
rect 17838 8990 17890 9042
rect 17890 8990 17892 9042
rect 17836 8988 17892 8990
rect 16380 5516 16436 5572
rect 18956 5516 19012 5572
rect 16828 5068 16884 5124
rect 16828 4562 16884 4564
rect 16828 4510 16830 4562
rect 16830 4510 16882 4562
rect 16882 4510 16884 4562
rect 16828 4508 16884 4510
rect 18732 4562 18788 4564
rect 18732 4510 18734 4562
rect 18734 4510 18786 4562
rect 18786 4510 18788 4562
rect 18732 4508 18788 4510
rect 19180 4508 19236 4564
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20076 9212 20132 9268
rect 20412 10050 20468 10052
rect 20412 9998 20414 10050
rect 20414 9998 20466 10050
rect 20466 9998 20468 10050
rect 20412 9996 20468 9998
rect 20860 9996 20916 10052
rect 21084 9266 21140 9268
rect 21084 9214 21086 9266
rect 21086 9214 21138 9266
rect 21138 9214 21140 9266
rect 21084 9212 21140 9214
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 22092 12684 22148 12740
rect 21644 12124 21700 12180
rect 21868 11900 21924 11956
rect 24220 13746 24276 13748
rect 24220 13694 24222 13746
rect 24222 13694 24274 13746
rect 24274 13694 24276 13746
rect 24220 13692 24276 13694
rect 22204 12178 22260 12180
rect 22204 12126 22206 12178
rect 22206 12126 22258 12178
rect 22258 12126 22260 12178
rect 22204 12124 22260 12126
rect 22428 11954 22484 11956
rect 22428 11902 22430 11954
rect 22430 11902 22482 11954
rect 22482 11902 22484 11954
rect 22428 11900 22484 11902
rect 25900 15202 25956 15204
rect 25900 15150 25902 15202
rect 25902 15150 25954 15202
rect 25954 15150 25956 15202
rect 25900 15148 25956 15150
rect 24556 11340 24612 11396
rect 25116 11282 25172 11284
rect 25116 11230 25118 11282
rect 25118 11230 25170 11282
rect 25170 11230 25172 11282
rect 25116 11228 25172 11230
rect 24444 10834 24500 10836
rect 24444 10782 24446 10834
rect 24446 10782 24498 10834
rect 24498 10782 24500 10834
rect 24444 10780 24500 10782
rect 24668 10834 24724 10836
rect 24668 10782 24670 10834
rect 24670 10782 24722 10834
rect 24722 10782 24724 10834
rect 24668 10780 24724 10782
rect 24220 10722 24276 10724
rect 24220 10670 24222 10722
rect 24222 10670 24274 10722
rect 24274 10670 24276 10722
rect 24220 10668 24276 10670
rect 24668 9548 24724 9604
rect 25004 10892 25060 10948
rect 25452 11394 25508 11396
rect 25452 11342 25454 11394
rect 25454 11342 25506 11394
rect 25506 11342 25508 11394
rect 25452 11340 25508 11342
rect 25564 10834 25620 10836
rect 25564 10782 25566 10834
rect 25566 10782 25618 10834
rect 25618 10782 25620 10834
rect 25564 10780 25620 10782
rect 28700 19906 28756 19908
rect 28700 19854 28702 19906
rect 28702 19854 28754 19906
rect 28754 19854 28756 19906
rect 28700 19852 28756 19854
rect 29932 19852 29988 19908
rect 29260 19794 29316 19796
rect 29260 19742 29262 19794
rect 29262 19742 29314 19794
rect 29314 19742 29316 19794
rect 29260 19740 29316 19742
rect 29260 19346 29316 19348
rect 29260 19294 29262 19346
rect 29262 19294 29314 19346
rect 29314 19294 29316 19346
rect 29260 19292 29316 19294
rect 30044 19964 30100 20020
rect 31276 23996 31332 24052
rect 32060 24050 32116 24052
rect 32060 23998 32062 24050
rect 32062 23998 32114 24050
rect 32114 23998 32116 24050
rect 32060 23996 32116 23998
rect 32396 26796 32452 26852
rect 33292 26796 33348 26852
rect 32508 26236 32564 26292
rect 33516 26236 33572 26292
rect 33180 26178 33236 26180
rect 33180 26126 33182 26178
rect 33182 26126 33234 26178
rect 33234 26126 33236 26178
rect 33180 26124 33236 26126
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 36428 31388 36484 31444
rect 34972 30098 35028 30100
rect 34972 30046 34974 30098
rect 34974 30046 35026 30098
rect 35026 30046 35028 30098
rect 34972 30044 35028 30046
rect 37660 34972 37716 35028
rect 36876 32786 36932 32788
rect 36876 32734 36878 32786
rect 36878 32734 36930 32786
rect 36930 32734 36932 32786
rect 36876 32732 36932 32734
rect 37212 33180 37268 33236
rect 37324 32844 37380 32900
rect 36764 32562 36820 32564
rect 36764 32510 36766 32562
rect 36766 32510 36818 32562
rect 36818 32510 36820 32562
rect 36764 32508 36820 32510
rect 37548 32562 37604 32564
rect 37548 32510 37550 32562
rect 37550 32510 37602 32562
rect 37602 32510 37604 32562
rect 37548 32508 37604 32510
rect 37548 31948 37604 32004
rect 37436 31724 37492 31780
rect 36988 31388 37044 31444
rect 35644 29820 35700 29876
rect 34860 29148 34916 29204
rect 36316 29932 36372 29988
rect 34972 28418 35028 28420
rect 34972 28366 34974 28418
rect 34974 28366 35026 28418
rect 35026 28366 35028 28418
rect 34972 28364 35028 28366
rect 34748 25564 34804 25620
rect 32620 25116 32676 25172
rect 29932 19180 29988 19236
rect 30380 19964 30436 20020
rect 31388 20018 31444 20020
rect 31388 19966 31390 20018
rect 31390 19966 31442 20018
rect 31442 19966 31444 20018
rect 31388 19964 31444 19966
rect 30156 18956 30212 19012
rect 29484 18844 29540 18900
rect 31164 19010 31220 19012
rect 31164 18958 31166 19010
rect 31166 18958 31218 19010
rect 31218 18958 31220 19010
rect 31164 18956 31220 18958
rect 32060 19234 32116 19236
rect 32060 19182 32062 19234
rect 32062 19182 32114 19234
rect 32114 19182 32116 19234
rect 32060 19180 32116 19182
rect 32172 19122 32228 19124
rect 32172 19070 32174 19122
rect 32174 19070 32226 19122
rect 32226 19070 32228 19122
rect 32172 19068 32228 19070
rect 31388 18844 31444 18900
rect 32396 18284 32452 18340
rect 29260 16156 29316 16212
rect 28700 15874 28756 15876
rect 28700 15822 28702 15874
rect 28702 15822 28754 15874
rect 28754 15822 28756 15874
rect 28700 15820 28756 15822
rect 29372 17052 29428 17108
rect 29372 15820 29428 15876
rect 28028 15426 28084 15428
rect 28028 15374 28030 15426
rect 28030 15374 28082 15426
rect 28082 15374 28084 15426
rect 28028 15372 28084 15374
rect 31948 16210 32004 16212
rect 31948 16158 31950 16210
rect 31950 16158 32002 16210
rect 32002 16158 32004 16210
rect 31948 16156 32004 16158
rect 32508 15202 32564 15204
rect 32508 15150 32510 15202
rect 32510 15150 32562 15202
rect 32562 15150 32564 15202
rect 32508 15148 32564 15150
rect 34524 24556 34580 24612
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35980 28642 36036 28644
rect 35980 28590 35982 28642
rect 35982 28590 36034 28642
rect 36034 28590 36036 28642
rect 35980 28588 36036 28590
rect 36428 29820 36484 29876
rect 36988 30098 37044 30100
rect 36988 30046 36990 30098
rect 36990 30046 37042 30098
rect 37042 30046 37044 30098
rect 36988 30044 37044 30046
rect 37324 30098 37380 30100
rect 37324 30046 37326 30098
rect 37326 30046 37378 30098
rect 37378 30046 37380 30098
rect 37324 30044 37380 30046
rect 36652 29596 36708 29652
rect 36988 28364 37044 28420
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 36652 26908 36708 26964
rect 37324 26796 37380 26852
rect 36764 26402 36820 26404
rect 36764 26350 36766 26402
rect 36766 26350 36818 26402
rect 36818 26350 36820 26402
rect 36764 26348 36820 26350
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35980 25618 36036 25620
rect 35980 25566 35982 25618
rect 35982 25566 36034 25618
rect 36034 25566 36036 25618
rect 35980 25564 36036 25566
rect 36988 25564 37044 25620
rect 35868 24892 35924 24948
rect 34972 24444 35028 24500
rect 35532 24722 35588 24724
rect 35532 24670 35534 24722
rect 35534 24670 35586 24722
rect 35586 24670 35588 24722
rect 35532 24668 35588 24670
rect 34860 22988 34916 23044
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35420 23042 35476 23044
rect 35420 22990 35422 23042
rect 35422 22990 35474 23042
rect 35474 22990 35476 23042
rect 35420 22988 35476 22990
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 20076 35252 20132
rect 37772 29596 37828 29652
rect 40124 38946 40180 38948
rect 40124 38894 40126 38946
rect 40126 38894 40178 38946
rect 40178 38894 40180 38946
rect 40124 38892 40180 38894
rect 40460 37996 40516 38052
rect 41020 38050 41076 38052
rect 41020 37998 41022 38050
rect 41022 37998 41074 38050
rect 41074 37998 41076 38050
rect 41020 37996 41076 37998
rect 42140 38220 42196 38276
rect 41916 37996 41972 38052
rect 39676 37772 39732 37828
rect 41244 37884 41300 37940
rect 40572 37826 40628 37828
rect 40572 37774 40574 37826
rect 40574 37774 40626 37826
rect 40626 37774 40628 37826
rect 40572 37772 40628 37774
rect 38108 36988 38164 37044
rect 38220 37154 38276 37156
rect 38220 37102 38222 37154
rect 38222 37102 38274 37154
rect 38274 37102 38276 37154
rect 38220 37100 38276 37102
rect 37996 33122 38052 33124
rect 37996 33070 37998 33122
rect 37998 33070 38050 33122
rect 38050 33070 38052 33122
rect 37996 33068 38052 33070
rect 38332 34972 38388 35028
rect 38892 34972 38948 35028
rect 41132 37212 41188 37268
rect 42700 37938 42756 37940
rect 42700 37886 42702 37938
rect 42702 37886 42754 37938
rect 42754 37886 42756 37938
rect 42700 37884 42756 37886
rect 43148 37938 43204 37940
rect 43148 37886 43150 37938
rect 43150 37886 43202 37938
rect 43202 37886 43204 37938
rect 43148 37884 43204 37886
rect 44044 37884 44100 37940
rect 40572 35026 40628 35028
rect 40572 34974 40574 35026
rect 40574 34974 40626 35026
rect 40626 34974 40628 35026
rect 40572 34972 40628 34974
rect 41020 34972 41076 35028
rect 41804 34972 41860 35028
rect 39788 32956 39844 33012
rect 40348 32284 40404 32340
rect 40012 31836 40068 31892
rect 38220 31724 38276 31780
rect 39004 31724 39060 31780
rect 38108 29932 38164 29988
rect 38220 29650 38276 29652
rect 38220 29598 38222 29650
rect 38222 29598 38274 29650
rect 38274 29598 38276 29650
rect 38220 29596 38276 29598
rect 37548 26962 37604 26964
rect 37548 26910 37550 26962
rect 37550 26910 37602 26962
rect 37602 26910 37604 26962
rect 37548 26908 37604 26910
rect 37772 26850 37828 26852
rect 37772 26798 37774 26850
rect 37774 26798 37826 26850
rect 37826 26798 37828 26850
rect 37772 26796 37828 26798
rect 38332 26348 38388 26404
rect 39676 31388 39732 31444
rect 42588 37826 42644 37828
rect 42588 37774 42590 37826
rect 42590 37774 42642 37826
rect 42642 37774 42644 37826
rect 42588 37772 42644 37774
rect 42140 37212 42196 37268
rect 43820 35026 43876 35028
rect 43820 34974 43822 35026
rect 43822 34974 43874 35026
rect 43874 34974 43876 35026
rect 43820 34972 43876 34974
rect 39340 30268 39396 30324
rect 39116 30098 39172 30100
rect 39116 30046 39118 30098
rect 39118 30046 39170 30098
rect 39170 30046 39172 30098
rect 39116 30044 39172 30046
rect 40348 30994 40404 30996
rect 40348 30942 40350 30994
rect 40350 30942 40402 30994
rect 40402 30942 40404 30994
rect 40348 30940 40404 30942
rect 41132 30994 41188 30996
rect 41132 30942 41134 30994
rect 41134 30942 41186 30994
rect 41186 30942 41188 30994
rect 41132 30940 41188 30942
rect 40124 30268 40180 30324
rect 39452 29932 39508 29988
rect 41804 32284 41860 32340
rect 42252 32284 42308 32340
rect 41692 29932 41748 29988
rect 40348 29260 40404 29316
rect 41244 27916 41300 27972
rect 39228 26348 39284 26404
rect 39900 25004 39956 25060
rect 38780 24722 38836 24724
rect 38780 24670 38782 24722
rect 38782 24670 38834 24722
rect 38834 24670 38836 24722
rect 38780 24668 38836 24670
rect 41692 27970 41748 27972
rect 41692 27918 41694 27970
rect 41694 27918 41746 27970
rect 41746 27918 41748 27970
rect 41692 27916 41748 27918
rect 41804 27804 41860 27860
rect 41244 26796 41300 26852
rect 41132 26178 41188 26180
rect 41132 26126 41134 26178
rect 41134 26126 41186 26178
rect 41186 26126 41188 26178
rect 41132 26124 41188 26126
rect 40236 24668 40292 24724
rect 40348 24556 40404 24612
rect 41580 27580 41636 27636
rect 41580 27132 41636 27188
rect 41804 27244 41860 27300
rect 40908 25004 40964 25060
rect 41132 25116 41188 25172
rect 40908 24556 40964 24612
rect 39452 22092 39508 22148
rect 37548 20802 37604 20804
rect 37548 20750 37550 20802
rect 37550 20750 37602 20802
rect 37602 20750 37604 20802
rect 37548 20748 37604 20750
rect 38780 20748 38836 20804
rect 36092 20300 36148 20356
rect 35084 19964 35140 20020
rect 35644 20130 35700 20132
rect 35644 20078 35646 20130
rect 35646 20078 35698 20130
rect 35698 20078 35700 20130
rect 35644 20076 35700 20078
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 33180 18338 33236 18340
rect 33180 18286 33182 18338
rect 33182 18286 33234 18338
rect 33234 18286 33236 18338
rect 33180 18284 33236 18286
rect 32956 17164 33012 17220
rect 32956 16940 33012 16996
rect 33180 17052 33236 17108
rect 32732 16156 32788 16212
rect 31836 14812 31892 14868
rect 25340 10722 25396 10724
rect 25340 10670 25342 10722
rect 25342 10670 25394 10722
rect 25394 10670 25396 10722
rect 25340 10668 25396 10670
rect 26348 11282 26404 11284
rect 26348 11230 26350 11282
rect 26350 11230 26402 11282
rect 26402 11230 26404 11282
rect 26348 11228 26404 11230
rect 26124 10780 26180 10836
rect 26684 10834 26740 10836
rect 26684 10782 26686 10834
rect 26686 10782 26738 10834
rect 26738 10782 26740 10834
rect 26684 10780 26740 10782
rect 26012 10668 26068 10724
rect 27020 10722 27076 10724
rect 27020 10670 27022 10722
rect 27022 10670 27074 10722
rect 27074 10670 27076 10722
rect 27020 10668 27076 10670
rect 28588 10668 28644 10724
rect 24892 9938 24948 9940
rect 24892 9886 24894 9938
rect 24894 9886 24946 9938
rect 24946 9886 24948 9938
rect 24892 9884 24948 9886
rect 26460 9938 26516 9940
rect 26460 9886 26462 9938
rect 26462 9886 26514 9938
rect 26514 9886 26516 9938
rect 26460 9884 26516 9886
rect 25788 9826 25844 9828
rect 25788 9774 25790 9826
rect 25790 9774 25842 9826
rect 25842 9774 25844 9826
rect 25788 9772 25844 9774
rect 23996 9266 24052 9268
rect 23996 9214 23998 9266
rect 23998 9214 24050 9266
rect 24050 9214 24052 9266
rect 23996 9212 24052 9214
rect 24556 9154 24612 9156
rect 24556 9102 24558 9154
rect 24558 9102 24610 9154
rect 24610 9102 24612 9154
rect 24556 9100 24612 9102
rect 25004 8988 25060 9044
rect 24668 8930 24724 8932
rect 24668 8878 24670 8930
rect 24670 8878 24722 8930
rect 24722 8878 24724 8930
rect 24668 8876 24724 8878
rect 25452 8876 25508 8932
rect 21756 6466 21812 6468
rect 21756 6414 21758 6466
rect 21758 6414 21810 6466
rect 21810 6414 21812 6466
rect 21756 6412 21812 6414
rect 23436 6412 23492 6468
rect 20412 4956 20468 5012
rect 31612 13746 31668 13748
rect 31612 13694 31614 13746
rect 31614 13694 31666 13746
rect 31666 13694 31668 13746
rect 31612 13692 31668 13694
rect 31612 11564 31668 11620
rect 31612 11394 31668 11396
rect 31612 11342 31614 11394
rect 31614 11342 31666 11394
rect 31666 11342 31668 11394
rect 31612 11340 31668 11342
rect 31276 11004 31332 11060
rect 29708 10780 29764 10836
rect 31948 11564 32004 11620
rect 31836 11452 31892 11508
rect 31724 11004 31780 11060
rect 33404 15148 33460 15204
rect 33068 14812 33124 14868
rect 32396 13746 32452 13748
rect 32396 13694 32398 13746
rect 32398 13694 32450 13746
rect 32450 13694 32452 13746
rect 32396 13692 32452 13694
rect 32060 11340 32116 11396
rect 32396 11452 32452 11508
rect 29260 9772 29316 9828
rect 25900 9548 25956 9604
rect 25676 9042 25732 9044
rect 25676 8990 25678 9042
rect 25678 8990 25730 9042
rect 25730 8990 25732 9042
rect 25676 8988 25732 8990
rect 26124 9154 26180 9156
rect 26124 9102 26126 9154
rect 26126 9102 26178 9154
rect 26178 9102 26180 9154
rect 26124 9100 26180 9102
rect 26572 9154 26628 9156
rect 26572 9102 26574 9154
rect 26574 9102 26626 9154
rect 26626 9102 26628 9154
rect 26572 9100 26628 9102
rect 28140 9100 28196 9156
rect 32732 11394 32788 11396
rect 32732 11342 32734 11394
rect 32734 11342 32786 11394
rect 32786 11342 32788 11394
rect 32732 11340 32788 11342
rect 32956 11394 33012 11396
rect 32956 11342 32958 11394
rect 32958 11342 33010 11394
rect 33010 11342 33012 11394
rect 32956 11340 33012 11342
rect 37548 20076 37604 20132
rect 35980 20018 36036 20020
rect 35980 19966 35982 20018
rect 35982 19966 36034 20018
rect 36034 19966 36036 20018
rect 35980 19964 36036 19966
rect 38892 20300 38948 20356
rect 39004 19964 39060 20020
rect 35756 18284 35812 18340
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34860 16828 34916 16884
rect 37996 19234 38052 19236
rect 37996 19182 37998 19234
rect 37998 19182 38050 19234
rect 38050 19182 38052 19234
rect 37996 19180 38052 19182
rect 38668 19234 38724 19236
rect 38668 19182 38670 19234
rect 38670 19182 38722 19234
rect 38722 19182 38724 19234
rect 38668 19180 38724 19182
rect 35756 16828 35812 16884
rect 36428 17164 36484 17220
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35756 13916 35812 13972
rect 35756 13746 35812 13748
rect 35756 13694 35758 13746
rect 35758 13694 35810 13746
rect 35810 13694 35812 13746
rect 35756 13692 35812 13694
rect 35868 13804 35924 13860
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34636 11340 34692 11396
rect 36204 13580 36260 13636
rect 36204 11394 36260 11396
rect 36204 11342 36206 11394
rect 36206 11342 36258 11394
rect 36258 11342 36260 11394
rect 36204 11340 36260 11342
rect 32620 11116 32676 11172
rect 34524 11170 34580 11172
rect 34524 11118 34526 11170
rect 34526 11118 34578 11170
rect 34578 11118 34580 11170
rect 34524 11116 34580 11118
rect 34188 11004 34244 11060
rect 35756 11004 35812 11060
rect 32508 10780 32564 10836
rect 33180 10834 33236 10836
rect 33180 10782 33182 10834
rect 33182 10782 33234 10834
rect 33234 10782 33236 10834
rect 33180 10780 33236 10782
rect 35084 10834 35140 10836
rect 35084 10782 35086 10834
rect 35086 10782 35138 10834
rect 35138 10782 35140 10834
rect 35084 10780 35140 10782
rect 35532 10780 35588 10836
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 31388 9548 31444 9604
rect 37548 17666 37604 17668
rect 37548 17614 37550 17666
rect 37550 17614 37602 17666
rect 37602 17614 37604 17666
rect 37548 17612 37604 17614
rect 37100 17164 37156 17220
rect 38108 16828 38164 16884
rect 36428 14530 36484 14532
rect 36428 14478 36430 14530
rect 36430 14478 36482 14530
rect 36482 14478 36484 14530
rect 36428 14476 36484 14478
rect 36764 13916 36820 13972
rect 36540 13746 36596 13748
rect 36540 13694 36542 13746
rect 36542 13694 36594 13746
rect 36594 13694 36596 13746
rect 36540 13692 36596 13694
rect 37436 13858 37492 13860
rect 37436 13806 37438 13858
rect 37438 13806 37490 13858
rect 37490 13806 37492 13858
rect 37436 13804 37492 13806
rect 37324 13746 37380 13748
rect 37324 13694 37326 13746
rect 37326 13694 37378 13746
rect 37378 13694 37380 13746
rect 37324 13692 37380 13694
rect 37212 13580 37268 13636
rect 37660 14476 37716 14532
rect 37996 13804 38052 13860
rect 37660 12908 37716 12964
rect 37548 12012 37604 12068
rect 36428 11452 36484 11508
rect 36988 11170 37044 11172
rect 36988 11118 36990 11170
rect 36990 11118 37042 11170
rect 37042 11118 37044 11170
rect 36988 11116 37044 11118
rect 36316 10780 36372 10836
rect 37660 11452 37716 11508
rect 37548 11394 37604 11396
rect 37548 11342 37550 11394
rect 37550 11342 37602 11394
rect 37602 11342 37604 11394
rect 37548 11340 37604 11342
rect 37100 9548 37156 9604
rect 30940 8988 30996 9044
rect 35084 9042 35140 9044
rect 35084 8990 35086 9042
rect 35086 8990 35138 9042
rect 35138 8990 35140 9042
rect 35084 8988 35140 8990
rect 39564 17778 39620 17780
rect 39564 17726 39566 17778
rect 39566 17726 39618 17778
rect 39618 17726 39620 17778
rect 39564 17724 39620 17726
rect 40908 24050 40964 24052
rect 40908 23998 40910 24050
rect 40910 23998 40962 24050
rect 40962 23998 40964 24050
rect 40908 23996 40964 23998
rect 41468 24444 41524 24500
rect 43596 30322 43652 30324
rect 43596 30270 43598 30322
rect 43598 30270 43650 30322
rect 43650 30270 43652 30322
rect 43596 30268 43652 30270
rect 42140 27244 42196 27300
rect 42028 26124 42084 26180
rect 43932 27186 43988 27188
rect 43932 27134 43934 27186
rect 43934 27134 43986 27186
rect 43986 27134 43988 27186
rect 43932 27132 43988 27134
rect 41916 24444 41972 24500
rect 43708 24444 43764 24500
rect 41692 23996 41748 24052
rect 40460 22146 40516 22148
rect 40460 22094 40462 22146
rect 40462 22094 40514 22146
rect 40514 22094 40516 22146
rect 40460 22092 40516 22094
rect 40908 22092 40964 22148
rect 39676 17612 39732 17668
rect 39676 16940 39732 16996
rect 39900 17724 39956 17780
rect 40236 17106 40292 17108
rect 40236 17054 40238 17106
rect 40238 17054 40290 17106
rect 40290 17054 40292 17106
rect 40236 17052 40292 17054
rect 40124 16994 40180 16996
rect 40124 16942 40126 16994
rect 40126 16942 40178 16994
rect 40178 16942 40180 16994
rect 40124 16940 40180 16942
rect 40908 17724 40964 17780
rect 41580 17724 41636 17780
rect 41468 17106 41524 17108
rect 41468 17054 41470 17106
rect 41470 17054 41522 17106
rect 41522 17054 41524 17106
rect 41468 17052 41524 17054
rect 41244 16994 41300 16996
rect 41244 16942 41246 16994
rect 41246 16942 41298 16994
rect 41298 16942 41300 16994
rect 41244 16940 41300 16942
rect 39900 13970 39956 13972
rect 39900 13918 39902 13970
rect 39902 13918 39954 13970
rect 39954 13918 39956 13970
rect 39900 13916 39956 13918
rect 40348 13634 40404 13636
rect 40348 13582 40350 13634
rect 40350 13582 40402 13634
rect 40402 13582 40404 13634
rect 40348 13580 40404 13582
rect 38444 13020 38500 13076
rect 40124 13074 40180 13076
rect 40124 13022 40126 13074
rect 40126 13022 40178 13074
rect 40178 13022 40180 13074
rect 40124 13020 40180 13022
rect 40236 12348 40292 12404
rect 43820 17778 43876 17780
rect 43820 17726 43822 17778
rect 43822 17726 43874 17778
rect 43874 17726 43876 17778
rect 43820 17724 43876 17726
rect 41020 13916 41076 13972
rect 41356 13580 41412 13636
rect 41020 12962 41076 12964
rect 41020 12910 41022 12962
rect 41022 12910 41074 12962
rect 41074 12910 41076 12962
rect 41020 12908 41076 12910
rect 43932 13634 43988 13636
rect 43932 13582 43934 13634
rect 43934 13582 43986 13634
rect 43986 13582 43988 13634
rect 43932 13580 43988 13582
rect 41020 12402 41076 12404
rect 41020 12350 41022 12402
rect 41022 12350 41074 12402
rect 41074 12350 41076 12402
rect 41020 12348 41076 12350
rect 38444 12012 38500 12068
rect 38332 9042 38388 9044
rect 38332 8990 38334 9042
rect 38334 8990 38386 9042
rect 38386 8990 38388 9042
rect 38332 8988 38388 8990
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 24108 5122 24164 5124
rect 24108 5070 24110 5122
rect 24110 5070 24162 5122
rect 24162 5070 24164 5122
rect 24108 5068 24164 5070
rect 24780 5068 24836 5124
rect 22204 4956 22260 5012
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
<< metal3 >>
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 13234 41916 13244 41972
rect 13300 41916 14476 41972
rect 14532 41916 14542 41972
rect 23202 41916 23212 41972
rect 23268 41916 28700 41972
rect 28756 41916 28766 41972
rect 31378 41916 31388 41972
rect 31444 41916 32508 41972
rect 32564 41916 32574 41972
rect 20850 41804 20860 41860
rect 20916 41804 22092 41860
rect 22148 41804 22158 41860
rect 24658 41804 24668 41860
rect 24724 41804 25900 41860
rect 25956 41804 25966 41860
rect 28466 41804 28476 41860
rect 28532 41804 29708 41860
rect 29764 41804 29774 41860
rect 36082 41804 36092 41860
rect 36148 41804 37324 41860
rect 37380 41804 37390 41860
rect 39890 41804 39900 41860
rect 39956 41804 41132 41860
rect 41188 41804 41198 41860
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 5170 40908 5180 40964
rect 5236 40908 6300 40964
rect 6356 40908 10780 40964
rect 10836 40908 13916 40964
rect 13972 40908 13982 40964
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 10434 40572 10444 40628
rect 10500 40572 32620 40628
rect 32676 40572 34188 40628
rect 34244 40572 34254 40628
rect 8082 40460 8092 40516
rect 8148 40460 10220 40516
rect 10276 40460 10286 40516
rect 3266 40348 3276 40404
rect 3332 40348 5180 40404
rect 5236 40348 5246 40404
rect 6178 40348 6188 40404
rect 6244 40348 8764 40404
rect 8820 40348 8830 40404
rect 14018 40348 14028 40404
rect 14084 40348 17052 40404
rect 17108 40348 17612 40404
rect 17668 40348 19740 40404
rect 19796 40348 20076 40404
rect 20132 40348 20142 40404
rect 25330 40348 25340 40404
rect 25396 40348 28476 40404
rect 28532 40348 28542 40404
rect 33394 40348 33404 40404
rect 33460 40348 33470 40404
rect 33404 40292 33460 40348
rect 3714 40236 3724 40292
rect 3780 40236 6412 40292
rect 6468 40236 6478 40292
rect 13570 40236 13580 40292
rect 13636 40236 24892 40292
rect 24948 40236 24958 40292
rect 31490 40236 31500 40292
rect 31556 40236 34972 40292
rect 35028 40236 36876 40292
rect 36932 40236 37996 40292
rect 38052 40236 38062 40292
rect 5842 40124 5852 40180
rect 5908 40124 13468 40180
rect 13524 40124 13534 40180
rect 28354 40124 28364 40180
rect 28420 40124 39788 40180
rect 39844 40124 39854 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 10098 39788 10108 39844
rect 10164 39788 11228 39844
rect 11284 39788 11900 39844
rect 11956 39788 11966 39844
rect 9090 39676 9100 39732
rect 9156 39676 11788 39732
rect 11844 39676 11854 39732
rect 34402 39676 34412 39732
rect 34468 39676 41580 39732
rect 41636 39676 41646 39732
rect 9202 39564 9212 39620
rect 9268 39564 10220 39620
rect 10276 39564 10286 39620
rect 40338 39564 40348 39620
rect 40404 39564 41468 39620
rect 41524 39564 41534 39620
rect 6962 39452 6972 39508
rect 7028 39452 7644 39508
rect 7700 39452 10780 39508
rect 10836 39452 10846 39508
rect 11900 39452 21084 39508
rect 21140 39452 21150 39508
rect 40450 39452 40460 39508
rect 40516 39452 41692 39508
rect 41748 39452 41758 39508
rect 11900 39396 11956 39452
rect 6290 39340 6300 39396
rect 6356 39340 7532 39396
rect 7588 39340 8316 39396
rect 8372 39340 8382 39396
rect 8642 39340 8652 39396
rect 8708 39340 8718 39396
rect 9874 39340 9884 39396
rect 9940 39340 11956 39396
rect 12114 39340 12124 39396
rect 12180 39340 28252 39396
rect 28308 39340 29260 39396
rect 29316 39340 29326 39396
rect 8316 39172 8372 39340
rect 8652 39284 8708 39340
rect 8652 39228 18172 39284
rect 18228 39228 18238 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 8316 39116 9100 39172
rect 9156 39116 9548 39172
rect 9604 39116 9614 39172
rect 7298 39004 7308 39060
rect 7364 39004 7868 39060
rect 7924 39004 8540 39060
rect 8596 39004 8606 39060
rect 12114 39004 12124 39060
rect 12180 39004 13916 39060
rect 13972 39004 13982 39060
rect 37986 39004 37996 39060
rect 38052 39004 39228 39060
rect 39284 39004 41132 39060
rect 41188 39004 41198 39060
rect 2594 38892 2604 38948
rect 2660 38892 8876 38948
rect 8932 38892 9660 38948
rect 9716 38892 9726 38948
rect 10770 38892 10780 38948
rect 10836 38892 11676 38948
rect 11732 38892 11742 38948
rect 38322 38892 38332 38948
rect 38388 38892 40124 38948
rect 40180 38892 40190 38948
rect 8978 38780 8988 38836
rect 9044 38780 9884 38836
rect 9940 38780 10556 38836
rect 10612 38780 10622 38836
rect 10780 38780 11228 38836
rect 11284 38780 11294 38836
rect 10780 38612 10836 38780
rect 10098 38556 10108 38612
rect 10164 38556 10836 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 42130 38220 42140 38276
rect 42196 38220 42206 38276
rect 42140 38052 42196 38220
rect 40450 37996 40460 38052
rect 40516 37996 41020 38052
rect 41076 37996 41086 38052
rect 41906 37996 41916 38052
rect 41972 37996 42196 38052
rect 21858 37884 21868 37940
rect 21924 37884 24892 37940
rect 24948 37884 24958 37940
rect 39676 37884 41244 37940
rect 41300 37884 42700 37940
rect 42756 37884 43148 37940
rect 43204 37884 43214 37940
rect 43652 37884 44044 37940
rect 44100 37884 44110 37940
rect 39676 37828 39732 37884
rect 43652 37828 43708 37884
rect 11442 37772 11452 37828
rect 11508 37772 12124 37828
rect 12180 37772 12190 37828
rect 25778 37772 25788 37828
rect 25844 37772 26348 37828
rect 26404 37772 39676 37828
rect 39732 37772 39742 37828
rect 40562 37772 40572 37828
rect 40628 37772 42588 37828
rect 42644 37772 43708 37828
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 24322 37324 24332 37380
rect 24388 37324 25564 37380
rect 25620 37324 25630 37380
rect 27570 37324 27580 37380
rect 27636 37324 28476 37380
rect 28532 37324 30268 37380
rect 30324 37324 30828 37380
rect 30884 37324 31724 37380
rect 31780 37324 31790 37380
rect 22978 37212 22988 37268
rect 23044 37212 24220 37268
rect 24276 37212 25228 37268
rect 25284 37212 25294 37268
rect 38612 37212 41132 37268
rect 41188 37212 42140 37268
rect 42196 37212 42206 37268
rect 38612 37156 38668 37212
rect 38210 37100 38220 37156
rect 38276 37100 38668 37156
rect 24546 36988 24556 37044
rect 24612 36988 37436 37044
rect 37492 36988 37772 37044
rect 37828 36988 38108 37044
rect 38164 36988 38174 37044
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 30370 36540 30380 36596
rect 30436 36540 30446 36596
rect 30380 36484 30436 36540
rect 17266 36428 17276 36484
rect 17332 36428 19068 36484
rect 19124 36428 19134 36484
rect 20514 36428 20524 36484
rect 20580 36428 24220 36484
rect 24276 36428 25564 36484
rect 25620 36428 25630 36484
rect 29474 36428 29484 36484
rect 29540 36428 30828 36484
rect 30884 36428 30894 36484
rect 15586 36316 15596 36372
rect 15652 36316 16940 36372
rect 16996 36316 17006 36372
rect 26786 36316 26796 36372
rect 26852 36316 29148 36372
rect 29204 36316 29214 36372
rect 4946 36204 4956 36260
rect 5012 36204 7196 36260
rect 7252 36204 9660 36260
rect 9716 36204 9726 36260
rect 16146 36204 16156 36260
rect 16212 36204 17724 36260
rect 17780 36204 17790 36260
rect 25666 36204 25676 36260
rect 25732 36204 26572 36260
rect 26628 36204 26908 36260
rect 26964 36204 26974 36260
rect 27458 36204 27468 36260
rect 27524 36204 28364 36260
rect 28420 36204 28430 36260
rect 17490 36092 17500 36148
rect 17556 36092 18060 36148
rect 18116 36092 19628 36148
rect 19684 36092 19694 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 2594 35756 2604 35812
rect 2660 35756 7644 35812
rect 7700 35756 7710 35812
rect 11218 35756 11228 35812
rect 11284 35756 16268 35812
rect 16324 35756 16334 35812
rect 18162 35756 18172 35812
rect 18228 35756 18620 35812
rect 18676 35756 20076 35812
rect 20132 35756 30380 35812
rect 30436 35756 30446 35812
rect 16370 35644 16380 35700
rect 16436 35644 17388 35700
rect 17444 35644 17454 35700
rect 17826 35644 17836 35700
rect 17892 35644 18732 35700
rect 18788 35644 19180 35700
rect 19236 35644 23660 35700
rect 23716 35644 23726 35700
rect 4722 35420 4732 35476
rect 4788 35420 9324 35476
rect 9380 35420 9390 35476
rect 10322 35420 10332 35476
rect 10388 35420 11564 35476
rect 11620 35420 14588 35476
rect 14644 35420 14654 35476
rect 14914 35420 14924 35476
rect 14980 35420 15708 35476
rect 15764 35420 16492 35476
rect 16548 35420 16558 35476
rect 17154 35420 17164 35476
rect 17220 35420 18620 35476
rect 18676 35420 18686 35476
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 10434 35196 10444 35252
rect 10500 35196 11116 35252
rect 11172 35196 14140 35252
rect 14196 35196 14206 35252
rect 7970 35084 7980 35140
rect 8036 35084 11396 35140
rect 15922 35084 15932 35140
rect 15988 35084 17724 35140
rect 17780 35084 17790 35140
rect 11340 35028 11396 35084
rect 4834 34972 4844 35028
rect 4900 34972 10220 35028
rect 10276 34972 10286 35028
rect 11330 34972 11340 35028
rect 11396 34972 11406 35028
rect 14690 34972 14700 35028
rect 14756 34972 15596 35028
rect 15652 34972 15662 35028
rect 36642 34972 36652 35028
rect 36708 34972 37660 35028
rect 37716 34972 38332 35028
rect 38388 34972 38892 35028
rect 38948 34972 40572 35028
rect 40628 34972 41020 35028
rect 41076 34972 41086 35028
rect 41794 34972 41804 35028
rect 41860 34972 43820 35028
rect 43876 34972 43886 35028
rect 10098 34860 10108 34916
rect 10164 34860 11116 34916
rect 11172 34860 11182 34916
rect 15362 34860 15372 34916
rect 15428 34860 16828 34916
rect 16884 34860 16894 34916
rect 30258 34860 30268 34916
rect 30324 34860 33516 34916
rect 33572 34860 33582 34916
rect 7074 34748 7084 34804
rect 7140 34748 14364 34804
rect 14420 34748 14430 34804
rect 25778 34748 25788 34804
rect 25844 34748 27356 34804
rect 27412 34748 27422 34804
rect 10098 34636 10108 34692
rect 10164 34636 10892 34692
rect 10948 34636 12348 34692
rect 12404 34636 15372 34692
rect 15428 34636 15438 34692
rect 23762 34636 23772 34692
rect 23828 34636 25676 34692
rect 25732 34636 25742 34692
rect 26002 34636 26012 34692
rect 26068 34636 27692 34692
rect 27748 34636 27758 34692
rect 9090 34524 9100 34580
rect 9156 34524 10444 34580
rect 10500 34524 10510 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 9538 34300 9548 34356
rect 9604 34300 10556 34356
rect 10612 34300 11340 34356
rect 11396 34300 11676 34356
rect 11732 34300 11742 34356
rect 31266 34300 31276 34356
rect 31332 34300 32060 34356
rect 32116 34300 33068 34356
rect 33124 34300 33134 34356
rect 27122 34188 27132 34244
rect 27188 34188 27916 34244
rect 27972 34188 27982 34244
rect 30380 34188 31612 34244
rect 31668 34188 31836 34244
rect 31892 34188 31902 34244
rect 30380 34132 30436 34188
rect 7074 34076 7084 34132
rect 7140 34076 14140 34132
rect 14196 34076 14206 34132
rect 26338 34076 26348 34132
rect 26404 34076 26908 34132
rect 26964 34076 27244 34132
rect 27300 34076 27310 34132
rect 27458 34076 27468 34132
rect 27524 34076 28028 34132
rect 28084 34076 30436 34132
rect 1922 33964 1932 34020
rect 1988 33964 4284 34020
rect 4340 33964 5180 34020
rect 5236 33964 7532 34020
rect 7588 33964 7598 34020
rect 14354 33852 14364 33908
rect 14420 33852 15260 33908
rect 15316 33852 15326 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 10210 33516 10220 33572
rect 10276 33516 10668 33572
rect 10724 33516 11452 33572
rect 11508 33516 17052 33572
rect 17108 33516 17118 33572
rect 17826 33404 17836 33460
rect 17892 33404 23100 33460
rect 23156 33404 23166 33460
rect 32946 33292 32956 33348
rect 33012 33292 36092 33348
rect 36148 33292 36158 33348
rect 23874 33180 23884 33236
rect 23940 33180 24668 33236
rect 24724 33180 24734 33236
rect 31602 33180 31612 33236
rect 31668 33180 32732 33236
rect 32788 33180 32798 33236
rect 35746 33180 35756 33236
rect 35812 33180 37212 33236
rect 37268 33180 37278 33236
rect 11666 33068 11676 33124
rect 11732 33068 12908 33124
rect 12964 33068 12974 33124
rect 26786 33068 26796 33124
rect 26852 33068 27468 33124
rect 27524 33068 27534 33124
rect 32386 33068 32396 33124
rect 32452 33068 34412 33124
rect 34468 33068 37996 33124
rect 38052 33068 38062 33124
rect 27122 32956 27132 33012
rect 27188 32956 28364 33012
rect 28420 32956 35420 33012
rect 35476 32956 39788 33012
rect 39844 32956 39854 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 36306 32844 36316 32900
rect 36372 32844 37324 32900
rect 37380 32844 37390 32900
rect 25106 32732 25116 32788
rect 25172 32732 31052 32788
rect 31108 32732 35532 32788
rect 35588 32732 36876 32788
rect 36932 32732 36942 32788
rect 15250 32508 15260 32564
rect 15316 32508 16940 32564
rect 16996 32508 17006 32564
rect 22866 32508 22876 32564
rect 22932 32508 23884 32564
rect 23940 32508 23950 32564
rect 24098 32508 24108 32564
rect 24164 32508 26684 32564
rect 26740 32508 26750 32564
rect 30258 32508 30268 32564
rect 30324 32508 31612 32564
rect 31668 32508 32284 32564
rect 32340 32508 32350 32564
rect 35970 32508 35980 32564
rect 36036 32508 36764 32564
rect 36820 32508 37548 32564
rect 37604 32508 37614 32564
rect 26562 32396 26572 32452
rect 26628 32396 27020 32452
rect 27076 32396 30044 32452
rect 30100 32396 30110 32452
rect 40338 32284 40348 32340
rect 40404 32284 41804 32340
rect 41860 32284 42252 32340
rect 42308 32284 42318 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 27010 32060 27020 32116
rect 27076 32060 34748 32116
rect 34804 32060 34814 32116
rect 26852 31948 30828 32004
rect 30884 31948 30894 32004
rect 37538 31948 37548 32004
rect 37604 31948 38668 32004
rect 26852 31892 26908 31948
rect 38612 31892 38668 31948
rect 25554 31836 25564 31892
rect 25620 31836 26908 31892
rect 27570 31836 27580 31892
rect 27636 31836 28252 31892
rect 28308 31836 28318 31892
rect 38612 31836 40012 31892
rect 40068 31836 40078 31892
rect 27580 31780 27636 31836
rect 12898 31724 12908 31780
rect 12964 31724 13580 31780
rect 13636 31724 23492 31780
rect 26674 31724 26684 31780
rect 26740 31724 27636 31780
rect 37426 31724 37436 31780
rect 37492 31724 38220 31780
rect 38276 31724 39004 31780
rect 39060 31724 39070 31780
rect 2930 31612 2940 31668
rect 2996 31612 4172 31668
rect 4228 31612 4238 31668
rect 13010 31612 13020 31668
rect 13076 31612 15148 31668
rect 15204 31612 18956 31668
rect 19012 31612 19022 31668
rect 2146 31500 2156 31556
rect 2212 31500 5740 31556
rect 5796 31500 7532 31556
rect 7588 31500 7598 31556
rect 14018 31500 14028 31556
rect 14084 31500 20748 31556
rect 20804 31500 21644 31556
rect 21700 31500 21710 31556
rect 23436 31444 23492 31724
rect 26450 31612 26460 31668
rect 26516 31612 27132 31668
rect 27188 31612 27198 31668
rect 24098 31500 24108 31556
rect 24164 31500 25564 31556
rect 25620 31500 25630 31556
rect 30034 31500 30044 31556
rect 30100 31500 30716 31556
rect 30772 31500 33628 31556
rect 33684 31500 33694 31556
rect 23426 31388 23436 31444
rect 23492 31388 36428 31444
rect 36484 31388 36988 31444
rect 37044 31388 39676 31444
rect 39732 31388 39742 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 30706 31052 30716 31108
rect 30772 31052 31500 31108
rect 31556 31052 31566 31108
rect 15922 30940 15932 30996
rect 15988 30940 17948 30996
rect 18004 30940 20188 30996
rect 30146 30940 30156 30996
rect 30212 30940 32508 30996
rect 32564 30940 33404 30996
rect 33460 30940 33470 30996
rect 40338 30940 40348 30996
rect 40404 30940 41132 30996
rect 41188 30940 41198 30996
rect 7522 30828 7532 30884
rect 7588 30828 9660 30884
rect 9716 30828 10892 30884
rect 10948 30828 10958 30884
rect 16818 30828 16828 30884
rect 16884 30828 17500 30884
rect 17556 30828 17566 30884
rect 20132 30828 20188 30940
rect 20244 30828 28588 30884
rect 28644 30828 28654 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 14354 30268 14364 30324
rect 14420 30268 14924 30324
rect 14980 30268 16156 30324
rect 16212 30268 16222 30324
rect 18946 30268 18956 30324
rect 19012 30268 19628 30324
rect 19684 30268 19694 30324
rect 21634 30268 21644 30324
rect 21700 30268 22540 30324
rect 22596 30268 22606 30324
rect 28578 30268 28588 30324
rect 28644 30268 30156 30324
rect 30212 30268 30222 30324
rect 39330 30268 39340 30324
rect 39396 30268 40124 30324
rect 40180 30268 43596 30324
rect 43652 30268 43662 30324
rect 29698 30156 29708 30212
rect 29764 30156 30604 30212
rect 30660 30156 30670 30212
rect 15698 30044 15708 30100
rect 15764 30044 18284 30100
rect 18340 30044 18350 30100
rect 28802 30044 28812 30100
rect 28868 30044 32060 30100
rect 32116 30044 33516 30100
rect 33572 30044 33582 30100
rect 34962 30044 34972 30100
rect 35028 30044 36988 30100
rect 37044 30044 37054 30100
rect 37314 30044 37324 30100
rect 37380 30044 39116 30100
rect 39172 30044 39182 30100
rect 36306 29932 36316 29988
rect 36372 29932 38108 29988
rect 38164 29932 39452 29988
rect 39508 29932 41692 29988
rect 41748 29932 41758 29988
rect 33618 29820 33628 29876
rect 33684 29820 35644 29876
rect 35700 29820 36428 29876
rect 36484 29820 36494 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 6850 29596 6860 29652
rect 6916 29596 11228 29652
rect 11284 29596 11294 29652
rect 11442 29596 11452 29652
rect 11508 29596 11900 29652
rect 11956 29596 14028 29652
rect 14084 29596 14094 29652
rect 36642 29596 36652 29652
rect 36708 29596 37772 29652
rect 37828 29596 38220 29652
rect 38276 29596 38668 29652
rect 38612 29316 38668 29596
rect 29474 29260 29484 29316
rect 29540 29260 30380 29316
rect 30436 29260 30446 29316
rect 38612 29260 40348 29316
rect 40404 29260 40414 29316
rect 32722 29148 32732 29204
rect 32788 29148 34860 29204
rect 34916 29148 34926 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 23202 28924 23212 28980
rect 23268 28924 26236 28980
rect 26292 28924 31948 28980
rect 32004 28924 34636 28980
rect 34692 28924 34702 28980
rect 2594 28812 2604 28868
rect 2660 28812 4508 28868
rect 4564 28812 4574 28868
rect 8372 28812 12852 28868
rect 26002 28812 26012 28868
rect 26068 28812 29820 28868
rect 29876 28812 29886 28868
rect 8372 28756 8428 28812
rect 12796 28756 12852 28812
rect 4274 28700 4284 28756
rect 4340 28700 5740 28756
rect 5796 28700 5806 28756
rect 6402 28700 6412 28756
rect 6468 28700 6972 28756
rect 7028 28700 8428 28756
rect 11666 28700 11676 28756
rect 11732 28700 12572 28756
rect 12628 28700 12638 28756
rect 12786 28700 12796 28756
rect 12852 28700 12862 28756
rect 20290 28700 20300 28756
rect 20356 28700 21308 28756
rect 21364 28700 21812 28756
rect 21970 28700 21980 28756
rect 22036 28700 22988 28756
rect 23044 28700 23996 28756
rect 24052 28700 24062 28756
rect 21756 28644 21812 28700
rect 9538 28588 9548 28644
rect 9604 28588 10332 28644
rect 10388 28588 11452 28644
rect 11508 28588 11518 28644
rect 12898 28588 12908 28644
rect 12964 28588 15148 28644
rect 15204 28588 16716 28644
rect 16772 28588 16782 28644
rect 17266 28588 17276 28644
rect 17332 28588 21532 28644
rect 21588 28588 21598 28644
rect 21756 28588 22316 28644
rect 22372 28588 23100 28644
rect 23156 28588 23166 28644
rect 29922 28588 29932 28644
rect 29988 28588 32508 28644
rect 32564 28588 32574 28644
rect 34626 28588 34636 28644
rect 34692 28588 35980 28644
rect 36036 28588 36046 28644
rect 5058 28476 5068 28532
rect 5124 28476 7756 28532
rect 7812 28476 7822 28532
rect 15922 28476 15932 28532
rect 15988 28476 17388 28532
rect 17444 28476 17454 28532
rect 4050 28364 4060 28420
rect 4116 28364 5628 28420
rect 5684 28364 5694 28420
rect 11890 28364 11900 28420
rect 11956 28364 12460 28420
rect 12516 28364 12526 28420
rect 31938 28364 31948 28420
rect 32004 28364 34972 28420
rect 35028 28364 36988 28420
rect 37044 28364 37054 28420
rect 4610 28252 4620 28308
rect 4676 28252 5516 28308
rect 5572 28252 5582 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4946 28140 4956 28196
rect 5012 28140 5404 28196
rect 5460 28140 5470 28196
rect 4834 28028 4844 28084
rect 4900 28028 5628 28084
rect 5684 28028 9996 28084
rect 10052 28028 10062 28084
rect 22642 28028 22652 28084
rect 22708 28028 23660 28084
rect 23716 28028 25340 28084
rect 25396 28028 28588 28084
rect 28644 28028 28812 28084
rect 28868 28028 28878 28084
rect 11890 27916 11900 27972
rect 11956 27916 15372 27972
rect 15428 27916 16492 27972
rect 16548 27916 16558 27972
rect 17154 27916 17164 27972
rect 17220 27916 17230 27972
rect 41234 27916 41244 27972
rect 41300 27916 41692 27972
rect 41748 27916 41758 27972
rect 17164 27860 17220 27916
rect 11666 27804 11676 27860
rect 11732 27804 15148 27860
rect 15204 27804 16604 27860
rect 16660 27804 17220 27860
rect 28578 27804 28588 27860
rect 28644 27804 28924 27860
rect 28980 27804 30156 27860
rect 30212 27804 30222 27860
rect 41580 27804 41804 27860
rect 41860 27804 41870 27860
rect 17154 27692 17164 27748
rect 17220 27692 19740 27748
rect 19796 27692 19806 27748
rect 28130 27692 28140 27748
rect 28196 27692 29372 27748
rect 29428 27692 29438 27748
rect 41580 27636 41636 27804
rect 41570 27580 41580 27636
rect 41636 27580 41646 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 41794 27244 41804 27300
rect 41860 27244 42140 27300
rect 42196 27244 42206 27300
rect 8754 27132 8764 27188
rect 8820 27132 10892 27188
rect 10948 27132 12124 27188
rect 12180 27132 17724 27188
rect 17780 27132 17790 27188
rect 41570 27132 41580 27188
rect 41636 27132 43932 27188
rect 43988 27132 43998 27188
rect 8978 27020 8988 27076
rect 9044 27020 9884 27076
rect 9940 27020 9950 27076
rect 12562 27020 12572 27076
rect 12628 27020 14140 27076
rect 14196 27020 14206 27076
rect 15362 27020 15372 27076
rect 15428 27020 17164 27076
rect 17220 27020 17230 27076
rect 30818 27020 30828 27076
rect 30884 27020 32844 27076
rect 32900 27020 32910 27076
rect 11554 26908 11564 26964
rect 11620 26908 12684 26964
rect 12740 26908 12750 26964
rect 29362 26908 29372 26964
rect 29428 26908 30716 26964
rect 30772 26908 30782 26964
rect 36642 26908 36652 26964
rect 36708 26908 37548 26964
rect 37604 26908 37614 26964
rect 14466 26796 14476 26852
rect 14532 26796 22652 26852
rect 22708 26796 22718 26852
rect 23874 26796 23884 26852
rect 23940 26796 26124 26852
rect 26180 26796 26190 26852
rect 31826 26796 31836 26852
rect 31892 26796 32396 26852
rect 32452 26796 33292 26852
rect 33348 26796 33358 26852
rect 37314 26796 37324 26852
rect 37380 26796 37772 26852
rect 37828 26796 41244 26852
rect 41300 26796 41310 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 5282 26460 5292 26516
rect 5348 26460 6412 26516
rect 6468 26460 6478 26516
rect 12226 26460 12236 26516
rect 12292 26460 13132 26516
rect 13188 26460 18732 26516
rect 18788 26460 21644 26516
rect 21700 26460 23100 26516
rect 23156 26460 23166 26516
rect 5842 26348 5852 26404
rect 5908 26348 6076 26404
rect 6132 26348 10780 26404
rect 10836 26348 11900 26404
rect 11956 26348 11966 26404
rect 36754 26348 36764 26404
rect 36820 26348 38332 26404
rect 38388 26348 39228 26404
rect 39284 26348 39294 26404
rect 4610 26236 4620 26292
rect 4676 26236 6300 26292
rect 6356 26236 6366 26292
rect 10546 26236 10556 26292
rect 10612 26236 11452 26292
rect 11508 26236 11518 26292
rect 13570 26236 13580 26292
rect 13636 26236 15708 26292
rect 15764 26236 16604 26292
rect 16660 26236 17388 26292
rect 17444 26236 17454 26292
rect 32498 26236 32508 26292
rect 32564 26236 33516 26292
rect 33572 26236 33582 26292
rect 32050 26124 32060 26180
rect 32116 26124 33180 26180
rect 33236 26124 33246 26180
rect 41122 26124 41132 26180
rect 41188 26124 42028 26180
rect 42084 26124 42094 26180
rect 4274 26012 4284 26068
rect 4340 26012 15148 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 15092 25844 15148 26012
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 15092 25788 20188 25844
rect 26002 25788 26012 25844
rect 26068 25788 30268 25844
rect 30324 25788 30334 25844
rect 9202 25676 9212 25732
rect 9268 25676 10444 25732
rect 10500 25676 10780 25732
rect 10836 25676 11004 25732
rect 11060 25676 11070 25732
rect 11330 25676 11340 25732
rect 11396 25676 12908 25732
rect 12964 25676 13580 25732
rect 13636 25676 13646 25732
rect 20132 25620 20188 25788
rect 8306 25564 8316 25620
rect 8372 25564 10556 25620
rect 10612 25564 10622 25620
rect 14018 25564 14028 25620
rect 14084 25564 14588 25620
rect 14644 25564 14654 25620
rect 20132 25564 25228 25620
rect 25284 25564 28924 25620
rect 28980 25564 28990 25620
rect 34738 25564 34748 25620
rect 34804 25564 35980 25620
rect 36036 25564 36988 25620
rect 37044 25564 37054 25620
rect 4834 25452 4844 25508
rect 4900 25452 5516 25508
rect 5572 25452 6188 25508
rect 6244 25452 7196 25508
rect 7252 25452 7262 25508
rect 8194 25452 8204 25508
rect 8260 25452 9548 25508
rect 9604 25452 9614 25508
rect 14354 25452 14364 25508
rect 14420 25452 15148 25508
rect 15204 25452 15214 25508
rect 23090 25452 23100 25508
rect 23156 25452 23772 25508
rect 23828 25452 24220 25508
rect 24276 25452 24286 25508
rect 5730 25340 5740 25396
rect 5796 25340 6412 25396
rect 6468 25340 11004 25396
rect 11060 25340 15708 25396
rect 15764 25340 15774 25396
rect 21410 25340 21420 25396
rect 21476 25340 23884 25396
rect 23940 25340 23950 25396
rect 4834 25228 4844 25284
rect 4900 25228 5852 25284
rect 5908 25228 5918 25284
rect 6178 25228 6188 25284
rect 6244 25228 10668 25284
rect 10724 25228 10734 25284
rect 23426 25228 23436 25284
rect 23492 25228 24892 25284
rect 24948 25228 25564 25284
rect 25620 25228 25630 25284
rect 27356 25116 32620 25172
rect 32676 25116 32686 25172
rect 39676 25116 41132 25172
rect 41188 25116 41198 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 5282 25004 5292 25060
rect 5348 25004 5908 25060
rect 9650 25004 9660 25060
rect 9716 25004 10556 25060
rect 10612 25004 11116 25060
rect 11172 25004 18060 25060
rect 18116 25004 18126 25060
rect 5852 24948 5908 25004
rect 4050 24892 4060 24948
rect 4116 24892 5068 24948
rect 5124 24892 5134 24948
rect 5842 24892 5852 24948
rect 5908 24892 7868 24948
rect 7924 24892 8764 24948
rect 8820 24892 8830 24948
rect 17714 24892 17724 24948
rect 17780 24892 20860 24948
rect 20916 24892 20926 24948
rect 24434 24892 24444 24948
rect 24500 24892 25340 24948
rect 25396 24892 26236 24948
rect 26292 24892 27132 24948
rect 27188 24892 27198 24948
rect 27356 24836 27412 25116
rect 39676 25060 39732 25116
rect 31266 25004 31276 25060
rect 31332 25004 39732 25060
rect 39890 25004 39900 25060
rect 39956 25004 40908 25060
rect 40964 25004 40974 25060
rect 6290 24780 6300 24836
rect 6356 24780 7644 24836
rect 7700 24780 7710 24836
rect 17490 24780 17500 24836
rect 17556 24780 26684 24836
rect 26740 24780 27412 24836
rect 27468 24892 35868 24948
rect 35924 24892 35934 24948
rect 27468 24724 27524 24892
rect 4610 24668 4620 24724
rect 4676 24668 4956 24724
rect 5012 24668 5022 24724
rect 5394 24668 5404 24724
rect 5460 24668 6076 24724
rect 6132 24668 6142 24724
rect 16594 24668 16604 24724
rect 16660 24668 17388 24724
rect 17444 24668 17454 24724
rect 20132 24668 22316 24724
rect 22372 24668 25900 24724
rect 25956 24668 27524 24724
rect 27580 24668 35364 24724
rect 35522 24668 35532 24724
rect 35588 24668 38780 24724
rect 38836 24668 40236 24724
rect 40292 24668 40302 24724
rect 20132 24612 20188 24668
rect 27580 24612 27636 24668
rect 35308 24612 35364 24668
rect 13234 24556 13244 24612
rect 13300 24556 20188 24612
rect 22082 24556 22092 24612
rect 22148 24556 22428 24612
rect 22484 24556 23996 24612
rect 24052 24556 24062 24612
rect 27570 24556 27580 24612
rect 27636 24556 27646 24612
rect 31490 24556 31500 24612
rect 31556 24556 34524 24612
rect 34580 24556 34590 24612
rect 35308 24556 40348 24612
rect 40404 24556 40908 24612
rect 40964 24556 40974 24612
rect 8306 24444 8316 24500
rect 8372 24444 10220 24500
rect 10276 24444 10286 24500
rect 24658 24444 24668 24500
rect 24724 24444 34972 24500
rect 35028 24444 35038 24500
rect 41458 24444 41468 24500
rect 41524 24444 41916 24500
rect 41972 24444 43708 24500
rect 43764 24444 43774 24500
rect 20850 24332 20860 24388
rect 20916 24332 21532 24388
rect 21588 24332 21598 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 8082 24220 8092 24276
rect 8148 24220 10668 24276
rect 10724 24220 17948 24276
rect 18004 24220 19516 24276
rect 19572 24220 19582 24276
rect 7746 24108 7756 24164
rect 7812 24108 21476 24164
rect 21420 24052 21476 24108
rect 20132 23996 21196 24052
rect 21252 23996 21262 24052
rect 21420 23996 25508 24052
rect 31266 23996 31276 24052
rect 31332 23996 32060 24052
rect 32116 23996 32126 24052
rect 40898 23996 40908 24052
rect 40964 23996 41692 24052
rect 41748 23996 41758 24052
rect 20132 23940 20188 23996
rect 25452 23940 25508 23996
rect 18274 23884 18284 23940
rect 18340 23884 20188 23940
rect 21522 23884 21532 23940
rect 21588 23884 22540 23940
rect 22596 23884 22606 23940
rect 25442 23884 25452 23940
rect 25508 23884 30156 23940
rect 30212 23884 30222 23940
rect 6066 23772 6076 23828
rect 6132 23772 7084 23828
rect 7140 23772 7150 23828
rect 16818 23772 16828 23828
rect 16884 23772 18732 23828
rect 18788 23772 18798 23828
rect 21858 23772 21868 23828
rect 21924 23772 22652 23828
rect 22708 23772 22718 23828
rect 2594 23660 2604 23716
rect 2660 23660 3724 23716
rect 3780 23660 3790 23716
rect 6290 23660 6300 23716
rect 6356 23660 6366 23716
rect 6300 23604 6356 23660
rect 3154 23548 3164 23604
rect 3220 23548 6356 23604
rect 8754 23548 8764 23604
rect 8820 23548 9996 23604
rect 10052 23548 10062 23604
rect 16818 23548 16828 23604
rect 16884 23548 17724 23604
rect 17780 23548 18284 23604
rect 18340 23548 18350 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 6514 23436 6524 23492
rect 6580 23436 7980 23492
rect 8036 23436 8046 23492
rect 9090 23212 9100 23268
rect 9156 23212 9548 23268
rect 9604 23212 14364 23268
rect 14420 23212 14430 23268
rect 14578 23212 14588 23268
rect 14644 23212 15260 23268
rect 15316 23212 15326 23268
rect 20178 22988 20188 23044
rect 20244 22988 21196 23044
rect 21252 22988 34860 23044
rect 34916 22988 35420 23044
rect 35476 22988 35486 23044
rect 16258 22876 16268 22932
rect 16324 22876 18620 22932
rect 18676 22876 18686 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 9986 22428 9996 22484
rect 10052 22428 16492 22484
rect 16548 22428 18508 22484
rect 18564 22428 18574 22484
rect 4722 22316 4732 22372
rect 4788 22316 5292 22372
rect 5348 22316 7084 22372
rect 7140 22316 7150 22372
rect 7634 22316 7644 22372
rect 7700 22316 8652 22372
rect 8708 22316 8718 22372
rect 1922 22204 1932 22260
rect 1988 22204 5516 22260
rect 5572 22204 5582 22260
rect 26786 22204 26796 22260
rect 26852 22204 28588 22260
rect 28644 22204 28654 22260
rect 2258 22092 2268 22148
rect 2324 22092 21532 22148
rect 21588 22092 21598 22148
rect 39442 22092 39452 22148
rect 39508 22092 40460 22148
rect 40516 22092 40908 22148
rect 40964 22092 40974 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 8306 21644 8316 21700
rect 8372 21644 13692 21700
rect 13748 21644 13758 21700
rect 6738 21532 6748 21588
rect 6804 21532 7420 21588
rect 7476 21532 7486 21588
rect 11442 21532 11452 21588
rect 11508 21532 12124 21588
rect 12180 21532 12190 21588
rect 5394 21420 5404 21476
rect 5460 21420 6412 21476
rect 6468 21420 11788 21476
rect 11844 21420 11854 21476
rect 15362 21308 15372 21364
rect 15428 21308 16268 21364
rect 16324 21308 16334 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 16594 20748 16604 20804
rect 16660 20748 17388 20804
rect 17444 20748 17454 20804
rect 37538 20748 37548 20804
rect 37604 20748 38780 20804
rect 38836 20748 38846 20804
rect 7410 20636 7420 20692
rect 7476 20636 11340 20692
rect 11396 20636 11406 20692
rect 15250 20636 15260 20692
rect 15316 20636 16716 20692
rect 16772 20636 16782 20692
rect 12562 20524 12572 20580
rect 12628 20524 15148 20580
rect 15092 20468 15148 20524
rect 16716 20524 20076 20580
rect 20132 20524 20142 20580
rect 16716 20468 16772 20524
rect 12674 20412 12684 20468
rect 12740 20412 14252 20468
rect 14308 20412 14588 20468
rect 14644 20412 14654 20468
rect 15092 20412 16716 20468
rect 16772 20412 16782 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 36082 20300 36092 20356
rect 36148 20300 38892 20356
rect 38948 20300 38958 20356
rect 10770 20188 10780 20244
rect 10836 20188 12236 20244
rect 12292 20188 12302 20244
rect 23090 20188 23100 20244
rect 23156 20188 23548 20244
rect 23604 20188 25788 20244
rect 25844 20188 25854 20244
rect 7746 20076 7756 20132
rect 7812 20076 9436 20132
rect 9492 20076 9502 20132
rect 9986 20076 9996 20132
rect 10052 20076 12348 20132
rect 12404 20076 12414 20132
rect 35186 20076 35196 20132
rect 35252 20076 35644 20132
rect 35700 20076 37548 20132
rect 37604 20076 37614 20132
rect 10546 19964 10556 20020
rect 10612 19964 12908 20020
rect 12964 19964 12974 20020
rect 25778 19964 25788 20020
rect 25844 19964 27132 20020
rect 27188 19964 27198 20020
rect 30034 19964 30044 20020
rect 30100 19964 30380 20020
rect 30436 19964 31388 20020
rect 31444 19964 31454 20020
rect 35074 19964 35084 20020
rect 35140 19964 35980 20020
rect 36036 19964 39004 20020
rect 39060 19964 39070 20020
rect 28690 19852 28700 19908
rect 28756 19852 29932 19908
rect 29988 19852 29998 19908
rect 10098 19740 10108 19796
rect 10164 19740 10892 19796
rect 10948 19740 10958 19796
rect 22866 19740 22876 19796
rect 22932 19740 23660 19796
rect 23716 19740 23726 19796
rect 26674 19740 26684 19796
rect 26740 19740 29260 19796
rect 29316 19740 29326 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 27122 19292 27132 19348
rect 27188 19292 29260 19348
rect 29316 19292 29326 19348
rect 29922 19180 29932 19236
rect 29988 19180 32060 19236
rect 32116 19180 32126 19236
rect 37986 19180 37996 19236
rect 38052 19180 38668 19236
rect 38724 19180 38734 19236
rect 17266 19068 17276 19124
rect 17332 19068 27244 19124
rect 27300 19068 27310 19124
rect 31892 19068 32172 19124
rect 32228 19068 32238 19124
rect 11890 18956 11900 19012
rect 11956 18956 16268 19012
rect 16324 18956 16334 19012
rect 30146 18956 30156 19012
rect 30212 18956 31164 19012
rect 31220 18956 31230 19012
rect 31892 18900 31948 19068
rect 9426 18844 9436 18900
rect 9492 18844 12124 18900
rect 12180 18844 12190 18900
rect 29474 18844 29484 18900
rect 29540 18844 31388 18900
rect 31444 18844 31948 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 9650 18732 9660 18788
rect 9716 18732 13804 18788
rect 13860 18732 15148 18788
rect 15092 18564 15148 18732
rect 8194 18508 8204 18564
rect 8260 18508 10444 18564
rect 10500 18508 10510 18564
rect 15092 18508 15708 18564
rect 15764 18508 16156 18564
rect 16212 18508 16222 18564
rect 9874 18396 9884 18452
rect 9940 18396 14700 18452
rect 14756 18396 15148 18452
rect 15362 18396 15372 18452
rect 15428 18396 17276 18452
rect 17332 18396 17342 18452
rect 21634 18396 21644 18452
rect 21700 18396 22092 18452
rect 22148 18396 22988 18452
rect 23044 18396 23054 18452
rect 15092 18340 15148 18396
rect 6962 18284 6972 18340
rect 7028 18284 10108 18340
rect 10164 18284 10174 18340
rect 15092 18284 16156 18340
rect 16212 18284 18732 18340
rect 18788 18284 18798 18340
rect 19506 18284 19516 18340
rect 19572 18284 20860 18340
rect 20916 18284 20926 18340
rect 32386 18284 32396 18340
rect 32452 18284 33180 18340
rect 33236 18284 35756 18340
rect 35812 18284 35822 18340
rect 14130 18172 14140 18228
rect 14196 18172 16492 18228
rect 16548 18172 21868 18228
rect 21924 18172 21934 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 39554 17724 39564 17780
rect 39620 17724 39900 17780
rect 39956 17724 40908 17780
rect 40964 17724 40974 17780
rect 41570 17724 41580 17780
rect 41636 17724 43820 17780
rect 43876 17724 43886 17780
rect 37538 17612 37548 17668
rect 37604 17612 39676 17668
rect 39732 17612 39742 17668
rect 8978 17500 8988 17556
rect 9044 17500 10108 17556
rect 10164 17500 10174 17556
rect 10658 17500 10668 17556
rect 10724 17500 11452 17556
rect 11508 17500 11518 17556
rect 17714 17500 17724 17556
rect 17780 17500 19404 17556
rect 19460 17500 19470 17556
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 32946 17164 32956 17220
rect 33012 17164 36428 17220
rect 36484 17164 37100 17220
rect 37156 17164 37166 17220
rect 10322 17052 10332 17108
rect 10388 17052 11340 17108
rect 11396 17052 11406 17108
rect 29362 17052 29372 17108
rect 29428 17052 33180 17108
rect 33236 17052 33246 17108
rect 40226 17052 40236 17108
rect 40292 17052 41468 17108
rect 41524 17052 41534 17108
rect 4386 16940 4396 16996
rect 4452 16940 9100 16996
rect 9156 16940 9166 16996
rect 11890 16940 11900 16996
rect 11956 16940 13804 16996
rect 13860 16940 13870 16996
rect 16930 16940 16940 16996
rect 16996 16940 17388 16996
rect 17444 16940 17454 16996
rect 17602 16940 17612 16996
rect 17668 16940 17948 16996
rect 18004 16940 32956 16996
rect 33012 16940 33022 16996
rect 39666 16940 39676 16996
rect 39732 16940 40124 16996
rect 40180 16940 41244 16996
rect 41300 16940 41310 16996
rect 1922 16828 1932 16884
rect 1988 16828 3612 16884
rect 3668 16828 3678 16884
rect 4834 16828 4844 16884
rect 4900 16828 9548 16884
rect 9604 16828 10220 16884
rect 10276 16828 10286 16884
rect 13346 16828 13356 16884
rect 13412 16828 14028 16884
rect 14084 16828 16156 16884
rect 16212 16828 17836 16884
rect 17892 16828 17902 16884
rect 20290 16828 20300 16884
rect 20356 16828 26012 16884
rect 26068 16828 26078 16884
rect 34850 16828 34860 16884
rect 34916 16828 35756 16884
rect 35812 16828 38108 16884
rect 38164 16828 38174 16884
rect 24220 16772 24276 16828
rect 6514 16716 6524 16772
rect 6580 16716 8988 16772
rect 9044 16716 9054 16772
rect 9874 16716 9884 16772
rect 9940 16716 13132 16772
rect 13188 16716 13198 16772
rect 24210 16716 24220 16772
rect 24276 16716 24286 16772
rect 11442 16604 11452 16660
rect 11508 16604 12348 16660
rect 12404 16604 12414 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 10994 16380 11004 16436
rect 11060 16380 11070 16436
rect 11004 16324 11060 16380
rect 3332 16268 11060 16324
rect 3332 16212 3388 16268
rect 2594 16156 2604 16212
rect 2660 16156 3388 16212
rect 5730 16156 5740 16212
rect 5796 16156 6972 16212
rect 7028 16156 7038 16212
rect 8978 16156 8988 16212
rect 9044 16156 12124 16212
rect 12180 16156 13020 16212
rect 13076 16156 13086 16212
rect 17266 16156 17276 16212
rect 17332 16156 19292 16212
rect 19348 16156 19358 16212
rect 29250 16156 29260 16212
rect 29316 16156 31948 16212
rect 32004 16156 32732 16212
rect 32788 16156 32798 16212
rect 9762 16044 9772 16100
rect 9828 16044 10220 16100
rect 10276 16044 11116 16100
rect 11172 16044 11676 16100
rect 11732 16044 11742 16100
rect 12450 16044 12460 16100
rect 12516 16044 13132 16100
rect 13188 16044 13198 16100
rect 24210 16044 24220 16100
rect 24276 16044 25732 16100
rect 25676 15988 25732 16044
rect 12226 15932 12236 15988
rect 12292 15932 12302 15988
rect 12786 15932 12796 15988
rect 12852 15932 20860 15988
rect 20916 15932 20926 15988
rect 22418 15932 22428 15988
rect 22484 15932 23324 15988
rect 23380 15932 24556 15988
rect 24612 15932 24622 15988
rect 24882 15932 24892 15988
rect 24948 15932 25452 15988
rect 25508 15932 25518 15988
rect 25666 15932 25676 15988
rect 25732 15932 25742 15988
rect 12236 15876 12292 15932
rect 9762 15820 9772 15876
rect 9828 15820 14588 15876
rect 14644 15820 14654 15876
rect 19282 15820 19292 15876
rect 19348 15820 28700 15876
rect 28756 15820 29372 15876
rect 29428 15820 29438 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 16146 15484 16156 15540
rect 16212 15484 18060 15540
rect 18116 15484 18126 15540
rect 19506 15484 19516 15540
rect 19572 15484 22820 15540
rect 16594 15372 16604 15428
rect 16660 15372 17388 15428
rect 17444 15372 17454 15428
rect 18834 15372 18844 15428
rect 18900 15372 19964 15428
rect 20020 15372 21084 15428
rect 21140 15372 21532 15428
rect 21588 15372 21868 15428
rect 21924 15372 21934 15428
rect 22764 15316 22820 15484
rect 23100 15484 23548 15540
rect 23604 15484 24108 15540
rect 24164 15484 24444 15540
rect 24500 15484 26012 15540
rect 26068 15484 26078 15540
rect 23100 15316 23156 15484
rect 25330 15372 25340 15428
rect 25396 15372 28028 15428
rect 28084 15372 28094 15428
rect 17714 15260 17724 15316
rect 17780 15260 18620 15316
rect 18676 15260 18686 15316
rect 22754 15260 22764 15316
rect 22820 15260 22830 15316
rect 23090 15260 23100 15316
rect 23156 15260 23166 15316
rect 23314 15260 23324 15316
rect 23380 15260 24220 15316
rect 24276 15260 24286 15316
rect 22764 15204 22820 15260
rect 15250 15148 15260 15204
rect 15316 15148 17612 15204
rect 17668 15148 17678 15204
rect 18050 15148 18060 15204
rect 18116 15148 20412 15204
rect 20468 15148 20478 15204
rect 21858 15148 21868 15204
rect 21924 15148 23436 15204
rect 23492 15148 23502 15204
rect 23986 15148 23996 15204
rect 24052 15148 24444 15204
rect 24500 15148 25900 15204
rect 25956 15148 25966 15204
rect 32498 15148 32508 15204
rect 32564 15148 33404 15204
rect 33460 15148 33470 15204
rect 19292 15092 19348 15148
rect 20412 15092 20468 15148
rect 19282 15036 19292 15092
rect 19348 15036 19358 15092
rect 20412 15036 24780 15092
rect 24836 15036 24846 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 31826 14812 31836 14868
rect 31892 14812 33068 14868
rect 33124 14812 33134 14868
rect 16258 14700 16268 14756
rect 16324 14700 16716 14756
rect 16772 14700 16782 14756
rect 16482 14588 16492 14644
rect 16548 14588 17612 14644
rect 17668 14588 18060 14644
rect 18116 14588 18126 14644
rect 14914 14476 14924 14532
rect 14980 14476 15484 14532
rect 15540 14476 15932 14532
rect 15988 14476 15998 14532
rect 17154 14476 17164 14532
rect 17220 14476 18172 14532
rect 18228 14476 18844 14532
rect 18900 14476 18910 14532
rect 36418 14476 36428 14532
rect 36484 14476 37660 14532
rect 37716 14476 37726 14532
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 10098 13916 10108 13972
rect 10164 13916 10556 13972
rect 10612 13916 10622 13972
rect 11330 13916 11340 13972
rect 11396 13916 14812 13972
rect 14868 13916 15596 13972
rect 15652 13916 16940 13972
rect 16996 13916 17006 13972
rect 35746 13916 35756 13972
rect 35812 13916 36764 13972
rect 36820 13916 36830 13972
rect 39890 13916 39900 13972
rect 39956 13916 41020 13972
rect 41076 13916 41086 13972
rect 35858 13804 35868 13860
rect 35924 13804 37436 13860
rect 37492 13804 37996 13860
rect 38052 13804 38062 13860
rect 23314 13692 23324 13748
rect 23380 13692 24220 13748
rect 24276 13692 24286 13748
rect 31602 13692 31612 13748
rect 31668 13692 32396 13748
rect 32452 13692 35756 13748
rect 35812 13692 35822 13748
rect 36530 13692 36540 13748
rect 36596 13692 37324 13748
rect 37380 13692 37390 13748
rect 4162 13580 4172 13636
rect 4228 13580 9660 13636
rect 9716 13580 9726 13636
rect 36194 13580 36204 13636
rect 36260 13580 37212 13636
rect 37268 13580 37278 13636
rect 40338 13580 40348 13636
rect 40404 13580 41356 13636
rect 41412 13580 43932 13636
rect 43988 13580 43998 13636
rect 9202 13468 9212 13524
rect 9268 13468 9996 13524
rect 10052 13468 10062 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 8642 13244 8652 13300
rect 8708 13244 9996 13300
rect 10052 13244 10062 13300
rect 8082 13132 8092 13188
rect 8148 13132 9660 13188
rect 9716 13132 9726 13188
rect 10434 13132 10444 13188
rect 10500 13132 11116 13188
rect 11172 13132 11182 13188
rect 9762 13020 9772 13076
rect 9828 13020 9838 13076
rect 38434 13020 38444 13076
rect 38500 13020 40124 13076
rect 40180 13020 40190 13076
rect 9772 12852 9828 13020
rect 10098 12908 10108 12964
rect 10164 12908 10444 12964
rect 10500 12908 10510 12964
rect 21410 12908 21420 12964
rect 21476 12908 21980 12964
rect 22036 12908 22046 12964
rect 37650 12908 37660 12964
rect 37716 12908 41020 12964
rect 41076 12908 41086 12964
rect 8866 12796 8876 12852
rect 8932 12796 11452 12852
rect 11508 12796 11518 12852
rect 21746 12796 21756 12852
rect 21812 12796 21822 12852
rect 7970 12684 7980 12740
rect 8036 12684 8316 12740
rect 8372 12684 9100 12740
rect 9156 12684 9166 12740
rect 11106 12684 11116 12740
rect 11172 12684 17164 12740
rect 17220 12684 17230 12740
rect 11116 12628 11172 12684
rect 9202 12572 9212 12628
rect 9268 12572 10556 12628
rect 10612 12572 11172 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 6402 12348 6412 12404
rect 6468 12348 7980 12404
rect 8036 12348 8046 12404
rect 4834 12236 4844 12292
rect 4900 12236 10780 12292
rect 10836 12236 11116 12292
rect 11172 12236 11182 12292
rect 21756 12180 21812 12796
rect 21980 12740 22036 12908
rect 21980 12684 22092 12740
rect 22148 12684 22158 12740
rect 40226 12348 40236 12404
rect 40292 12348 41020 12404
rect 41076 12348 41086 12404
rect 9090 12124 9100 12180
rect 9156 12124 9548 12180
rect 9604 12124 9614 12180
rect 21634 12124 21644 12180
rect 21700 12124 22204 12180
rect 22260 12124 22270 12180
rect 37538 12012 37548 12068
rect 37604 12012 38444 12068
rect 38500 12012 38510 12068
rect 1922 11900 1932 11956
rect 1988 11900 3500 11956
rect 3556 11900 5740 11956
rect 5796 11900 5806 11956
rect 21858 11900 21868 11956
rect 21924 11900 22428 11956
rect 22484 11900 22494 11956
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 9986 11676 9996 11732
rect 10052 11676 11228 11732
rect 11284 11676 11294 11732
rect 31602 11564 31612 11620
rect 31668 11564 31948 11620
rect 32004 11564 32014 11620
rect 5730 11452 5740 11508
rect 5796 11452 6972 11508
rect 7028 11452 7038 11508
rect 31826 11452 31836 11508
rect 31892 11452 32396 11508
rect 32452 11452 33012 11508
rect 36418 11452 36428 11508
rect 36484 11452 37660 11508
rect 37716 11452 37726 11508
rect 32956 11396 33012 11452
rect 2594 11340 2604 11396
rect 2660 11340 10220 11396
rect 10276 11340 10286 11396
rect 24546 11340 24556 11396
rect 24612 11340 25452 11396
rect 25508 11340 25518 11396
rect 31602 11340 31612 11396
rect 31668 11340 32060 11396
rect 32116 11340 32732 11396
rect 32788 11340 32798 11396
rect 32946 11340 32956 11396
rect 33012 11340 34636 11396
rect 34692 11340 34702 11396
rect 36194 11340 36204 11396
rect 36260 11340 37548 11396
rect 37604 11340 37614 11396
rect 12114 11228 12124 11284
rect 12180 11228 12684 11284
rect 12740 11228 12750 11284
rect 25106 11228 25116 11284
rect 25172 11228 26348 11284
rect 26404 11228 26414 11284
rect 8372 11116 8876 11172
rect 8932 11116 9996 11172
rect 10052 11116 10062 11172
rect 11778 11116 11788 11172
rect 11844 11116 12908 11172
rect 12964 11116 12974 11172
rect 32610 11116 32620 11172
rect 32676 11116 34524 11172
rect 34580 11116 36988 11172
rect 37044 11116 37054 11172
rect 8372 10612 8428 11116
rect 31266 11004 31276 11060
rect 31332 11004 31724 11060
rect 31780 11004 34188 11060
rect 34244 11004 35756 11060
rect 35812 11004 35822 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 24444 10892 25004 10948
rect 25060 10892 25070 10948
rect 24444 10836 24500 10892
rect 10210 10780 10220 10836
rect 10276 10780 10668 10836
rect 10724 10780 15372 10836
rect 15428 10780 16268 10836
rect 16324 10780 16334 10836
rect 17714 10780 17724 10836
rect 17780 10780 24444 10836
rect 24500 10780 24510 10836
rect 24658 10780 24668 10836
rect 24724 10780 25564 10836
rect 25620 10780 26124 10836
rect 26180 10780 26684 10836
rect 26740 10780 26750 10836
rect 29698 10780 29708 10836
rect 29764 10780 32508 10836
rect 32564 10780 33180 10836
rect 33236 10780 33246 10836
rect 35074 10780 35084 10836
rect 35140 10780 35532 10836
rect 35588 10780 36316 10836
rect 36372 10780 36382 10836
rect 12674 10668 12684 10724
rect 12740 10668 13580 10724
rect 13636 10668 13646 10724
rect 13906 10668 13916 10724
rect 13972 10668 20356 10724
rect 24210 10668 24220 10724
rect 24276 10668 25340 10724
rect 25396 10668 26012 10724
rect 26068 10668 26078 10724
rect 27010 10668 27020 10724
rect 27076 10668 28588 10724
rect 28644 10668 28654 10724
rect 20300 10612 20356 10668
rect 7858 10556 7868 10612
rect 7924 10556 7934 10612
rect 8194 10556 8204 10612
rect 8260 10556 8428 10612
rect 12898 10556 12908 10612
rect 12964 10556 18284 10612
rect 18340 10556 18350 10612
rect 20290 10556 20300 10612
rect 20356 10556 20366 10612
rect 7868 10500 7924 10556
rect 7868 10444 8876 10500
rect 8932 10444 14364 10500
rect 14420 10444 15260 10500
rect 15316 10444 15326 10500
rect 6962 10332 6972 10388
rect 7028 10332 8764 10388
rect 8820 10332 8830 10388
rect 12898 10332 12908 10388
rect 12964 10332 13692 10388
rect 13748 10332 13758 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 17826 9996 17836 10052
rect 17892 9996 19292 10052
rect 19348 9996 19358 10052
rect 19618 9996 19628 10052
rect 19684 9996 20412 10052
rect 20468 9996 20860 10052
rect 20916 9996 20926 10052
rect 24882 9884 24892 9940
rect 24948 9884 26460 9940
rect 26516 9884 26526 9940
rect 12450 9772 12460 9828
rect 12516 9772 13580 9828
rect 13636 9772 13646 9828
rect 13906 9772 13916 9828
rect 13972 9772 15036 9828
rect 15092 9772 15102 9828
rect 15362 9772 15372 9828
rect 15428 9772 15484 9828
rect 15540 9772 15550 9828
rect 15698 9772 15708 9828
rect 15764 9772 15820 9828
rect 15876 9772 15886 9828
rect 17378 9772 17388 9828
rect 17444 9772 17948 9828
rect 18004 9772 19068 9828
rect 19124 9772 19852 9828
rect 19908 9772 19918 9828
rect 25778 9772 25788 9828
rect 25844 9772 29260 9828
rect 29316 9772 29326 9828
rect 15036 9716 15092 9772
rect 15036 9660 15372 9716
rect 15428 9660 15438 9716
rect 15586 9660 15596 9716
rect 15652 9660 15662 9716
rect 15596 9604 15652 9660
rect 7746 9548 7756 9604
rect 7812 9548 8540 9604
rect 8596 9548 8606 9604
rect 14802 9548 14812 9604
rect 14868 9548 15708 9604
rect 15764 9548 16492 9604
rect 16548 9548 17948 9604
rect 18004 9548 18014 9604
rect 24658 9548 24668 9604
rect 24724 9548 25900 9604
rect 25956 9548 25966 9604
rect 31378 9548 31388 9604
rect 31444 9548 37100 9604
rect 37156 9548 37166 9604
rect 9762 9436 9772 9492
rect 9828 9436 12796 9492
rect 12852 9436 15820 9492
rect 15876 9436 15886 9492
rect 16706 9436 16716 9492
rect 16772 9436 18620 9492
rect 18676 9436 18686 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 15138 9324 15148 9380
rect 15204 9324 15708 9380
rect 15764 9324 15774 9380
rect 12338 9212 12348 9268
rect 12404 9212 12908 9268
rect 12964 9212 12974 9268
rect 15586 9212 15596 9268
rect 15652 9212 17612 9268
rect 17668 9212 17678 9268
rect 20066 9212 20076 9268
rect 20132 9212 21084 9268
rect 21140 9212 23996 9268
rect 24052 9212 24062 9268
rect 13570 9100 13580 9156
rect 13636 9100 14700 9156
rect 14756 9100 24388 9156
rect 24546 9100 24556 9156
rect 24612 9100 26124 9156
rect 26180 9100 26190 9156
rect 26562 9100 26572 9156
rect 26628 9100 28140 9156
rect 28196 9100 28206 9156
rect 24332 9044 24388 9100
rect 15670 8988 15708 9044
rect 15764 8988 15774 9044
rect 16706 8988 16716 9044
rect 16772 8988 17836 9044
rect 17892 8988 17902 9044
rect 24332 8988 25004 9044
rect 25060 8988 25676 9044
rect 25732 8988 30940 9044
rect 30996 8988 31006 9044
rect 35074 8988 35084 9044
rect 35140 8988 38332 9044
rect 38388 8988 38398 9044
rect 24658 8876 24668 8932
rect 24724 8876 25452 8932
rect 25508 8876 25518 8932
rect 15698 8764 15708 8820
rect 15764 8764 16268 8820
rect 16324 8764 16334 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 5618 8316 5628 8372
rect 5684 8316 7532 8372
rect 7588 8316 7598 8372
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 9650 7532 9660 7588
rect 9716 7532 12572 7588
rect 12628 7532 12638 7588
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 12562 6412 12572 6468
rect 12628 6412 13580 6468
rect 13636 6412 13646 6468
rect 21746 6412 21756 6468
rect 21812 6412 23436 6468
rect 23492 6412 23502 6468
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 16370 5516 16380 5572
rect 16436 5516 18956 5572
rect 19012 5516 19022 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 13570 5068 13580 5124
rect 13636 5068 15372 5124
rect 15428 5068 15438 5124
rect 16146 5068 16156 5124
rect 16212 5068 16828 5124
rect 16884 5068 16894 5124
rect 24098 5068 24108 5124
rect 24164 5068 24780 5124
rect 24836 5068 24846 5124
rect 20402 4956 20412 5012
rect 20468 4956 22204 5012
rect 22260 4956 22270 5012
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 16818 4508 16828 4564
rect 16884 4508 18732 4564
rect 18788 4508 19180 4564
rect 19236 4508 19246 4564
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 15372 10780 15428 10836
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 15372 9772 15428 9828
rect 15820 9772 15876 9828
rect 15708 9548 15764 9604
rect 15820 9436 15876 9492
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 15708 8988 15764 9044
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 42396
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 19808 42364 20128 42396
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 15372 10836 15428 10846
rect 15372 9828 15428 10780
rect 15372 9762 15428 9772
rect 15820 9828 15876 9838
rect 15708 9604 15764 9614
rect 15708 9044 15764 9548
rect 15820 9492 15876 9772
rect 15820 9426 15876 9436
rect 19808 9436 20128 10948
rect 15708 8978 15764 8988
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 41580 35488 42396
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _342_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8624 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _343_
timestamp 1698431365
transform -1 0 29680 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _344_
timestamp 1698431365
transform -1 0 32368 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _345_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27664 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _346_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24528 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _347_
timestamp 1698431365
transform -1 0 28224 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _348_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25424 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _349_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25536 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _350_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31584 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _351_
timestamp 1698431365
transform -1 0 20832 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _352_
timestamp 1698431365
transform -1 0 18256 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _353_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10080 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _354_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _355_
timestamp 1698431365
transform -1 0 15568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _356_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14672 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _357_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16352 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _358_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7280 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _359_
timestamp 1698431365
transform 1 0 6160 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _360_
timestamp 1698431365
transform 1 0 6832 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _361_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31920 0 1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _362_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38528 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _363_
timestamp 1698431365
transform 1 0 37408 0 1 14112
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _364_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35616 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _365_
timestamp 1698431365
transform 1 0 10416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _366_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _367_
timestamp 1698431365
transform 1 0 18368 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _368_
timestamp 1698431365
transform 1 0 26096 0 -1 14112
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _369_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9744 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _370_
timestamp 1698431365
transform -1 0 9184 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _371_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _372_
timestamp 1698431365
transform -1 0 17360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _373_
timestamp 1698431365
transform 1 0 6608 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _374_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11984 0 1 18816
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _375_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _376_
timestamp 1698431365
transform 1 0 7840 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _377_
timestamp 1698431365
transform -1 0 16912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _378_
timestamp 1698431365
transform 1 0 12096 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _379_
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _380_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11088 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _381_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15680 0 -1 20384
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _382_
timestamp 1698431365
transform -1 0 9296 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _383_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _384_
timestamp 1698431365
transform -1 0 15120 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _385_
timestamp 1698431365
transform 1 0 9968 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _386_
timestamp 1698431365
transform -1 0 11984 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _387_
timestamp 1698431365
transform 1 0 10416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _388_
timestamp 1698431365
transform -1 0 12880 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _389_
timestamp 1698431365
transform 1 0 11984 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _390_
timestamp 1698431365
transform 1 0 15232 0 1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _391_
timestamp 1698431365
transform 1 0 15008 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _392_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _393_
timestamp 1698431365
transform -1 0 24864 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _394_
timestamp 1698431365
transform -1 0 18928 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _395_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17584 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _396_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15344 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _397_
timestamp 1698431365
transform 1 0 14000 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _398_
timestamp 1698431365
transform -1 0 15120 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _399_
timestamp 1698431365
transform -1 0 7392 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _400_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18368 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _401_
timestamp 1698431365
transform -1 0 18256 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _402_
timestamp 1698431365
transform -1 0 19376 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _403_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17696 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _404_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16688 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _405_
timestamp 1698431365
transform -1 0 17920 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _406_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16912 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _407_
timestamp 1698431365
transform -1 0 11088 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _408_
timestamp 1698431365
transform -1 0 11648 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _409_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10080 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _410_
timestamp 1698431365
transform -1 0 15792 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _411_
timestamp 1698431365
transform -1 0 15344 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _412_
timestamp 1698431365
transform -1 0 10192 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _413_
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _414_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _415_
timestamp 1698431365
transform -1 0 8176 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _416_
timestamp 1698431365
transform -1 0 7952 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _417_
timestamp 1698431365
transform 1 0 6160 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _418_
timestamp 1698431365
transform 1 0 10304 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _419_
timestamp 1698431365
transform -1 0 10528 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _420_
timestamp 1698431365
transform 1 0 6944 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _421_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9632 0 1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _422_
timestamp 1698431365
transform 1 0 10080 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _423_
timestamp 1698431365
transform -1 0 11648 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _424_
timestamp 1698431365
transform -1 0 9184 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _425_
timestamp 1698431365
transform -1 0 10304 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _426_
timestamp 1698431365
transform -1 0 9408 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _427_
timestamp 1698431365
transform 1 0 11648 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _428_
timestamp 1698431365
transform 1 0 7504 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _429_
timestamp 1698431365
transform 1 0 9968 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _430_
timestamp 1698431365
transform 1 0 7952 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _431_
timestamp 1698431365
transform 1 0 11424 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _432_
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _433_
timestamp 1698431365
transform 1 0 11200 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _434_
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _435_
timestamp 1698431365
transform 1 0 37072 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _436_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _437_
timestamp 1698431365
transform 1 0 38528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _438_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37744 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _439_
timestamp 1698431365
transform 1 0 41104 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _440_
timestamp 1698431365
transform 1 0 23968 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _441_
timestamp 1698431365
transform 1 0 26992 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _442_
timestamp 1698431365
transform 1 0 39984 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _443_
timestamp 1698431365
transform 1 0 40208 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _444_
timestamp 1698431365
transform 1 0 41328 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _445_
timestamp 1698431365
transform -1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _446_
timestamp 1698431365
transform -1 0 41328 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _447_
timestamp 1698431365
transform -1 0 15792 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _448_
timestamp 1698431365
transform -1 0 40656 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _449_
timestamp 1698431365
transform -1 0 38640 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _450_
timestamp 1698431365
transform -1 0 37968 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _451_
timestamp 1698431365
transform 1 0 40656 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _452_
timestamp 1698431365
transform 1 0 41552 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _453_
timestamp 1698431365
transform -1 0 36624 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _454_
timestamp 1698431365
transform 1 0 26096 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _455_
timestamp 1698431365
transform -1 0 37632 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _456_
timestamp 1698431365
transform 1 0 35840 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _457_
timestamp 1698431365
transform -1 0 37968 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _458_
timestamp 1698431365
transform -1 0 34720 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _459_
timestamp 1698431365
transform 1 0 35728 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _460_
timestamp 1698431365
transform -1 0 36176 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _461_
timestamp 1698431365
transform -1 0 33600 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _462_
timestamp 1698431365
transform 1 0 31696 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _463_
timestamp 1698431365
transform 1 0 31248 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _464_
timestamp 1698431365
transform 1 0 31136 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _465_
timestamp 1698431365
transform -1 0 33152 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _466_
timestamp 1698431365
transform -1 0 32032 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _467_
timestamp 1698431365
transform -1 0 32144 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _468_
timestamp 1698431365
transform -1 0 26208 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _469_
timestamp 1698431365
transform -1 0 31808 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _470_
timestamp 1698431365
transform -1 0 30912 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _471_
timestamp 1698431365
transform -1 0 23744 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _472_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30464 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _473_
timestamp 1698431365
transform -1 0 26880 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _474_
timestamp 1698431365
transform -1 0 35168 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _475_
timestamp 1698431365
transform -1 0 26768 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _476_
timestamp 1698431365
transform 1 0 31808 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _477_
timestamp 1698431365
transform 1 0 32480 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _478_
timestamp 1698431365
transform 1 0 37632 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _479_
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _480_
timestamp 1698431365
transform 1 0 35504 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _481_
timestamp 1698431365
transform -1 0 37744 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _482_
timestamp 1698431365
transform 1 0 35616 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _483_
timestamp 1698431365
transform -1 0 23968 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _484_
timestamp 1698431365
transform 1 0 25536 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _485_
timestamp 1698431365
transform 1 0 29792 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _486_
timestamp 1698431365
transform -1 0 31920 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _487_
timestamp 1698431365
transform 1 0 34496 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _488_
timestamp 1698431365
transform -1 0 31360 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _489_
timestamp 1698431365
transform 1 0 30576 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _490_
timestamp 1698431365
transform 1 0 35840 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _491_
timestamp 1698431365
transform -1 0 38304 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _492_
timestamp 1698431365
transform 1 0 36624 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _493_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _494_
timestamp 1698431365
transform 1 0 31248 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _495_
timestamp 1698431365
transform 1 0 32144 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _496_
timestamp 1698431365
transform -1 0 32144 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _497_
timestamp 1698431365
transform 1 0 24640 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _498_
timestamp 1698431365
transform -1 0 32144 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _499_
timestamp 1698431365
transform 1 0 30464 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _500_
timestamp 1698431365
transform -1 0 31136 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _501_
timestamp 1698431365
transform -1 0 31472 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _502_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _503_
timestamp 1698431365
transform 1 0 40656 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _504_
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _505_
timestamp 1698431365
transform 1 0 31248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _506_
timestamp 1698431365
transform -1 0 31024 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _507_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31472 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _508_
timestamp 1698431365
transform -1 0 33040 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _509_
timestamp 1698431365
transform -1 0 29568 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _510_
timestamp 1698431365
transform 1 0 29568 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _511_
timestamp 1698431365
transform -1 0 39648 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _512_
timestamp 1698431365
transform -1 0 35504 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _513_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _514_
timestamp 1698431365
transform -1 0 42000 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _515_
timestamp 1698431365
transform 1 0 39872 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _516_
timestamp 1698431365
transform 1 0 39872 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _517_
timestamp 1698431365
transform 1 0 41104 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _518_
timestamp 1698431365
transform -1 0 42672 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _519_
timestamp 1698431365
transform 1 0 41440 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _520_
timestamp 1698431365
transform 1 0 41328 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _521_
timestamp 1698431365
transform -1 0 42448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _522_
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _523_
timestamp 1698431365
transform -1 0 26768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _524_
timestamp 1698431365
transform -1 0 42112 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _525_
timestamp 1698431365
transform 1 0 41552 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _526_
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _527_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _528_
timestamp 1698431365
transform 1 0 41104 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _529_
timestamp 1698431365
transform -1 0 42000 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _530_
timestamp 1698431365
transform -1 0 38976 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _531_
timestamp 1698431365
transform -1 0 38080 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _532_
timestamp 1698431365
transform 1 0 25200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _533_
timestamp 1698431365
transform -1 0 37184 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _534_
timestamp 1698431365
transform -1 0 36624 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _535_
timestamp 1698431365
transform 1 0 34944 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _536_
timestamp 1698431365
transform 1 0 40320 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _537_
timestamp 1698431365
transform 1 0 39872 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _538_
timestamp 1698431365
transform 1 0 41440 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _539_
timestamp 1698431365
transform 1 0 40880 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _540_
timestamp 1698431365
transform -1 0 42896 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _541_
timestamp 1698431365
transform -1 0 42336 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _542_
timestamp 1698431365
transform 1 0 16016 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _543_
timestamp 1698431365
transform 1 0 18256 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _544_
timestamp 1698431365
transform 1 0 16128 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _545_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _546_
timestamp 1698431365
transform 1 0 23744 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _547_
timestamp 1698431365
transform -1 0 18144 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _548_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19712 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _549_
timestamp 1698431365
transform 1 0 16128 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _550_
timestamp 1698431365
transform 1 0 16128 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _551_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _552_
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _553_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22288 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _554_
timestamp 1698431365
transform -1 0 16352 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _555_
timestamp 1698431365
transform 1 0 18368 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _556_
timestamp 1698431365
transform 1 0 19824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _557_
timestamp 1698431365
transform -1 0 18368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _558_
timestamp 1698431365
transform -1 0 16688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _559_
timestamp 1698431365
transform -1 0 15792 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _560_
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _561_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _562_
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _563_
timestamp 1698431365
transform -1 0 14336 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _564_
timestamp 1698431365
transform -1 0 21392 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _565_
timestamp 1698431365
transform -1 0 15120 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _566_
timestamp 1698431365
transform -1 0 13776 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _567_
timestamp 1698431365
transform 1 0 11872 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _568_
timestamp 1698431365
transform 1 0 11200 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _569_
timestamp 1698431365
transform -1 0 12096 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _570_
timestamp 1698431365
transform -1 0 17920 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _571_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10416 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _572_
timestamp 1698431365
transform 1 0 8512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _573_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _574_
timestamp 1698431365
transform 1 0 8848 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _575_
timestamp 1698431365
transform -1 0 8848 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _576_
timestamp 1698431365
transform 1 0 8512 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _577_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _578_
timestamp 1698431365
transform 1 0 7392 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _579_
timestamp 1698431365
transform -1 0 9072 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _580_
timestamp 1698431365
transform 1 0 8624 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _581_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _582_
timestamp 1698431365
transform -1 0 8624 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _583_
timestamp 1698431365
transform 1 0 8288 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _584_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _585_
timestamp 1698431365
transform 1 0 11648 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _586_
timestamp 1698431365
transform -1 0 11872 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _587_
timestamp 1698431365
transform 1 0 9744 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _588_
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _589_
timestamp 1698431365
transform -1 0 12768 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _590_
timestamp 1698431365
transform 1 0 11984 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _591_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11872 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _592_
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _593_
timestamp 1698431365
transform 1 0 13440 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _594_
timestamp 1698431365
transform 1 0 15456 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _595_
timestamp 1698431365
transform -1 0 16240 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _596_
timestamp 1698431365
transform -1 0 15232 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _597_
timestamp 1698431365
transform 1 0 14672 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _598_
timestamp 1698431365
transform -1 0 18592 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _599_
timestamp 1698431365
transform -1 0 17696 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _600_
timestamp 1698431365
transform 1 0 17584 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _601_
timestamp 1698431365
transform -1 0 17920 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _602_
timestamp 1698431365
transform 1 0 16464 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _603_
timestamp 1698431365
transform -1 0 20720 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _604_
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _605_
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _606_
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _607_
timestamp 1698431365
transform -1 0 21840 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _608_
timestamp 1698431365
transform 1 0 19936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _609_
timestamp 1698431365
transform 1 0 19152 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _610_
timestamp 1698431365
transform 1 0 22064 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _611_
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _612_
timestamp 1698431365
transform 1 0 21392 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _613_
timestamp 1698431365
transform -1 0 22288 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _614_
timestamp 1698431365
transform -1 0 22064 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _615_
timestamp 1698431365
transform 1 0 21504 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _616_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _617_
timestamp 1698431365
transform -1 0 26544 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _618_
timestamp 1698431365
transform -1 0 23520 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _619_
timestamp 1698431365
transform 1 0 21728 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _620_
timestamp 1698431365
transform -1 0 23744 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _621_
timestamp 1698431365
transform -1 0 23408 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _622_
timestamp 1698431365
transform 1 0 24416 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _623_
timestamp 1698431365
transform 1 0 23408 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _624_
timestamp 1698431365
transform 1 0 23856 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _625_
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _626_
timestamp 1698431365
transform -1 0 27216 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _627_
timestamp 1698431365
transform 1 0 25312 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _628_
timestamp 1698431365
transform 1 0 23744 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _629_
timestamp 1698431365
transform 1 0 25872 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _630_
timestamp 1698431365
transform -1 0 25312 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _631_
timestamp 1698431365
transform 1 0 25200 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _632_
timestamp 1698431365
transform 1 0 24640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _633_
timestamp 1698431365
transform -1 0 26768 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _634_
timestamp 1698431365
transform 1 0 24080 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _635_
timestamp 1698431365
transform 1 0 24192 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _636_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _637_
timestamp 1698431365
transform 1 0 14672 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _638_
timestamp 1698431365
transform -1 0 16688 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _639_
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _640_
timestamp 1698431365
transform -1 0 16016 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _641_
timestamp 1698431365
transform -1 0 15792 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _642_
timestamp 1698431365
transform -1 0 17584 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _643_
timestamp 1698431365
transform -1 0 23408 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _644_
timestamp 1698431365
transform -1 0 22064 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _645_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _646_
timestamp 1698431365
transform 1 0 12768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _647_
timestamp 1698431365
transform -1 0 12880 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _648_
timestamp 1698431365
transform -1 0 12992 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _649_
timestamp 1698431365
transform -1 0 12432 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _650_
timestamp 1698431365
transform -1 0 12096 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _651_
timestamp 1698431365
transform 1 0 10416 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _652_
timestamp 1698431365
transform 1 0 10752 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _653_
timestamp 1698431365
transform 1 0 10976 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _654_
timestamp 1698431365
transform -1 0 16240 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _655_
timestamp 1698431365
transform -1 0 11424 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _656_
timestamp 1698431365
transform 1 0 7168 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _657_
timestamp 1698431365
transform -1 0 6384 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _658_
timestamp 1698431365
transform 1 0 6944 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _659_
timestamp 1698431365
transform 1 0 6048 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _660_
timestamp 1698431365
transform -1 0 5488 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _661_
timestamp 1698431365
transform -1 0 5600 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _662_
timestamp 1698431365
transform -1 0 5040 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _663_
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _664_
timestamp 1698431365
transform -1 0 4480 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _665_
timestamp 1698431365
transform -1 0 5040 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _666_
timestamp 1698431365
transform 1 0 5040 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _667_
timestamp 1698431365
transform 1 0 5712 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _668_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _669_
timestamp 1698431365
transform -1 0 4480 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _670_
timestamp 1698431365
transform -1 0 5936 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _671_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _672_
timestamp 1698431365
transform -1 0 5264 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _673_
timestamp 1698431365
transform -1 0 26096 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _674_
timestamp 1698431365
transform -1 0 22064 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _675_
timestamp 1698431365
transform -1 0 27440 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _676_
timestamp 1698431365
transform 1 0 26208 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _677_
timestamp 1698431365
transform 1 0 26544 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _678_
timestamp 1698431365
transform 1 0 27440 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _679_
timestamp 1698431365
transform -1 0 24416 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _680_
timestamp 1698431365
transform -1 0 22064 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _681_
timestamp 1698431365
transform 1 0 23856 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _682_
timestamp 1698431365
transform 1 0 25984 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _683_
timestamp 1698431365
transform -1 0 25984 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _684_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _685_
timestamp 1698431365
transform 1 0 2800 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _686_
timestamp 1698431365
transform 1 0 10528 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _687_
timestamp 1698431365
transform 1 0 20160 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _688_
timestamp 1698431365
transform 1 0 28336 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _689_
timestamp 1698431365
transform 1 0 33264 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _690_
timestamp 1698431365
transform 1 0 13776 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _691_
timestamp 1698431365
transform 1 0 35952 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _692_
timestamp 1698431365
transform 1 0 35616 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _693_
timestamp 1698431365
transform 1 0 40768 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _694_
timestamp 1698431365
transform 1 0 40880 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _695_
timestamp 1698431365
transform 1 0 34608 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _696_
timestamp 1698431365
transform 1 0 34832 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _697_
timestamp 1698431365
transform 1 0 29456 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _698_
timestamp 1698431365
transform 1 0 29456 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _699_
timestamp 1698431365
transform -1 0 32592 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _700_
timestamp 1698431365
transform 1 0 25648 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _701_
timestamp 1698431365
transform 1 0 1680 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _702_
timestamp 1698431365
transform 1 0 1680 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _703_
timestamp 1698431365
transform 1 0 4032 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _704_
timestamp 1698431365
transform 1 0 34384 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _705_
timestamp 1698431365
transform 1 0 30016 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _706_
timestamp 1698431365
transform -1 0 38640 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _707_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31248 0 1 39200
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _708_
timestamp 1698431365
transform 1 0 28560 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _709_
timestamp 1698431365
transform -1 0 35504 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _710_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _711_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _712_
timestamp 1698431365
transform -1 0 37968 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _713_
timestamp 1698431365
transform 1 0 40544 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _714_
timestamp 1698431365
transform 1 0 40880 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _715_
timestamp 1698431365
transform 1 0 40768 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _716_
timestamp 1698431365
transform 1 0 40656 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _717_
timestamp 1698431365
transform 1 0 35280 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _718_
timestamp 1698431365
transform -1 0 41440 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _719_
timestamp 1698431365
transform 1 0 40992 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _720_
timestamp 1698431365
transform -1 0 23184 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _721_
timestamp 1698431365
transform -1 0 21840 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _722_
timestamp 1698431365
transform 1 0 1680 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _723_
timestamp 1698431365
transform 1 0 3472 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _724_
timestamp 1698431365
transform 1 0 3248 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _725_
timestamp 1698431365
transform -1 0 8736 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _726_
timestamp 1698431365
transform 1 0 1680 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _727_
timestamp 1698431365
transform -1 0 12768 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _728_
timestamp 1698431365
transform 1 0 13328 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _729_
timestamp 1698431365
transform 1 0 15568 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _730_
timestamp 1698431365
transform 1 0 18928 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _731_
timestamp 1698431365
transform -1 0 24416 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _732_
timestamp 1698431365
transform 1 0 22736 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _733_
timestamp 1698431365
transform -1 0 29008 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _734_
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _735_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _736_
timestamp 1698431365
transform -1 0 19264 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _737_
timestamp 1698431365
transform -1 0 22848 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _738_
timestamp 1698431365
transform -1 0 12656 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _739_
timestamp 1698431365
transform 1 0 5936 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _740_
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _741_
timestamp 1698431365
transform 1 0 1680 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _742_
timestamp 1698431365
transform 1 0 2016 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _743_
timestamp 1698431365
transform 1 0 1680 0 -1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _744_
timestamp 1698431365
transform 1 0 19936 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _745_
timestamp 1698431365
transform 1 0 27328 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _746_
timestamp 1698431365
transform 1 0 19824 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _747_
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__B
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A1
timestamp 1698431365
transform 1 0 14112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A1
timestamp 1698431365
transform 1 0 11424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A2
timestamp 1698431365
transform -1 0 12432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A1
timestamp 1698431365
transform -1 0 10528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A1
timestamp 1698431365
transform 1 0 10192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A2
timestamp 1698431365
transform 1 0 10080 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A1
timestamp 1698431365
transform -1 0 12208 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__I
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__I
timestamp 1698431365
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__A1
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__I
timestamp 1698431365
transform 1 0 23072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__A1
timestamp 1698431365
transform 1 0 39984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__I
timestamp 1698431365
transform -1 0 14896 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__A1
timestamp 1698431365
transform 1 0 37072 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__B
timestamp 1698431365
transform -1 0 35840 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__A1
timestamp 1698431365
transform 1 0 35056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__B
timestamp 1698431365
transform -1 0 31696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A1
timestamp 1698431365
transform 1 0 30912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__B
timestamp 1698431365
transform 1 0 30016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__I
timestamp 1698431365
transform -1 0 23072 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__A1
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__I
timestamp 1698431365
transform 1 0 35392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__I
timestamp 1698431365
transform 1 0 26992 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__I
timestamp 1698431365
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__I
timestamp 1698431365
transform 1 0 22624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__I
timestamp 1698431365
transform 1 0 30688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A1
timestamp 1698431365
transform 1 0 30128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__I
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__B
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__A1
timestamp 1698431365
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__I
timestamp 1698431365
transform 1 0 39648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__C
timestamp 1698431365
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__I
timestamp 1698431365
transform 1 0 26992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__A2
timestamp 1698431365
transform 1 0 41328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__C
timestamp 1698431365
transform 1 0 40880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__C
timestamp 1698431365
transform 1 0 35840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__I
timestamp 1698431365
transform 1 0 34720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__A2
timestamp 1698431365
transform -1 0 40320 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A2
timestamp 1698431365
transform 1 0 39648 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__A2
timestamp 1698431365
transform -1 0 39872 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__A2
timestamp 1698431365
transform 1 0 43120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__I
timestamp 1698431365
transform 1 0 18032 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A1
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__A1
timestamp 1698431365
transform -1 0 18032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__B
timestamp 1698431365
transform 1 0 19936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__549__A2
timestamp 1698431365
transform 1 0 15904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__553__B
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__I
timestamp 1698431365
transform 1 0 17024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__A2
timestamp 1698431365
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__561__A2
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__A1
timestamp 1698431365
transform 1 0 20160 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__A2
timestamp 1698431365
transform 1 0 12880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__I
timestamp 1698431365
transform 1 0 10976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__A2
timestamp 1698431365
transform 1 0 10640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__B
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__A2
timestamp 1698431365
transform 1 0 12992 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__C
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__A2
timestamp 1698431365
transform 1 0 16240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__B
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__C
timestamp 1698431365
transform 1 0 17584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__I
timestamp 1698431365
transform 1 0 18816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__A2
timestamp 1698431365
transform 1 0 21056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__609__C
timestamp 1698431365
transform -1 0 19152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__614__C
timestamp 1698431365
transform -1 0 22288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__616__I
timestamp 1698431365
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__621__A1
timestamp 1698431365
transform -1 0 22736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__625__B
timestamp 1698431365
transform 1 0 24192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__A2
timestamp 1698431365
transform 1 0 24528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__635__A2
timestamp 1698431365
transform 1 0 23968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__636__C
timestamp 1698431365
transform -1 0 25088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__639__B
timestamp 1698431365
transform 1 0 17472 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__644__B
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__A1
timestamp 1698431365
transform 1 0 13104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__652__B2
timestamp 1698431365
transform -1 0 12208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__653__A1
timestamp 1698431365
transform 1 0 11872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__658__A1
timestamp 1698431365
transform 1 0 7728 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__663__A1
timestamp 1698431365
transform 1 0 5824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__664__A1
timestamp 1698431365
transform -1 0 3696 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__668__C
timestamp 1698431365
transform -1 0 7056 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__671__A3
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__672__A1
timestamp 1698431365
transform -1 0 5600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__A2
timestamp 1698431365
transform 1 0 26320 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__A1
timestamp 1698431365
transform -1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__A2
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__676__A3
timestamp 1698431365
transform -1 0 27216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__677__A1
timestamp 1698431365
transform -1 0 27552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__680__A1
timestamp 1698431365
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__A1
timestamp 1698431365
transform 1 0 27104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__B
timestamp 1698431365
transform 1 0 27552 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__684__CLK
timestamp 1698431365
transform 1 0 17024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__685__CLK
timestamp 1698431365
transform 1 0 6272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__CLK
timestamp 1698431365
transform -1 0 14000 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__687__CLK
timestamp 1698431365
transform -1 0 20160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__688__CLK
timestamp 1698431365
transform 1 0 31808 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__688__D
timestamp 1698431365
transform -1 0 28336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__CLK
timestamp 1698431365
transform -1 0 36960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__D
timestamp 1698431365
transform -1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__690__CLK
timestamp 1698431365
transform -1 0 17696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__691__CLK
timestamp 1698431365
transform 1 0 39424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__692__CLK
timestamp 1698431365
transform 1 0 39088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__693__CLK
timestamp 1698431365
transform 1 0 39536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__694__CLK
timestamp 1698431365
transform 1 0 39872 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__695__CLK
timestamp 1698431365
transform 1 0 38080 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__696__CLK
timestamp 1698431365
transform 1 0 38304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__697__CLK
timestamp 1698431365
transform 1 0 32704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__699__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__700__CLK
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__702__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__703__CLK
timestamp 1698431365
transform 1 0 7504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__704__CLK
timestamp 1698431365
transform 1 0 37632 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__705__CLK
timestamp 1698431365
transform 1 0 33488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__706__CLK
timestamp 1698431365
transform 1 0 38864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__CLK
timestamp 1698431365
transform 1 0 34944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__CLK
timestamp 1698431365
transform 1 0 32032 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__CLK
timestamp 1698431365
transform -1 0 35952 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__CLK
timestamp 1698431365
transform -1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__CLK
timestamp 1698431365
transform 1 0 38192 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__CLK
timestamp 1698431365
transform 1 0 40320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__714__CLK
timestamp 1698431365
transform 1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__715__CLK
timestamp 1698431365
transform 1 0 40544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__CLK
timestamp 1698431365
transform 1 0 40432 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__717__CLK
timestamp 1698431365
transform 1 0 38752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__718__CLK
timestamp 1698431365
transform 1 0 37968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__719__CLK
timestamp 1698431365
transform 1 0 39200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__720__CLK
timestamp 1698431365
transform -1 0 23632 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__721__CLK
timestamp 1698431365
transform 1 0 22064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__722__CLK
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__723__CLK
timestamp 1698431365
transform 1 0 6944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__724__CLK
timestamp 1698431365
transform 1 0 6944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__725__CLK
timestamp 1698431365
transform -1 0 9184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__726__CLK
timestamp 1698431365
transform 1 0 5712 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__727__CLK
timestamp 1698431365
transform 1 0 13552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__728__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__729__CLK
timestamp 1698431365
transform 1 0 15344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__730__CLK
timestamp 1698431365
transform 1 0 18704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__731__CLK
timestamp 1698431365
transform -1 0 24864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__CLK
timestamp 1698431365
transform 1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__733__CLK
timestamp 1698431365
transform 1 0 29232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__CLK
timestamp 1698431365
transform 1 0 29232 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__735__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__736__CLK
timestamp 1698431365
transform -1 0 19712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__CLK
timestamp 1698431365
transform 1 0 23632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__738__CLK
timestamp 1698431365
transform -1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__739__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__740__CLK
timestamp 1698431365
transform 1 0 5936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__741__CLK
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__742__CLK
timestamp 1698431365
transform 1 0 5712 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__743__CLK
timestamp 1698431365
transform 1 0 5824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__744__CLK
timestamp 1698431365
transform 1 0 19712 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__745__CLK
timestamp 1698431365
transform 1 0 30800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__746__CLK
timestamp 1698431365
transform 1 0 19600 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__747__CLK
timestamp 1698431365
transform -1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 21616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 15344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 19376 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 17920 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 20160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output10_I
timestamp 1698431365
transform 1 0 39760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 15120 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1698431365
transform -1 0 16128 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1698431365
transform -1 0 20160 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1698431365
transform 1 0 33376 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1698431365
transform 1 0 33264 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_376 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_104 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_106 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13216 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_154
timestamp 1698431365
transform 1 0 18592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_186 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22176 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_202
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_123
timestamp 1698431365
transform 1 0 15120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_156
timestamp 1698431365
transform 1 0 18816 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_172
timestamp 1698431365
transform 1 0 20608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_206
timestamp 1698431365
transform 1 0 24416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_210
timestamp 1698431365
transform 1 0 24864 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_383
timestamp 1698431365
transform 1 0 44240 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_189
timestamp 1698431365
transform 1 0 22512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_205
timestamp 1698431365
transform 1 0 24304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_241
timestamp 1698431365
transform 1 0 28336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_245
timestamp 1698431365
transform 1 0 28784 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_277
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_102
timestamp 1698431365
transform 1 0 12768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_111
timestamp 1698431365
transform 1 0 13776 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_143
timestamp 1698431365
transform 1 0 17360 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_147
timestamp 1698431365
transform 1 0 17808 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_154
timestamp 1698431365
transform 1 0 18592 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_170
timestamp 1698431365
transform 1 0 20384 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_179
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_184
timestamp 1698431365
transform 1 0 21952 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_216
timestamp 1698431365
transform 1 0 25536 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_232
timestamp 1698431365
transform 1 0 27328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_240
timestamp 1698431365
transform 1 0 28224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_383
timestamp 1698431365
transform 1 0 44240 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_66
timestamp 1698431365
transform 1 0 8736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_70
timestamp 1698431365
transform 1 0 9184 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_102
timestamp 1698431365
transform 1 0 12768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_212
timestamp 1698431365
transform 1 0 25088 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_88
timestamp 1698431365
transform 1 0 11200 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_92
timestamp 1698431365
transform 1 0 11648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_94
timestamp 1698431365
transform 1 0 11872 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_103
timestamp 1698431365
transform 1 0 12880 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_125
timestamp 1698431365
transform 1 0 15344 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_131
timestamp 1698431365
transform 1 0 16016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_133
timestamp 1698431365
transform 1 0 16240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_151
timestamp 1698431365
transform 1 0 18256 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_159
timestamp 1698431365
transform 1 0 19152 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_163
timestamp 1698431365
transform 1 0 19600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_165
timestamp 1698431365
transform 1 0 19824 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_174
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_178
timestamp 1698431365
transform 1 0 21280 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_194
timestamp 1698431365
transform 1 0 23072 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_227
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_259
timestamp 1698431365
transform 1 0 30352 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_275
timestamp 1698431365
transform 1 0 32144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_298
timestamp 1698431365
transform 1 0 34720 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_328
timestamp 1698431365
transform 1 0 38080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_332
timestamp 1698431365
transform 1 0 38528 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_348
timestamp 1698431365
transform 1 0 40320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_68
timestamp 1698431365
transform 1 0 8960 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_84
timestamp 1698431365
transform 1 0 10752 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_92
timestamp 1698431365
transform 1 0 11648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_111
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_133
timestamp 1698431365
transform 1 0 16240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_152
timestamp 1698431365
transform 1 0 18368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_156
timestamp 1698431365
transform 1 0 18816 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_193
timestamp 1698431365
transform 1 0 22960 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_201
timestamp 1698431365
transform 1 0 23856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_205
timestamp 1698431365
transform 1 0 24304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_207
timestamp 1698431365
transform 1 0 24528 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_251
timestamp 1698431365
transform 1 0 29456 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_259
timestamp 1698431365
transform 1 0 30352 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_263
timestamp 1698431365
transform 1 0 30800 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_274
timestamp 1698431365
transform 1 0 32032 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_306
timestamp 1698431365
transform 1 0 35616 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_383
timestamp 1698431365
transform 1 0 44240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_50
timestamp 1698431365
transform 1 0 6944 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_54
timestamp 1698431365
transform 1 0 7392 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_56
timestamp 1698431365
transform 1 0 7616 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_65
timestamp 1698431365
transform 1 0 8624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_81
timestamp 1698431365
transform 1 0 10416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_85
timestamp 1698431365
transform 1 0 10864 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_93
timestamp 1698431365
transform 1 0 11760 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_102
timestamp 1698431365
transform 1 0 12768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_106
timestamp 1698431365
transform 1 0 13216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_114
timestamp 1698431365
transform 1 0 14112 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_122
timestamp 1698431365
transform 1 0 15008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_126
timestamp 1698431365
transform 1 0 15456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_130
timestamp 1698431365
transform 1 0 15904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_132
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_135
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_144
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_147
timestamp 1698431365
transform 1 0 17808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_149
timestamp 1698431365
transform 1 0 18032 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_187
timestamp 1698431365
transform 1 0 22288 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_221
timestamp 1698431365
transform 1 0 26096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_231
timestamp 1698431365
transform 1 0 27216 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_247
timestamp 1698431365
transform 1 0 29008 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_286
timestamp 1698431365
transform 1 0 33376 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_294
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_298
timestamp 1698431365
transform 1 0 34720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_300
timestamp 1698431365
transform 1 0 34944 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_311
timestamp 1698431365
transform 1 0 36176 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_343
timestamp 1698431365
transform 1 0 39760 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_347
timestamp 1698431365
transform 1 0 40208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_41
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_57
timestamp 1698431365
transform 1 0 7728 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_70
timestamp 1698431365
transform 1 0 9184 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_86
timestamp 1698431365
transform 1 0 10976 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_90
timestamp 1698431365
transform 1 0 11424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_98
timestamp 1698431365
transform 1 0 12320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1698431365
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_148
timestamp 1698431365
transform 1 0 17920 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_164
timestamp 1698431365
transform 1 0 19712 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_183
timestamp 1698431365
transform 1 0 21840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_187
timestamp 1698431365
transform 1 0 22288 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_203
timestamp 1698431365
transform 1 0 24080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_224
timestamp 1698431365
transform 1 0 26432 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_240
timestamp 1698431365
transform 1 0 28224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_263
timestamp 1698431365
transform 1 0 30800 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_265
timestamp 1698431365
transform 1 0 31024 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_284
timestamp 1698431365
transform 1 0 33152 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_298
timestamp 1698431365
transform 1 0 34720 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_306
timestamp 1698431365
transform 1 0 35616 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_327
timestamp 1698431365
transform 1 0 37968 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_359
timestamp 1698431365
transform 1 0 41552 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_375
timestamp 1698431365
transform 1 0 43344 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_383
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_14
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_16
timestamp 1698431365
transform 1 0 3136 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_48
timestamp 1698431365
transform 1 0 6720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_52
timestamp 1698431365
transform 1 0 7168 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_60
timestamp 1698431365
transform 1 0 8064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_62
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_112
timestamp 1698431365
transform 1 0 13888 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_128
timestamp 1698431365
transform 1 0 15680 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_174
timestamp 1698431365
transform 1 0 20832 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_193
timestamp 1698431365
transform 1 0 22960 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_314
timestamp 1698431365
transform 1 0 36512 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_318
timestamp 1698431365
transform 1 0 36960 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_333
timestamp 1698431365
transform 1 0 38640 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_357
timestamp 1698431365
transform 1 0 41328 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_373
timestamp 1698431365
transform 1 0 43120 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_381
timestamp 1698431365
transform 1 0 44016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_383
timestamp 1698431365
transform 1 0 44240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_53
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_57
timestamp 1698431365
transform 1 0 7728 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_73
timestamp 1698431365
transform 1 0 9520 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_94
timestamp 1698431365
transform 1 0 11872 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_197
timestamp 1698431365
transform 1 0 23408 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_229
timestamp 1698431365
transform 1 0 26992 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_333
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_341
timestamp 1698431365
transform 1 0 39536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_365
timestamp 1698431365
transform 1 0 42224 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_383
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_34
timestamp 1698431365
transform 1 0 5152 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_50
timestamp 1698431365
transform 1 0 6944 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_58
timestamp 1698431365
transform 1 0 7840 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_82
timestamp 1698431365
transform 1 0 10528 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_114
timestamp 1698431365
transform 1 0 14112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_118
timestamp 1698431365
transform 1 0 14560 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_129
timestamp 1698431365
transform 1 0 15792 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_174
timestamp 1698431365
transform 1 0 20832 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_178
timestamp 1698431365
transform 1 0 21280 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_184
timestamp 1698431365
transform 1 0 21952 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_258
timestamp 1698431365
transform 1 0 30240 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_266
timestamp 1698431365
transform 1 0 31136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_268
timestamp 1698431365
transform 1 0 31360 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_298
timestamp 1698431365
transform 1 0 34720 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_324
timestamp 1698431365
transform 1 0 37632 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_340
timestamp 1698431365
transform 1 0 39424 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_382
timestamp 1698431365
transform 1 0 44128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_53
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_61
timestamp 1698431365
transform 1 0 8176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_63
timestamp 1698431365
transform 1 0 8400 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_68
timestamp 1698431365
transform 1 0 8960 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_84
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_94
timestamp 1698431365
transform 1 0 11872 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_102
timestamp 1698431365
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_137
timestamp 1698431365
transform 1 0 16688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_152
timestamp 1698431365
transform 1 0 18368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_158
timestamp 1698431365
transform 1 0 19040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_162
timestamp 1698431365
transform 1 0 19488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_170
timestamp 1698431365
transform 1 0 20384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_193
timestamp 1698431365
transform 1 0 22960 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_203
timestamp 1698431365
transform 1 0 24080 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_235
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_263
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_275
timestamp 1698431365
transform 1 0 32144 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_279
timestamp 1698431365
transform 1 0 32592 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_282
timestamp 1698431365
transform 1 0 32928 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_298
timestamp 1698431365
transform 1 0 34720 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_306
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_308
timestamp 1698431365
transform 1 0 35840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_321
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_359
timestamp 1698431365
transform 1 0 41552 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_375
timestamp 1698431365
transform 1 0 43344 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_383
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_81
timestamp 1698431365
transform 1 0 10416 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_97
timestamp 1698431365
transform 1 0 12208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_101
timestamp 1698431365
transform 1 0 12656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_105
timestamp 1698431365
transform 1 0 13104 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_151
timestamp 1698431365
transform 1 0 18256 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_164
timestamp 1698431365
transform 1 0 19712 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_179
timestamp 1698431365
transform 1 0 21392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_181
timestamp 1698431365
transform 1 0 21616 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_198
timestamp 1698431365
transform 1 0 23520 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_200
timestamp 1698431365
transform 1 0 23744 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_247
timestamp 1698431365
transform 1 0 29008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_288
timestamp 1698431365
transform 1 0 33600 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_296
timestamp 1698431365
transform 1 0 34496 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_326
timestamp 1698431365
transform 1 0 37856 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698431365
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_41
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_57
timestamp 1698431365
transform 1 0 7728 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_65
timestamp 1698431365
transform 1 0 8624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_77
timestamp 1698431365
transform 1 0 9968 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_93
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_157
timestamp 1698431365
transform 1 0 18928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_161
timestamp 1698431365
transform 1 0 19376 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_169
timestamp 1698431365
transform 1 0 20272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698431365
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_189
timestamp 1698431365
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_200
timestamp 1698431365
transform 1 0 23744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_225
timestamp 1698431365
transform 1 0 26544 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_297
timestamp 1698431365
transform 1 0 34608 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_313
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_383
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_18
timestamp 1698431365
transform 1 0 3360 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_48
timestamp 1698431365
transform 1 0 6720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_52
timestamp 1698431365
transform 1 0 7168 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_82
timestamp 1698431365
transform 1 0 10528 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_96
timestamp 1698431365
transform 1 0 12096 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_116
timestamp 1698431365
transform 1 0 14336 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_124
timestamp 1698431365
transform 1 0 15232 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_150
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_182
timestamp 1698431365
transform 1 0 21728 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_198
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_336
timestamp 1698431365
transform 1 0 38976 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_344
timestamp 1698431365
transform 1 0 39872 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_354
timestamp 1698431365
transform 1 0 40992 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_361
timestamp 1698431365
transform 1 0 41776 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_377
timestamp 1698431365
transform 1 0 43568 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_381
timestamp 1698431365
transform 1 0 44016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_383
timestamp 1698431365
transform 1 0 44240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_61
timestamp 1698431365
transform 1 0 8176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_65
timestamp 1698431365
transform 1 0 8624 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_93
timestamp 1698431365
transform 1 0 11760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_95
timestamp 1698431365
transform 1 0 11984 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_100
timestamp 1698431365
transform 1 0 12544 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_123
timestamp 1698431365
transform 1 0 15120 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_127
timestamp 1698431365
transform 1 0 15568 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_134
timestamp 1698431365
transform 1 0 16352 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_138
timestamp 1698431365
transform 1 0 16800 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_142
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_158
timestamp 1698431365
transform 1 0 19040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_166
timestamp 1698431365
transform 1 0 19936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698431365
transform 1 0 20384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_343
timestamp 1698431365
transform 1 0 39760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_381
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_383
timestamp 1698431365
transform 1 0 44240 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_123
timestamp 1698431365
transform 1 0 15120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_127
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698431365
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_187
timestamp 1698431365
transform 1 0 22288 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698431365
transform 1 0 24080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_222
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_238
timestamp 1698431365
transform 1 0 28000 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_246
timestamp 1698431365
transform 1 0 28896 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_286
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_302
timestamp 1698431365
transform 1 0 35168 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_335
timestamp 1698431365
transform 1 0 38864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_339
timestamp 1698431365
transform 1 0 39312 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_347
timestamp 1698431365
transform 1 0 40208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_356
timestamp 1698431365
transform 1 0 41216 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_363
timestamp 1698431365
transform 1 0 42000 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_379
timestamp 1698431365
transform 1 0 43792 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_383
timestamp 1698431365
transform 1 0 44240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_53
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_95
timestamp 1698431365
transform 1 0 11984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_123
timestamp 1698431365
transform 1 0 15120 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_131
timestamp 1698431365
transform 1 0 16016 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_145
timestamp 1698431365
transform 1 0 17584 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_161
timestamp 1698431365
transform 1 0 19376 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_169
timestamp 1698431365
transform 1 0 20272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_185
timestamp 1698431365
transform 1 0 22064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_189
timestamp 1698431365
transform 1 0 22512 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_220
timestamp 1698431365
transform 1 0 25984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_228
timestamp 1698431365
transform 1 0 26880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_240
timestamp 1698431365
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_255
timestamp 1698431365
transform 1 0 29904 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_272
timestamp 1698431365
transform 1 0 31808 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_310
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_321
timestamp 1698431365
transform 1 0 37296 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_340
timestamp 1698431365
transform 1 0 39424 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_372
timestamp 1698431365
transform 1 0 43008 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_380
timestamp 1698431365
transform 1 0 43904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_39
timestamp 1698431365
transform 1 0 5712 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_43
timestamp 1698431365
transform 1 0 6160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_59
timestamp 1698431365
transform 1 0 7952 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_84
timestamp 1698431365
transform 1 0 10752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_128
timestamp 1698431365
transform 1 0 15680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_130
timestamp 1698431365
transform 1 0 15904 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_174
timestamp 1698431365
transform 1 0 20832 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_182
timestamp 1698431365
transform 1 0 21728 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_186
timestamp 1698431365
transform 1 0 22176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_188
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_197
timestamp 1698431365
transform 1 0 23408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698431365
transform 1 0 24304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_216
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_246
timestamp 1698431365
transform 1 0 28896 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_260
timestamp 1698431365
transform 1 0 30464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_264
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_266
timestamp 1698431365
transform 1 0 31136 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698431365
transform 1 0 32144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_311
timestamp 1698431365
transform 1 0 36176 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_343
timestamp 1698431365
transform 1 0 39760 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_53
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_103
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_161
timestamp 1698431365
transform 1 0 19376 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_169
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698431365
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_279
timestamp 1698431365
transform 1 0 32592 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_306
timestamp 1698431365
transform 1 0 35616 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_357
timestamp 1698431365
transform 1 0 41328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_373
timestamp 1698431365
transform 1 0 43120 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_381
timestamp 1698431365
transform 1 0 44016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_34
timestamp 1698431365
transform 1 0 5152 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_42
timestamp 1698431365
transform 1 0 6048 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_49
timestamp 1698431365
transform 1 0 6832 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_57
timestamp 1698431365
transform 1 0 7728 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_65
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_76
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_78
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_158
timestamp 1698431365
transform 1 0 19040 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_195
timestamp 1698431365
transform 1 0 23184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_199
timestamp 1698431365
transform 1 0 23632 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698431365
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_298
timestamp 1698431365
transform 1 0 34720 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_306
timestamp 1698431365
transform 1 0 35616 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_308
timestamp 1698431365
transform 1 0 35840 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_338
timestamp 1698431365
transform 1 0 39200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_342
timestamp 1698431365
transform 1 0 39648 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698431365
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_41
timestamp 1698431365
transform 1 0 5936 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_81
timestamp 1698431365
transform 1 0 10416 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_97
timestamp 1698431365
transform 1 0 12208 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_131
timestamp 1698431365
transform 1 0 16016 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_148
timestamp 1698431365
transform 1 0 17920 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_164
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_231
timestamp 1698431365
transform 1 0 27216 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_239
timestamp 1698431365
transform 1 0 28112 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_380
timestamp 1698431365
transform 1 0 43904 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_26
timestamp 1698431365
transform 1 0 4256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_30
timestamp 1698431365
transform 1 0 4704 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_37
timestamp 1698431365
transform 1 0 5488 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698431365
transform 1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_96
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_100
timestamp 1698431365
transform 1 0 12544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_134
timestamp 1698431365
transform 1 0 16352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_175
timestamp 1698431365
transform 1 0 20944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_179
timestamp 1698431365
transform 1 0 21392 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_195
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_244
timestamp 1698431365
transform 1 0 28672 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_260
timestamp 1698431365
transform 1 0 30464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_264
timestamp 1698431365
transform 1 0 30912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_269
timestamp 1698431365
transform 1 0 31472 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_275
timestamp 1698431365
transform 1 0 32144 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_294
timestamp 1698431365
transform 1 0 34272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_302
timestamp 1698431365
transform 1 0 35168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_306
timestamp 1698431365
transform 1 0 35616 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_338
timestamp 1698431365
transform 1 0 39200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_356
timestamp 1698431365
transform 1 0 41216 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_358
timestamp 1698431365
transform 1 0 41440 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_363
timestamp 1698431365
transform 1 0 42000 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_379
timestamp 1698431365
transform 1 0 43792 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_383
timestamp 1698431365
transform 1 0 44240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_55
timestamp 1698431365
transform 1 0 7504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_59
timestamp 1698431365
transform 1 0 7952 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_91
timestamp 1698431365
transform 1 0 11536 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_99
timestamp 1698431365
transform 1 0 12432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_103
timestamp 1698431365
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_139
timestamp 1698431365
transform 1 0 16912 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_164
timestamp 1698431365
transform 1 0 19712 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_195
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_211
timestamp 1698431365
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_213
timestamp 1698431365
transform 1 0 25200 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_222
timestamp 1698431365
transform 1 0 26208 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698431365
transform 1 0 28000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_305
timestamp 1698431365
transform 1 0 35504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_309
timestamp 1698431365
transform 1 0 35952 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_349
timestamp 1698431365
transform 1 0 40432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_365
timestamp 1698431365
transform 1 0 42224 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_381
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_383
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_18
timestamp 1698431365
transform 1 0 3360 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_26
timestamp 1698431365
transform 1 0 4256 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_38
timestamp 1698431365
transform 1 0 5600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_42
timestamp 1698431365
transform 1 0 6048 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_54
timestamp 1698431365
transform 1 0 7392 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_64
timestamp 1698431365
transform 1 0 8512 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_85
timestamp 1698431365
transform 1 0 10864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_89
timestamp 1698431365
transform 1 0 11312 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_121
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_129
timestamp 1698431365
transform 1 0 15792 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_150
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_182
timestamp 1698431365
transform 1 0 21728 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_198
timestamp 1698431365
transform 1 0 23520 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_237
timestamp 1698431365
transform 1 0 27888 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_253
timestamp 1698431365
transform 1 0 29680 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_261
timestamp 1698431365
transform 1 0 30576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_265
timestamp 1698431365
transform 1 0 31024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_275
timestamp 1698431365
transform 1 0 32144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_298
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_302
timestamp 1698431365
transform 1 0 35168 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_332
timestamp 1698431365
transform 1 0 38528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_336
timestamp 1698431365
transform 1 0 38976 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_344
timestamp 1698431365
transform 1 0 39872 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_348
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_357
timestamp 1698431365
transform 1 0 41328 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_373
timestamp 1698431365
transform 1 0 43120 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_381
timestamp 1698431365
transform 1 0 44016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_383
timestamp 1698431365
transform 1 0 44240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_51
timestamp 1698431365
transform 1 0 7056 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_66
timestamp 1698431365
transform 1 0 8736 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_82
timestamp 1698431365
transform 1 0 10528 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_90
timestamp 1698431365
transform 1 0 11424 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_98
timestamp 1698431365
transform 1 0 12320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_102
timestamp 1698431365
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_121
timestamp 1698431365
transform 1 0 14896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_125
timestamp 1698431365
transform 1 0 15344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_133
timestamp 1698431365
transform 1 0 16240 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_151
timestamp 1698431365
transform 1 0 18256 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_167
timestamp 1698431365
transform 1 0 20048 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_183
timestamp 1698431365
transform 1 0 21840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_187
timestamp 1698431365
transform 1 0 22288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_189
timestamp 1698431365
transform 1 0 22512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_192
timestamp 1698431365
transform 1 0 22848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_222
timestamp 1698431365
transform 1 0 26208 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_269
timestamp 1698431365
transform 1 0 31472 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_301
timestamp 1698431365
transform 1 0 35056 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_323
timestamp 1698431365
transform 1 0 37520 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_331
timestamp 1698431365
transform 1 0 38416 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_346
timestamp 1698431365
transform 1 0 40096 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_350
timestamp 1698431365
transform 1 0 40544 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_357
timestamp 1698431365
transform 1 0 41328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_373
timestamp 1698431365
transform 1 0 43120 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_383
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_18
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_22
timestamp 1698431365
transform 1 0 3808 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_43
timestamp 1698431365
transform 1 0 6160 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_59
timestamp 1698431365
transform 1 0 7952 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_78
timestamp 1698431365
transform 1 0 10080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_80
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_89
timestamp 1698431365
transform 1 0 11312 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_99
timestamp 1698431365
transform 1 0 12432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_101
timestamp 1698431365
transform 1 0 12656 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_110
timestamp 1698431365
transform 1 0 13664 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_118
timestamp 1698431365
transform 1 0 14560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_120
timestamp 1698431365
transform 1 0 14784 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_127
timestamp 1698431365
transform 1 0 15568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_131
timestamp 1698431365
transform 1 0 16016 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_148
timestamp 1698431365
transform 1 0 17920 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_150
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_157
timestamp 1698431365
transform 1 0 18928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_189
timestamp 1698431365
transform 1 0 22512 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_290
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_306
timestamp 1698431365
transform 1 0 35616 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_320
timestamp 1698431365
transform 1 0 37184 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_336
timestamp 1698431365
transform 1 0 38976 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_344
timestamp 1698431365
transform 1 0 39872 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_354
timestamp 1698431365
transform 1 0 40992 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_367
timestamp 1698431365
transform 1 0 42448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_383
timestamp 1698431365
transform 1 0 44240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_47
timestamp 1698431365
transform 1 0 6608 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_63
timestamp 1698431365
transform 1 0 8400 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_71
timestamp 1698431365
transform 1 0 9296 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_83
timestamp 1698431365
transform 1 0 10640 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_93
timestamp 1698431365
transform 1 0 11760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_97
timestamp 1698431365
transform 1 0 12208 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_131
timestamp 1698431365
transform 1 0 16016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_143
timestamp 1698431365
transform 1 0 17360 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_259
timestamp 1698431365
transform 1 0 30352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_265
timestamp 1698431365
transform 1 0 31024 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_269
timestamp 1698431365
transform 1 0 31472 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_275
timestamp 1698431365
transform 1 0 32144 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_307
timestamp 1698431365
transform 1 0 35728 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698431365
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_328
timestamp 1698431365
transform 1 0 38080 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_344
timestamp 1698431365
transform 1 0 39872 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_348
timestamp 1698431365
transform 1 0 40320 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_350
timestamp 1698431365
transform 1 0 40544 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_34
timestamp 1698431365
transform 1 0 5152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_41
timestamp 1698431365
transform 1 0 5936 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_57
timestamp 1698431365
transform 1 0 7728 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_65
timestamp 1698431365
transform 1 0 8624 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_88
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_96
timestamp 1698431365
transform 1 0 12096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_103
timestamp 1698431365
transform 1 0 12880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_107
timestamp 1698431365
transform 1 0 13328 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_158
timestamp 1698431365
transform 1 0 19040 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_162
timestamp 1698431365
transform 1 0 19488 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_197
timestamp 1698431365
transform 1 0 23408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_201
timestamp 1698431365
transform 1 0 23856 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_241
timestamp 1698431365
transform 1 0 28336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_245
timestamp 1698431365
transform 1 0 28784 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_253
timestamp 1698431365
transform 1 0 29680 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_259
timestamp 1698431365
transform 1 0 30352 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_275
timestamp 1698431365
transform 1 0 32144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_356
timestamp 1698431365
transform 1 0 41216 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_367
timestamp 1698431365
transform 1 0 42448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_383
timestamp 1698431365
transform 1 0 44240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_18
timestamp 1698431365
transform 1 0 3360 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_26
timestamp 1698431365
transform 1 0 4256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_47
timestamp 1698431365
transform 1 0 6608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_51
timestamp 1698431365
transform 1 0 7056 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_83
timestamp 1698431365
transform 1 0 10640 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_87
timestamp 1698431365
transform 1 0 11088 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_89
timestamp 1698431365
transform 1 0 11312 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_115
timestamp 1698431365
transform 1 0 14224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_119
timestamp 1698431365
transform 1 0 14672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_121
timestamp 1698431365
transform 1 0 14896 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_145
timestamp 1698431365
transform 1 0 17584 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_161
timestamp 1698431365
transform 1 0 19376 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_169
timestamp 1698431365
transform 1 0 20272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698431365
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_189
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_227
timestamp 1698431365
transform 1 0 26768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_231
timestamp 1698431365
transform 1 0 27216 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_239
timestamp 1698431365
transform 1 0 28112 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_266
timestamp 1698431365
transform 1 0 31136 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_270
timestamp 1698431365
transform 1 0 31584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_283
timestamp 1698431365
transform 1 0 33040 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_291
timestamp 1698431365
transform 1 0 33936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_295
timestamp 1698431365
transform 1 0 34384 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_302
timestamp 1698431365
transform 1 0 35168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_306
timestamp 1698431365
transform 1 0 35616 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_34
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_38
timestamp 1698431365
transform 1 0 5600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_42
timestamp 1698431365
transform 1 0 6048 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_58
timestamp 1698431365
transform 1 0 7840 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_80
timestamp 1698431365
transform 1 0 10304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_84
timestamp 1698431365
transform 1 0 10752 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_92
timestamp 1698431365
transform 1 0 11648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_96
timestamp 1698431365
transform 1 0 12096 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_104
timestamp 1698431365
transform 1 0 12992 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_108
timestamp 1698431365
transform 1 0 13440 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_110
timestamp 1698431365
transform 1 0 13664 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_119
timestamp 1698431365
transform 1 0 14672 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_135
timestamp 1698431365
transform 1 0 16464 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_174
timestamp 1698431365
transform 1 0 20832 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_190
timestamp 1698431365
transform 1 0 22624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_200
timestamp 1698431365
transform 1 0 23744 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_205
timestamp 1698431365
transform 1 0 24304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_228
timestamp 1698431365
transform 1 0 26880 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_236
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_240
timestamp 1698431365
transform 1 0 28224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_242
timestamp 1698431365
transform 1 0 28448 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_272
timestamp 1698431365
transform 1 0 31808 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_327
timestamp 1698431365
transform 1 0 37968 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_331
timestamp 1698431365
transform 1 0 38416 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_347
timestamp 1698431365
transform 1 0 40208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_356
timestamp 1698431365
transform 1 0 41216 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_363
timestamp 1698431365
transform 1 0 42000 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_379
timestamp 1698431365
transform 1 0 43792 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_383
timestamp 1698431365
transform 1 0 44240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_69
timestamp 1698431365
transform 1 0 9072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_71
timestamp 1698431365
transform 1 0 9296 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_160
timestamp 1698431365
transform 1 0 19264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_164
timestamp 1698431365
transform 1 0 19712 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698431365
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_297
timestamp 1698431365
transform 1 0 34608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_299
timestamp 1698431365
transform 1 0 34832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_333
timestamp 1698431365
transform 1 0 38640 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_342
timestamp 1698431365
transform 1 0 39648 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_346
timestamp 1698431365
transform 1 0 40096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_379
timestamp 1698431365
transform 1 0 43792 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_383
timestamp 1698431365
transform 1 0 44240 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_18
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_22
timestamp 1698431365
transform 1 0 3808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_28
timestamp 1698431365
transform 1 0 4480 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_36
timestamp 1698431365
transform 1 0 5376 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_40
timestamp 1698431365
transform 1 0 5824 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_76
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_80
timestamp 1698431365
transform 1 0 10304 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_146
timestamp 1698431365
transform 1 0 17696 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_166
timestamp 1698431365
transform 1 0 19936 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_170
timestamp 1698431365
transform 1 0 20384 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_202
timestamp 1698431365
transform 1 0 23968 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_244
timestamp 1698431365
transform 1 0 28672 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_265
timestamp 1698431365
transform 1 0 31024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_272
timestamp 1698431365
transform 1 0 31808 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_284
timestamp 1698431365
transform 1 0 33152 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_335
timestamp 1698431365
transform 1 0 38864 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_343
timestamp 1698431365
transform 1 0 39760 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_354
timestamp 1698431365
transform 1 0 40992 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_363
timestamp 1698431365
transform 1 0 42000 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_379
timestamp 1698431365
transform 1 0 43792 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_383
timestamp 1698431365
transform 1 0 44240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_41
timestamp 1698431365
transform 1 0 5936 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_73
timestamp 1698431365
transform 1 0 9520 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_89
timestamp 1698431365
transform 1 0 11312 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_97
timestamp 1698431365
transform 1 0 12208 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_115
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_117
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_168
timestamp 1698431365
transform 1 0 20160 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_172
timestamp 1698431365
transform 1 0 20608 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_185
timestamp 1698431365
transform 1 0 22064 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_201
timestamp 1698431365
transform 1 0 23856 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_209
timestamp 1698431365
transform 1 0 24752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_211
timestamp 1698431365
transform 1 0 24976 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_228
timestamp 1698431365
transform 1 0 26880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_232
timestamp 1698431365
transform 1 0 27328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_236
timestamp 1698431365
transform 1 0 27776 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_253
timestamp 1698431365
transform 1 0 29680 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_260
timestamp 1698431365
transform 1 0 30464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_264
timestamp 1698431365
transform 1 0 30912 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_296
timestamp 1698431365
transform 1 0 34496 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_323
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_339
timestamp 1698431365
transform 1 0 39312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_341
timestamp 1698431365
transform 1 0 39536 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_350
timestamp 1698431365
transform 1 0 40544 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_382
timestamp 1698431365
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_104
timestamp 1698431365
transform 1 0 12992 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_120
timestamp 1698431365
transform 1 0 14784 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_128
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_158
timestamp 1698431365
transform 1 0 19040 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_162
timestamp 1698431365
transform 1 0 19488 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_216
timestamp 1698431365
transform 1 0 25536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_218
timestamp 1698431365
transform 1 0 25760 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_227
timestamp 1698431365
transform 1 0 26768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_231
timestamp 1698431365
transform 1 0 27216 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_325
timestamp 1698431365
transform 1 0 37744 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_341
timestamp 1698431365
transform 1 0 39536 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_365
timestamp 1698431365
transform 1 0 42224 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_381
timestamp 1698431365
transform 1 0 44016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_383
timestamp 1698431365
transform 1 0 44240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_69
timestamp 1698431365
transform 1 0 9072 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_77
timestamp 1698431365
transform 1 0 9968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_81
timestamp 1698431365
transform 1 0 10416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_85
timestamp 1698431365
transform 1 0 10864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_87
timestamp 1698431365
transform 1 0 11088 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_94
timestamp 1698431365
transform 1 0 11872 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_102
timestamp 1698431365
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_216
timestamp 1698431365
transform 1 0 25536 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_224
timestamp 1698431365
transform 1 0 26432 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_230
timestamp 1698431365
transform 1 0 27104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_234
timestamp 1698431365
transform 1 0 27552 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_242
timestamp 1698431365
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_259
timestamp 1698431365
transform 1 0 30352 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_273
timestamp 1698431365
transform 1 0 31920 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_277
timestamp 1698431365
transform 1 0 32368 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_283
timestamp 1698431365
transform 1 0 33040 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_291
timestamp 1698431365
transform 1 0 33936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_295
timestamp 1698431365
transform 1 0 34384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_297
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_330
timestamp 1698431365
transform 1 0 38304 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_346
timestamp 1698431365
transform 1 0 40096 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_354
timestamp 1698431365
transform 1 0 40992 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_358
timestamp 1698431365
transform 1 0 41440 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_367
timestamp 1698431365
transform 1 0 42448 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_383
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_18
timestamp 1698431365
transform 1 0 3360 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_22
timestamp 1698431365
transform 1 0 3808 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_53
timestamp 1698431365
transform 1 0 7280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_57
timestamp 1698431365
transform 1 0 7728 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_65
timestamp 1698431365
transform 1 0 8624 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_76
timestamp 1698431365
transform 1 0 9856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_88
timestamp 1698431365
transform 1 0 11200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_92
timestamp 1698431365
transform 1 0 11648 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_108
timestamp 1698431365
transform 1 0 13440 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_112
timestamp 1698431365
transform 1 0 13888 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_121
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_220
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_240
timestamp 1698431365
transform 1 0 28224 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_256
timestamp 1698431365
transform 1 0 30016 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_264
timestamp 1698431365
transform 1 0 30912 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_268
timestamp 1698431365
transform 1 0 31360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_270
timestamp 1698431365
transform 1 0 31584 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_277
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_298
timestamp 1698431365
transform 1 0 34720 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_302
timestamp 1698431365
transform 1 0 35168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_333
timestamp 1698431365
transform 1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_337
timestamp 1698431365
transform 1 0 39088 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_345
timestamp 1698431365
transform 1 0 39984 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_369
timestamp 1698431365
transform 1 0 42672 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_377
timestamp 1698431365
transform 1 0 43568 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_381
timestamp 1698431365
transform 1 0 44016 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_383
timestamp 1698431365
transform 1 0 44240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_53
timestamp 1698431365
transform 1 0 7280 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_61
timestamp 1698431365
transform 1 0 8176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_95
timestamp 1698431365
transform 1 0 11984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_99
timestamp 1698431365
transform 1 0 12432 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_103
timestamp 1698431365
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_111
timestamp 1698431365
transform 1 0 13776 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_113
timestamp 1698431365
transform 1 0 14000 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_123
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_132
timestamp 1698431365
transform 1 0 16128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_136
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_151
timestamp 1698431365
transform 1 0 18256 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_167
timestamp 1698431365
transform 1 0 20048 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_209
timestamp 1698431365
transform 1 0 24752 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_213
timestamp 1698431365
transform 1 0 25200 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_223
timestamp 1698431365
transform 1 0 26320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_227
timestamp 1698431365
transform 1 0 26768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_231
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_239
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_285
timestamp 1698431365
transform 1 0 33264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_289
timestamp 1698431365
transform 1 0 33712 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_305
timestamp 1698431365
transform 1 0 35504 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_349
timestamp 1698431365
transform 1 0 40432 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_32
timestamp 1698431365
transform 1 0 4928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_36
timestamp 1698431365
transform 1 0 5376 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_52
timestamp 1698431365
transform 1 0 7168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_54
timestamp 1698431365
transform 1 0 7392 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_61
timestamp 1698431365
transform 1 0 8176 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_92
timestamp 1698431365
transform 1 0 11648 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_108
timestamp 1698431365
transform 1 0 13440 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_116
timestamp 1698431365
transform 1 0 14336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_125
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_137
timestamp 1698431365
transform 1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_161
timestamp 1698431365
transform 1 0 19376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_174
timestamp 1698431365
transform 1 0 20832 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_356
timestamp 1698431365
transform 1 0 41216 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_364
timestamp 1698431365
transform 1 0 42112 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_380
timestamp 1698431365
transform 1 0 43904 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_49
timestamp 1698431365
transform 1 0 6832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_54
timestamp 1698431365
transform 1 0 7392 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_70
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_78
timestamp 1698431365
transform 1 0 10080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_82
timestamp 1698431365
transform 1 0 10528 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_98
timestamp 1698431365
transform 1 0 12320 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_102
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_123
timestamp 1698431365
transform 1 0 15120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_129
timestamp 1698431365
transform 1 0 15792 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_137
timestamp 1698431365
transform 1 0 16688 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_151
timestamp 1698431365
transform 1 0 18256 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_167
timestamp 1698431365
transform 1 0 20048 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_201
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_207
timestamp 1698431365
transform 1 0 24528 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_223
timestamp 1698431365
transform 1 0 26320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_239
timestamp 1698431365
transform 1 0 28112 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_253
timestamp 1698431365
transform 1 0 29680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_257
timestamp 1698431365
transform 1 0 30128 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_270
timestamp 1698431365
transform 1 0 31584 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_302
timestamp 1698431365
transform 1 0 35168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_310
timestamp 1698431365
transform 1 0 36064 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_321
timestamp 1698431365
transform 1 0 37296 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_323
timestamp 1698431365
transform 1 0 37520 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_326
timestamp 1698431365
transform 1 0 37856 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_358
timestamp 1698431365
transform 1 0 41440 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_374
timestamp 1698431365
transform 1 0 43232 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_382
timestamp 1698431365
transform 1 0 44128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_34
timestamp 1698431365
transform 1 0 5152 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_42
timestamp 1698431365
transform 1 0 6048 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_46
timestamp 1698431365
transform 1 0 6496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_54
timestamp 1698431365
transform 1 0 7392 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698431365
transform 1 0 19040 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_162
timestamp 1698431365
transform 1 0 19488 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_195
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_197
timestamp 1698431365
transform 1 0 23408 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_218
timestamp 1698431365
transform 1 0 25760 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_226
timestamp 1698431365
transform 1 0 26656 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_230
timestamp 1698431365
transform 1 0 27104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_261
timestamp 1698431365
transform 1 0 30576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_265
timestamp 1698431365
transform 1 0 31024 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_273
timestamp 1698431365
transform 1 0 31920 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1698431365
transform 1 0 32368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_290
timestamp 1698431365
transform 1 0 33824 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_294
timestamp 1698431365
transform 1 0 34272 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_332
timestamp 1698431365
transform 1 0 38528 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_348
timestamp 1698431365
transform 1 0 40320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_69
timestamp 1698431365
transform 1 0 9072 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_73
timestamp 1698431365
transform 1 0 9520 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_93
timestamp 1698431365
transform 1 0 11760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_97
timestamp 1698431365
transform 1 0 12208 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_221
timestamp 1698431365
transform 1 0 26096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_225
timestamp 1698431365
transform 1 0 26544 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_321
timestamp 1698431365
transform 1 0 37296 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_336
timestamp 1698431365
transform 1 0 38976 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_340
timestamp 1698431365
transform 1 0 39424 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_344
timestamp 1698431365
transform 1 0 39872 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_371
timestamp 1698431365
transform 1 0 42896 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_375
timestamp 1698431365
transform 1 0 43344 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_383
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_32
timestamp 1698431365
transform 1 0 4928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_36
timestamp 1698431365
transform 1 0 5376 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_52
timestamp 1698431365
transform 1 0 7168 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_54
timestamp 1698431365
transform 1 0 7392 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_60
timestamp 1698431365
transform 1 0 8064 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_64
timestamp 1698431365
transform 1 0 8512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_86
timestamp 1698431365
transform 1 0 10976 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_98
timestamp 1698431365
transform 1 0 12320 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_130
timestamp 1698431365
transform 1 0 15904 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_138
timestamp 1698431365
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_314
timestamp 1698431365
transform 1 0 36512 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_330
timestamp 1698431365
transform 1 0 38304 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_340
timestamp 1698431365
transform 1 0 39424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_349
timestamp 1698431365
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_383
timestamp 1698431365
transform 1 0 44240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_41
timestamp 1698431365
transform 1 0 5936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_66
timestamp 1698431365
transform 1 0 8736 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_80
timestamp 1698431365
transform 1 0 10304 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_97
timestamp 1698431365
transform 1 0 12208 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_117
timestamp 1698431365
transform 1 0 14448 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_133
timestamp 1698431365
transform 1 0 16240 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_137
timestamp 1698431365
transform 1 0 16688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_139
timestamp 1698431365
transform 1 0 16912 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_209
timestamp 1698431365
transform 1 0 24752 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_225
timestamp 1698431365
transform 1 0 26544 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_233
timestamp 1698431365
transform 1 0 27440 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_237
timestamp 1698431365
transform 1 0 27888 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_263
timestamp 1698431365
transform 1 0 30800 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_298
timestamp 1698431365
transform 1 0 34720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_302
timestamp 1698431365
transform 1 0 35168 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_310
timestamp 1698431365
transform 1 0 36064 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_325
timestamp 1698431365
transform 1 0 37744 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_366
timestamp 1698431365
transform 1 0 42336 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_10
timestamp 1698431365
transform 1 0 2464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_12
timestamp 1698431365
transform 1 0 2688 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_42
timestamp 1698431365
transform 1 0 6048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_46
timestamp 1698431365
transform 1 0 6496 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_62
timestamp 1698431365
transform 1 0 8288 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_146
timestamp 1698431365
transform 1 0 17696 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_162
timestamp 1698431365
transform 1 0 19488 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_197
timestamp 1698431365
transform 1 0 23408 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_205
timestamp 1698431365
transform 1 0 24304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_270
timestamp 1698431365
transform 1 0 31584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_274
timestamp 1698431365
transform 1 0 32032 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_284
timestamp 1698431365
transform 1 0 33152 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_314
timestamp 1698431365
transform 1 0 36512 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_318
timestamp 1698431365
transform 1 0 36960 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_113
timestamp 1698431365
transform 1 0 14000 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_145
timestamp 1698431365
transform 1 0 17584 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_161
timestamp 1698431365
transform 1 0 19376 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_169
timestamp 1698431365
transform 1 0 20272 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_173
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_243
timestamp 1698431365
transform 1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_333
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_341
timestamp 1698431365
transform 1 0 39536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_345
timestamp 1698431365
transform 1 0 39984 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_353
timestamp 1698431365
transform 1 0 40880 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_357
timestamp 1698431365
transform 1 0 41328 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_26
timestamp 1698431365
transform 1 0 4256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_30
timestamp 1698431365
transform 1 0 4704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_36
timestamp 1698431365
transform 1 0 5376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_38
timestamp 1698431365
transform 1 0 5600 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_45
timestamp 1698431365
transform 1 0 6384 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_61
timestamp 1698431365
transform 1 0 8176 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_65
timestamp 1698431365
transform 1 0 8624 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_70
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_79
timestamp 1698431365
transform 1 0 10192 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_95
timestamp 1698431365
transform 1 0 11984 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_99
timestamp 1698431365
transform 1 0 12432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_101
timestamp 1698431365
transform 1 0 12656 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_106
timestamp 1698431365
transform 1 0 13216 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_133
timestamp 1698431365
transform 1 0 16240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_135
timestamp 1698431365
transform 1 0 16464 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_138
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_140
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_167
timestamp 1698431365
transform 1 0 20048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_169
timestamp 1698431365
transform 1 0 20272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_174
timestamp 1698431365
transform 1 0 20832 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_201
timestamp 1698431365
transform 1 0 23856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_203
timestamp 1698431365
transform 1 0 24080 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_208
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_235
timestamp 1698431365
transform 1 0 27664 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_237
timestamp 1698431365
transform 1 0 27888 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_240
timestamp 1698431365
transform 1 0 28224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_242
timestamp 1698431365
transform 1 0 28448 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_269
timestamp 1698431365
transform 1 0 31472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_271
timestamp 1698431365
transform 1 0 31696 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_274
timestamp 1698431365
transform 1 0 32032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_303
timestamp 1698431365
transform 1 0 35280 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_305
timestamp 1698431365
transform 1 0 35504 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_308
timestamp 1698431365
transform 1 0 35840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_310
timestamp 1698431365
transform 1 0 36064 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_337
timestamp 1698431365
transform 1 0 39088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_339
timestamp 1698431365
transform 1 0 39312 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_342
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_344
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_371
timestamp 1698431365
transform 1 0 42896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_373
timestamp 1698431365
transform 1 0 43120 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_376
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform 1 0 9520 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 5712 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698431365
transform 1 0 17136 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698431365
transform 1 0 20944 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698431365
transform 1 0 28560 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698431365
transform 1 0 36176 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698431365
transform 1 0 39984 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform 1 0 41440 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_50 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 44576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 44576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 44576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 44576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 44576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 44576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 44576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 44576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 44576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 44576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 44576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 44576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 44576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 44576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 44576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 44576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 44576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 44576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 44576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 44576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 44576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 44576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 44576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 44576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 44576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 44576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 44576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 44576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 44576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 44576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 44576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 44576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 44576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 44576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 44576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 44576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 44576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 44576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 44576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 44576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 44576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 44576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 44576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_112
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_113
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_114
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_115
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_118
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_119
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_120
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_121
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_122
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_123
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_124
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_125
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_126
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_127
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_128
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_129
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_130
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_131
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_132
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_133
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_134
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_135
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_136
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_137
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_138
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_139
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_140
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_141
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_142
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_143
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_144
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_145
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_146
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_147
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_148
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_149
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_150
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_151
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_152
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_153
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_154
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_155
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_156
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_157
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_158
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_159
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_160
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_161
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_162
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_163
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_164
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_165
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_166
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_167
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_168
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_169
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_170
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_171
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_172
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_173
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_174
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_175
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_176
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_177
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_178
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_179
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_180
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_181
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_182
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_183
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_184
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_185
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_186
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_187
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_188
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_189
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_190
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_191
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_192
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_193
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_194
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_195
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_196
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_197
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_198
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_199
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_200
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_201
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_202
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_209
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_210
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_212
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_213
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_214
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_215
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_216
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_217
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_218
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_219
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_220
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_221
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_222
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_223
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_224
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_225
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_226
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_227
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_228
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_229
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_230
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_231
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_232
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_233
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_234
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_235
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_236
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_237
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_238
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_239
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_240
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_241
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_242
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_243
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_244
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_245
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_246
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_247
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_248
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_249
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_250
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_251
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_252
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_253
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_254
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_255
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_256
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_257
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_258
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_259
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_260
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_261
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_262
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_263
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_264
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_265
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_266
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_267
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_268
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_269
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_270
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_271
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_272
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_273
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_274
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_275
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_276
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_277
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_278
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_279
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_280
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_281
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_282
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_283
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_284
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_285
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_286
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_287
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_288
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_289
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_290
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_291
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_292
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_293
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_294
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_295
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_296
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_297
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_298
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_299
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_300
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_301
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_302
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_303
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_304
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_305
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_306
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_307
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_308
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_309
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_310
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_311
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_312
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_313
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_314
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_315
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_316
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_317
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_318
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_319
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_320
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_321
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_322
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_323
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_324
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_325
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_326
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_327
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_328
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_329
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_330
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_331
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_332
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_333
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_334
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_335
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_336
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_337
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_338
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_339
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_340
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_341
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_342
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_343
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_344
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_345
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_346
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_347
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_348
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_349
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_350
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_351
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_352
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_353
timestamp 1698431365
transform 1 0 12768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_354
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_355
timestamp 1698431365
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_356
timestamp 1698431365
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_357
timestamp 1698431365
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_358
timestamp 1698431365
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_359
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_360
timestamp 1698431365
transform 1 0 39424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_361
timestamp 1698431365
transform 1 0 43232 0 -1 42336
box -86 -86 310 870
<< labels >>
flabel metal2 s 9408 45200 9520 46000 0 FreeSans 448 90 0 0 io_in
port 0 nsew signal input
flabel metal2 s 13216 45200 13328 46000 0 FreeSans 448 90 0 0 io_out[0]
port 1 nsew signal tristate
flabel metal2 s 17024 45200 17136 46000 0 FreeSans 448 90 0 0 io_out[1]
port 2 nsew signal tristate
flabel metal2 s 20832 45200 20944 46000 0 FreeSans 448 90 0 0 io_out[2]
port 3 nsew signal tristate
flabel metal2 s 24640 45200 24752 46000 0 FreeSans 448 90 0 0 io_out[3]
port 4 nsew signal tristate
flabel metal2 s 28448 45200 28560 46000 0 FreeSans 448 90 0 0 io_out[4]
port 5 nsew signal tristate
flabel metal2 s 32256 45200 32368 46000 0 FreeSans 448 90 0 0 io_out[5]
port 6 nsew signal tristate
flabel metal2 s 36064 45200 36176 46000 0 FreeSans 448 90 0 0 io_out[6]
port 7 nsew signal tristate
flabel metal2 s 39872 45200 39984 46000 0 FreeSans 448 90 0 0 io_out[7]
port 8 nsew signal tristate
flabel metal2 s 43680 45200 43792 46000 0 FreeSans 448 90 0 0 io_out[8]
port 9 nsew signal tristate
flabel metal2 s 5600 45200 5712 46000 0 FreeSans 448 90 0 0 rst_n
port 10 nsew signal input
flabel metal4 s 4448 3076 4768 42396 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 35168 3076 35488 42396 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 19808 3076 20128 42396 0 FreeSans 1280 90 0 0 vss
port 12 nsew ground bidirectional
flabel metal2 s 1792 45200 1904 46000 0 FreeSans 448 90 0 0 wb_clk_i
port 13 nsew signal input
rlabel metal1 22960 41552 22960 41552 0 vdd
rlabel metal1 22960 42336 22960 42336 0 vss
rlabel metal2 6440 39984 6440 39984 0 _000_
rlabel metal2 11368 39984 11368 39984 0 _001_
rlabel metal2 21112 39872 21112 39872 0 _002_
rlabel metal2 29288 39872 29288 39872 0 _003_
rlabel metal2 34216 40544 34216 40544 0 _004_
rlabel metal2 18200 39368 18200 39368 0 _005_
rlabel metal2 14280 39872 14280 39872 0 _006_
rlabel metal2 37352 21168 37352 21168 0 _007_
rlabel metal2 36568 18088 36568 18088 0 _008_
rlabel metal2 41720 18032 41720 18032 0 _009_
rlabel metal2 42000 12824 42000 12824 0 _010_
rlabel metal2 36064 13944 36064 13944 0 _011_
rlabel metal2 35840 9128 35840 9128 0 _012_
rlabel metal2 31528 14896 31528 14896 0 _013_
rlabel metal2 30408 10248 30408 10248 0 _014_
rlabel metal2 31640 18592 31640 18592 0 _015_
rlabel metal2 26600 19600 26600 19600 0 _016_
rlabel metal2 9688 39256 9688 39256 0 _017_
rlabel metal3 5152 35784 5152 35784 0 _018_
rlabel metal3 6104 36232 6104 36232 0 _019_
rlabel metal2 35896 35280 35896 35280 0 _020_
rlabel metal2 30856 34160 30856 34160 0 _021_
rlabel metal2 37128 33712 37128 33712 0 _022_
rlabel metal2 32032 39480 32032 39480 0 _023_
rlabel metal2 30408 29064 30408 29064 0 _024_
rlabel metal2 34552 24304 34552 24304 0 _025_
rlabel metal2 29960 24808 29960 24808 0 _026_
rlabel metal2 26040 28392 26040 28392 0 _027_
rlabel metal2 37072 29512 37072 29512 0 _028_
rlabel metal2 41496 30744 41496 30744 0 _029_
rlabel metal2 41832 27216 41832 27216 0 _030_
rlabel metal2 41832 34104 41832 34104 0 _031_
rlabel metal2 41608 22680 41608 22680 0 _032_
rlabel metal2 36232 25032 36232 25032 0 _033_
rlabel metal3 41104 39480 41104 39480 0 _034_
rlabel metal2 42056 38192 42056 38192 0 _035_
rlabel metal2 22120 21672 22120 21672 0 _036_
rlabel metal2 19544 18032 19544 18032 0 _037_
rlabel metal3 2996 16184 2996 16184 0 _038_
rlabel metal3 6776 16968 6776 16968 0 _039_
rlabel metal2 4200 12936 4200 12936 0 _040_
rlabel metal2 7784 8960 7784 8960 0 _041_
rlabel metal2 10248 12040 10248 12040 0 _042_
rlabel metal2 11816 7532 11816 7532 0 _043_
rlabel metal2 14280 6412 14280 6412 0 _044_
rlabel metal2 16520 6272 16520 6272 0 _045_
rlabel metal2 19880 4480 19880 4480 0 _046_
rlabel metal2 23464 5824 23464 5824 0 _047_
rlabel metal2 23688 19544 23688 19544 0 _048_
rlabel metal3 26712 15400 26712 15400 0 _049_
rlabel metal3 25704 9912 25704 9912 0 _050_
rlabel metal2 26040 7448 26040 7448 0 _051_
rlabel metal3 17024 30072 17024 30072 0 _052_
rlabel metal2 21840 27944 21840 27944 0 _053_
rlabel metal2 12656 28616 12656 28616 0 _054_
rlabel metal2 6888 30240 6888 30240 0 _055_
rlabel metal2 3192 21840 3192 21840 0 _056_
rlabel metal2 2632 23072 2632 23072 0 _057_
rlabel metal2 4200 31416 4200 31416 0 _058_
rlabel metal3 3584 28840 3584 28840 0 _059_
rlabel metal2 21560 36904 21560 36904 0 _060_
rlabel metal2 27944 36904 27944 36904 0 _061_
rlabel metal2 21560 32200 21560 32200 0 _062_
rlabel metal2 25816 34440 25816 34440 0 _063_
rlabel metal2 22680 26208 22680 26208 0 _064_
rlabel metal2 26824 36400 26824 36400 0 _065_
rlabel metal3 27776 34104 27776 34104 0 _066_
rlabel metal2 27384 34552 27384 34552 0 _067_
rlabel metal2 24248 36568 24248 36568 0 _068_
rlabel metal2 27720 34496 27720 34496 0 _069_
rlabel metal2 23800 33992 23800 33992 0 _070_
rlabel metal2 17864 34048 17864 34048 0 _071_
rlabel metal2 20104 35728 20104 35728 0 _072_
rlabel metal2 18088 36232 18088 36232 0 _073_
rlabel metal2 16016 34776 16016 34776 0 _074_
rlabel metal2 9576 24696 9576 24696 0 _075_
rlabel metal2 12488 27832 12488 27832 0 _076_
rlabel metal2 15176 24304 15176 24304 0 _077_
rlabel metal2 13944 28028 13944 28028 0 _078_
rlabel metal2 16296 22680 16296 22680 0 _079_
rlabel metal2 7616 21784 7616 21784 0 _080_
rlabel metal2 6552 23632 6552 23632 0 _081_
rlabel metal2 18536 22736 18536 22736 0 _082_
rlabel metal2 35504 19768 35504 19768 0 _083_
rlabel metal3 35448 20104 35448 20104 0 _084_
rlabel metal2 35056 20664 35056 20664 0 _085_
rlabel metal2 20216 23128 20216 23128 0 _086_
rlabel metal2 17976 24416 17976 24416 0 _087_
rlabel metal2 17808 22344 17808 22344 0 _088_
rlabel metal2 16464 19096 16464 19096 0 _089_
rlabel metal2 27272 16520 27272 16520 0 _090_
rlabel metal2 10808 25536 10808 25536 0 _091_
rlabel metal2 8904 17920 8904 17920 0 _092_
rlabel metal3 10528 19768 10528 19768 0 _093_
rlabel metal2 15176 28112 15176 28112 0 _094_
rlabel metal3 8624 20104 8624 20104 0 _095_
rlabel metal2 16296 19096 16296 19096 0 _096_
rlabel metal2 16632 21056 16632 21056 0 _097_
rlabel metal2 8120 12600 8120 12600 0 _098_
rlabel metal2 16184 19208 16184 19208 0 _099_
rlabel metal2 12376 18984 12376 18984 0 _100_
rlabel metal2 10360 17920 10360 17920 0 _101_
rlabel metal2 10584 20272 10584 20272 0 _102_
rlabel metal2 16856 20776 16856 20776 0 _103_
rlabel metal2 8344 21280 8344 21280 0 _104_
rlabel metal2 13160 17808 13160 17808 0 _105_
rlabel metal2 13832 21224 13832 21224 0 _106_
rlabel metal2 10248 24024 10248 24024 0 _107_
rlabel metal2 11480 21672 11480 21672 0 _108_
rlabel metal2 10304 12936 10304 12936 0 _109_
rlabel metal2 12376 21112 12376 21112 0 _110_
rlabel metal2 15400 21056 15400 21056 0 _111_
rlabel metal2 17024 22344 17024 22344 0 _112_
rlabel metal2 16296 31556 16296 31556 0 _113_
rlabel metal2 26600 35280 26600 35280 0 _114_
rlabel metal2 23688 36400 23688 36400 0 _115_
rlabel metal2 17192 35280 17192 35280 0 _116_
rlabel metal2 15400 34944 15400 34944 0 _117_
rlabel metal2 14728 34944 14728 34944 0 _118_
rlabel metal2 14784 34328 14784 34328 0 _119_
rlabel metal2 7112 35560 7112 35560 0 _120_
rlabel metal2 6888 38052 6888 38052 0 _121_
rlabel metal3 16912 35672 16912 35672 0 _122_
rlabel metal3 16856 35112 16856 35112 0 _123_
rlabel metal2 19096 36176 19096 36176 0 _124_
rlabel metal3 16296 36344 16296 36344 0 _125_
rlabel metal2 16296 35672 16296 35672 0 _126_
rlabel metal2 17136 22456 17136 22456 0 _127_
rlabel metal2 15960 24976 15960 24976 0 _128_
rlabel metal2 10808 35392 10808 35392 0 _129_
rlabel metal2 10584 36960 10584 36960 0 _130_
rlabel metal3 6944 39368 6944 39368 0 _131_
rlabel metal2 15288 35952 15288 35952 0 _132_
rlabel metal2 11592 35168 11592 35168 0 _133_
rlabel metal2 10024 35000 10024 35000 0 _134_
rlabel metal2 10584 34216 10584 34216 0 _135_
rlabel metal2 8008 35392 8008 35392 0 _136_
rlabel metal3 9240 39480 9240 39480 0 _137_
rlabel metal2 11200 14616 11200 14616 0 _138_
rlabel metal2 10248 37856 10248 37856 0 _139_
rlabel metal2 10136 38360 10136 38360 0 _140_
rlabel metal2 11760 38808 11760 38808 0 _141_
rlabel metal2 9128 39760 9128 39760 0 _142_
rlabel metal2 8064 39032 8064 39032 0 _143_
rlabel metal3 13048 39032 13048 39032 0 _144_
rlabel metal2 23464 30408 23464 30408 0 _145_
rlabel metal2 37352 20664 37352 20664 0 _146_
rlabel metal2 17976 16912 17976 16912 0 _147_
rlabel metal3 40712 16968 40712 16968 0 _148_
rlabel metal2 41608 16856 41608 16856 0 _149_
rlabel metal3 24920 24920 24920 24920 0 _150_
rlabel metal2 27552 24584 27552 24584 0 _151_
rlabel metal2 40488 12488 40488 12488 0 _152_
rlabel metal2 40712 17920 40712 17920 0 _153_
rlabel metal2 40264 13160 40264 13160 0 _154_
rlabel metal2 40824 12656 40824 12656 0 _155_
rlabel metal2 30968 9296 30968 9296 0 _156_
rlabel metal2 38472 12712 38472 12712 0 _157_
rlabel metal2 35896 12544 35896 12544 0 _158_
rlabel metal2 37688 12656 37688 12656 0 _159_
rlabel metal2 41552 12824 41552 12824 0 _160_
rlabel metal3 36904 11368 36904 11368 0 _161_
rlabel metal2 26712 24696 26712 24696 0 _162_
rlabel metal3 36960 13720 36960 13720 0 _163_
rlabel metal3 35784 11144 35784 11144 0 _164_
rlabel metal2 31304 11144 31304 11144 0 _165_
rlabel metal2 36008 10864 36008 10864 0 _166_
rlabel metal2 31752 14560 31752 14560 0 _167_
rlabel metal2 31976 14168 31976 14168 0 _168_
rlabel metal2 31640 10584 31640 10584 0 _169_
rlabel metal2 31696 18984 31696 18984 0 _170_
rlabel metal2 30072 19936 30072 19936 0 _171_
rlabel metal3 27832 23912 27832 23912 0 _172_
rlabel metal2 31136 19208 31136 19208 0 _173_
rlabel metal2 21336 28672 21336 28672 0 _174_
rlabel metal2 26712 19600 26712 19600 0 _175_
rlabel metal2 26600 28672 26600 28672 0 _176_
rlabel metal2 26264 28728 26264 28728 0 _177_
rlabel metal2 33096 26684 33096 26684 0 _178_
rlabel metal3 34552 33320 34552 33320 0 _179_
rlabel metal2 39032 28616 39032 28616 0 _180_
rlabel metal2 24696 24528 24696 24528 0 _181_
rlabel metal2 40040 31192 40040 31192 0 _182_
rlabel metal2 37240 32984 37240 32984 0 _183_
rlabel metal2 25648 25256 25648 25256 0 _184_
rlabel metal2 25368 31752 25368 31752 0 _185_
rlabel metal2 30632 30576 30632 30576 0 _186_
rlabel metal2 31192 33320 31192 33320 0 _187_
rlabel metal3 36008 28392 36008 28392 0 _188_
rlabel metal2 30800 32760 30800 32760 0 _189_
rlabel metal2 39480 30016 39480 30016 0 _190_
rlabel metal2 37352 33376 37352 33376 0 _191_
rlabel metal2 37072 32760 37072 32760 0 _192_
rlabel metal2 31752 31864 31752 31864 0 _193_
rlabel metal2 32088 32424 32088 32424 0 _194_
rlabel metal2 4648 28000 4648 28000 0 _195_
rlabel metal2 31640 27720 31640 27720 0 _196_
rlabel metal2 30968 29792 30968 29792 0 _197_
rlabel metal2 31640 24472 31640 24472 0 _198_
rlabel metal2 40936 25704 40936 25704 0 _199_
rlabel metal2 31304 24976 31304 24976 0 _200_
rlabel metal2 31976 25480 31976 25480 0 _201_
rlabel metal2 30856 25760 30856 25760 0 _202_
rlabel metal2 29960 28560 29960 28560 0 _203_
rlabel metal2 29456 28840 29456 28840 0 _204_
rlabel metal3 38248 30072 38248 30072 0 _205_
rlabel metal3 36008 30072 36008 30072 0 _206_
rlabel metal2 41552 29624 41552 29624 0 _207_
rlabel metal3 40768 30968 40768 30968 0 _208_
rlabel metal2 41608 37856 41608 37856 0 _209_
rlabel metal2 41608 28616 41608 28616 0 _210_
rlabel metal2 41832 26656 41832 26656 0 _211_
rlabel metal2 42280 26936 42280 26936 0 _212_
rlabel metal2 42168 32984 42168 32984 0 _213_
rlabel metal2 25816 37912 25816 37912 0 _214_
rlabel metal2 41720 33824 41720 33824 0 _215_
rlabel metal2 40936 24920 40936 24920 0 _216_
rlabel metal2 41608 24248 41608 24248 0 _217_
rlabel metal2 41832 23296 41832 23296 0 _218_
rlabel metal2 37912 32648 37912 32648 0 _219_
rlabel metal3 37128 26936 37128 26936 0 _220_
rlabel metal2 6440 28672 6440 28672 0 _221_
rlabel metal2 36456 25872 36456 25872 0 _222_
rlabel metal2 39816 35392 39816 35392 0 _223_
rlabel metal2 40824 38136 40824 38136 0 _224_
rlabel metal2 40376 39312 40376 39312 0 _225_
rlabel metal2 41832 38080 41832 38080 0 _226_
rlabel metal2 42280 37912 42280 37912 0 _227_
rlabel metal3 22288 23800 22288 23800 0 _228_
rlabel metal2 21672 25984 21672 25984 0 _229_
rlabel metal2 21224 24696 21224 24696 0 _230_
rlabel metal2 23912 25816 23912 25816 0 _231_
rlabel metal2 22456 24248 22456 24248 0 _232_
rlabel metal3 17024 24696 17024 24696 0 _233_
rlabel metal2 16856 24248 16856 24248 0 _234_
rlabel metal2 16072 25872 16072 25872 0 _235_
rlabel metal2 16632 26320 16632 26320 0 _236_
rlabel metal2 20888 24472 20888 24472 0 _237_
rlabel metal3 22064 23912 22064 23912 0 _238_
rlabel metal3 17024 16856 17024 16856 0 _239_
rlabel metal2 21112 15344 21112 15344 0 _240_
rlabel metal2 18088 15232 18088 15232 0 _241_
rlabel metal3 17304 14616 17304 14616 0 _242_
rlabel metal3 15736 14504 15736 14504 0 _243_
rlabel metal3 16464 15176 16464 15176 0 _244_
rlabel metal3 17024 15400 17024 15400 0 _245_
rlabel metal2 17752 16520 17752 16520 0 _246_
rlabel metal3 12880 16968 12880 16968 0 _247_
rlabel metal2 20888 15736 20888 15736 0 _248_
rlabel metal3 10192 12824 10192 12824 0 _249_
rlabel metal2 12152 16128 12152 16128 0 _250_
rlabel metal2 12376 16408 12376 16408 0 _251_
rlabel metal3 10304 12936 10304 12936 0 _252_
rlabel metal2 9240 12656 9240 12656 0 _253_
rlabel metal2 8680 13496 8680 13496 0 _254_
rlabel metal2 8792 13272 8792 13272 0 _255_
rlabel metal2 9912 15904 9912 15904 0 _256_
rlabel metal2 8568 13216 8568 13216 0 _257_
rlabel metal2 9240 13272 9240 13272 0 _258_
rlabel metal2 8176 9912 8176 9912 0 _259_
rlabel metal2 8792 11704 8792 11704 0 _260_
rlabel metal2 9240 11368 9240 11368 0 _261_
rlabel metal2 8680 10024 8680 10024 0 _262_
rlabel metal2 8344 10248 8344 10248 0 _263_
rlabel metal2 12936 11312 12936 11312 0 _264_
rlabel metal2 12152 11312 12152 11312 0 _265_
rlabel metal2 11144 13104 11144 13104 0 _266_
rlabel metal2 13944 10640 13944 10640 0 _267_
rlabel metal2 12264 10192 12264 10192 0 _268_
rlabel metal2 12208 9240 12208 9240 0 _269_
rlabel metal2 16520 9380 16520 9380 0 _270_
rlabel metal3 14504 9800 14504 9800 0 _271_
rlabel metal2 16184 9688 16184 9688 0 _272_
rlabel metal2 15176 9184 15176 9184 0 _273_
rlabel metal2 14896 9128 14896 9128 0 _274_
rlabel metal2 18032 9128 18032 9128 0 _275_
rlabel metal2 17416 9296 17416 9296 0 _276_
rlabel metal2 17864 10136 17864 10136 0 _277_
rlabel metal2 17304 10024 17304 10024 0 _278_
rlabel metal3 20664 10024 20664 10024 0 _279_
rlabel metal3 22792 15400 22792 15400 0 _280_
rlabel metal2 18312 9240 18312 9240 0 _281_
rlabel metal2 21672 10864 21672 10864 0 _282_
rlabel metal2 20944 9016 20944 9016 0 _283_
rlabel metal2 20216 9632 20216 9632 0 _284_
rlabel metal2 22904 12656 22904 12656 0 _285_
rlabel metal2 23296 15288 23296 15288 0 _286_
rlabel metal2 21672 13160 21672 13160 0 _287_
rlabel metal2 21560 12376 21560 12376 0 _288_
rlabel metal2 21728 6664 21728 6664 0 _289_
rlabel metal3 22120 30296 22120 30296 0 _290_
rlabel metal3 25256 15512 25256 15512 0 _291_
rlabel metal2 22904 15512 22904 15512 0 _292_
rlabel metal3 23968 15960 23968 15960 0 _293_
rlabel metal2 23240 17976 23240 17976 0 _294_
rlabel metal3 25200 15960 25200 15960 0 _295_
rlabel metal2 23912 15008 23912 15008 0 _296_
rlabel metal2 24584 15568 24584 15568 0 _297_
rlabel metal3 25144 10808 25144 10808 0 _298_
rlabel metal2 25144 10080 25144 10080 0 _299_
rlabel metal2 24248 12096 24248 12096 0 _300_
rlabel metal3 25760 11256 25760 11256 0 _301_
rlabel metal2 24808 10472 24808 10472 0 _302_
rlabel metal2 25424 9800 25424 9800 0 _303_
rlabel metal3 25368 9128 25368 9128 0 _304_
rlabel metal2 25928 9296 25928 9296 0 _305_
rlabel metal2 25480 8960 25480 8960 0 _306_
rlabel metal2 15400 28168 15400 28168 0 _307_
rlabel metal2 15960 28896 15960 28896 0 _308_
rlabel metal2 15960 30408 15960 30408 0 _309_
rlabel metal2 15176 28672 15176 28672 0 _310_
rlabel metal3 19432 28616 19432 28616 0 _311_
rlabel metal2 22904 28392 22904 28392 0 _312_
rlabel metal2 12936 25984 12936 25984 0 _313_
rlabel metal2 11592 26992 11592 26992 0 _314_
rlabel metal2 12376 28336 12376 28336 0 _315_
rlabel metal2 10808 26320 10808 26320 0 _316_
rlabel metal2 10584 25928 10584 25928 0 _317_
rlabel metal2 11144 26600 11144 26600 0 _318_
rlabel metal2 11368 28168 11368 28168 0 _319_
rlabel metal3 8400 25368 8400 25368 0 _320_
rlabel metal2 6216 24584 6216 24584 0 _321_
rlabel metal3 6720 25480 6720 25480 0 _322_
rlabel metal2 6104 24528 6104 24528 0 _323_
rlabel metal2 7224 24080 7224 24080 0 _324_
rlabel metal2 4648 24752 4648 24752 0 _325_
rlabel metal3 4592 24920 4592 24920 0 _326_
rlabel metal2 4760 25144 4760 25144 0 _327_
rlabel metal2 4424 25536 4424 25536 0 _328_
rlabel metal3 4872 28392 4872 28392 0 _329_
rlabel metal2 5992 25928 5992 25928 0 _330_
rlabel metal2 5768 28000 5768 28000 0 _331_
rlabel metal2 4312 29792 4312 29792 0 _332_
rlabel metal2 5432 28112 5432 28112 0 _333_
rlabel metal3 6440 28504 6440 28504 0 _334_
rlabel metal2 21896 37296 21896 37296 0 _335_
rlabel metal2 27496 36568 27496 36568 0 _336_
rlabel metal2 26712 32872 26712 32872 0 _337_
rlabel metal2 27048 33488 27048 33488 0 _338_
rlabel metal2 21896 32088 21896 32088 0 _339_
rlabel metal2 24136 30576 24136 30576 0 _340_
rlabel metal2 25816 31808 25816 31808 0 _341_
rlabel metal2 10248 34944 10248 34944 0 bcd\[0\]
rlabel metal2 4760 35504 4760 35504 0 bcd\[1\]
rlabel metal2 7112 34048 7112 34048 0 bcd\[2\]
rlabel metal2 14952 30240 14952 30240 0 clkdiv\[0\]
rlabel metal2 17192 27384 17192 27384 0 clkdiv\[1\]
rlabel metal2 11480 28336 11480 28336 0 clkdiv\[2\]
rlabel metal3 9464 27048 9464 27048 0 clkdiv\[3\]
rlabel metal2 11816 20720 11816 20720 0 clkdiv\[4\]
rlabel metal2 7112 21168 7112 21168 0 clkdiv\[5\]
rlabel metal2 5880 28616 5880 28616 0 clkdiv\[6\]
rlabel metal2 4872 28952 4872 28952 0 clkdiv\[7\]
rlabel metal3 27720 22232 27720 22232 0 clknet_0_wb_clk_i
rlabel metal2 7000 11200 7000 11200 0 clknet_3_0__leaf_wb_clk_i
rlabel metal2 13608 4704 13608 4704 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 2184 30576 2184 30576 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 20328 40432 20328 40432 0 clknet_3_3__leaf_wb_clk_i
rlabel metal2 28672 6104 28672 6104 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 39032 20328 39032 20328 0 clknet_3_5__leaf_wb_clk_i
rlabel metal2 25368 27944 25368 27944 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 31528 39928 31528 39928 0 clknet_3_7__leaf_wb_clk_i
rlabel metal3 16744 20496 16744 20496 0 counter\[0\]
rlabel metal2 22232 5040 22232 5040 0 counter\[10\]
rlabel metal2 21112 5600 21112 5600 0 counter\[11\]
rlabel metal2 25816 17864 25816 17864 0 counter\[12\]
rlabel metal2 26096 15176 26096 15176 0 counter\[13\]
rlabel metal2 28616 11648 28616 11648 0 counter\[14\]
rlabel metal2 28448 9688 28448 9688 0 counter\[15\]
rlabel metal2 16184 17976 16184 17976 0 counter\[1\]
rlabel metal3 7224 16856 7224 16856 0 counter\[2\]
rlabel metal2 10136 17472 10136 17472 0 counter\[3\]
rlabel metal2 8008 12656 8008 12656 0 counter\[4\]
rlabel metal3 6608 8344 6608 8344 0 counter\[5\]
rlabel metal2 4872 11872 4872 11872 0 counter\[6\]
rlabel metal2 9688 7168 9688 7168 0 counter\[7\]
rlabel metal2 19096 5768 19096 5768 0 counter\[8\]
rlabel metal2 18648 5544 18648 5544 0 counter\[9\]
rlabel metal2 9576 41944 9576 41944 0 io_in
rlabel metal2 14504 41888 14504 41888 0 io_out[0]
rlabel metal2 17640 45304 17640 45304 0 io_out[1]
rlabel metal3 21504 41832 21504 41832 0 io_out[2]
rlabel metal3 25312 41832 25312 41832 0 io_out[3]
rlabel metal3 29120 41832 29120 41832 0 io_out[4]
rlabel metal2 32872 45304 32872 45304 0 io_out[5]
rlabel metal3 36736 41832 36736 41832 0 io_out[6]
rlabel metal3 40544 41832 40544 41832 0 io_out[7]
rlabel metal2 43736 43274 43736 43274 0 io_out[8]
rlabel metal2 24584 37072 24584 37072 0 lfsr\[0\]
rlabel metal2 41664 26488 41664 26488 0 lfsr\[10\]
rlabel metal2 41832 35336 41832 35336 0 lfsr\[11\]
rlabel metal2 43736 23464 43736 23464 0 lfsr\[12\]
rlabel metal2 39256 25984 39256 25984 0 lfsr\[13\]
rlabel metal3 39256 38920 39256 38920 0 lfsr\[14\]
rlabel metal2 44072 38304 44072 38304 0 lfsr\[15\]
rlabel metal2 32088 34216 32088 34216 0 lfsr\[1\]
rlabel metal2 25144 33096 25144 33096 0 lfsr\[2\]
rlabel metal2 31584 31080 31584 31080 0 lfsr\[4\]
rlabel metal2 33320 26656 33320 26656 0 lfsr\[5\]
rlabel metal2 31304 23632 31304 23632 0 lfsr\[6\]
rlabel metal2 29288 28280 29288 28280 0 lfsr\[7\]
rlabel metal2 34888 29232 34888 29232 0 lfsr\[8\]
rlabel metal2 40152 30688 40152 30688 0 lfsr\[9\]
rlabel metal2 38920 21448 38920 21448 0 m_clkdiv\[0\]
rlabel metal2 38696 18760 38696 18760 0 m_clkdiv\[1\]
rlabel metal2 41496 17416 41496 17416 0 m_clkdiv\[2\]
rlabel metal2 41384 14000 41384 14000 0 m_clkdiv\[3\]
rlabel metal2 37688 14784 37688 14784 0 m_clkdiv\[4\]
rlabel metal2 37688 11760 37688 11760 0 m_clkdiv\[5\]
rlabel metal2 33432 16072 33432 16072 0 m_clkdiv\[6\]
rlabel metal2 31864 11424 31864 11424 0 m_clkdiv\[7\]
rlabel metal2 31416 18928 31416 18928 0 m_clkdiv\[8\]
rlabel metal2 29960 19600 29960 19600 0 m_clkdiv\[9\]
rlabel metal2 9744 28056 9744 28056 0 net1
rlabel metal2 28280 40264 28280 40264 0 net10
rlabel metal3 38024 39704 38024 39704 0 net11
rlabel metal2 9520 34104 9520 34104 0 net2
rlabel metal2 5880 40208 5880 40208 0 net3
rlabel metal2 16856 41104 16856 41104 0 net4
rlabel metal2 20328 39816 20328 39816 0 net5
rlabel metal2 24920 41104 24920 41104 0 net6
rlabel metal2 23240 41104 23240 41104 0 net7
rlabel metal2 31416 41104 31416 41104 0 net8
rlabel metal2 36344 41104 36344 41104 0 net9
rlabel metal2 24192 36232 24192 36232 0 r_counter\[0\]
rlabel metal3 30184 36456 30184 36456 0 r_counter\[1\]
rlabel metal2 23912 32872 23912 32872 0 r_counter\[2\]
rlabel metal2 5880 42504 5880 42504 0 rst_n
rlabel metal2 21672 22344 21672 22344 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 46000 46000
<< end >>
