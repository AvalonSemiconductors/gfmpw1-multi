* NGSPICE file created from diceroll.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

.subckt diceroll io_in io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] rst_n vdd vss wb_clk_i
XFILLER_0_49_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_3__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_501_ lfsr\[7\] _182_ _202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_432_ m_clkdiv\[1\] m_clkdiv\[0\] _148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_363_ _080_ _084_ _088_ _089_ _090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_415_ _122_ _018_ _138_ _139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_346_ _064_ _070_ _072_ _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__679__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_680_ _006_ clknet_3_2__leaf_wb_clk_i net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__717__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_732_ _058_ clknet_3_3__leaf_wb_clk_i clkdiv\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_3_7__f_wb_clk_i clknet_0_wb_clk_i clknet_3_7__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_594_ counter\[10\] _275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_663_ _189_ _330_ _059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput7 net7 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_715_ _041_ clknet_3_0__leaf_wb_clk_i counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_577_ counter\[6\] _257_ _248_ _261_ _262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_646_ _316_ _314_ _312_ _309_ _318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_49_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_500_ _200_ _179_ _201_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_37_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_431_ _145_ _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_362_ net1 _089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_23_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_629_ _304_ _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_414_ _134_ _138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_345_ _071_ lfsr\[0\] _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__477__A1 _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__468__A1 _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_24_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_6__f_wb_clk_i clknet_0_wb_clk_i clknet_3_6__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__622__A1 _273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__613__A1 _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_731_ _057_ clknet_3_3__leaf_wb_clk_i clkdiv\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_662_ clkdiv\[7\] _327_ _329_ _233_ _330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_41_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_593_ _271_ _267_ _274_ _260_ _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_29_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput10 net10 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput8 net8 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_43_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_714_ _040_ clknet_3_0__leaf_wb_clk_i counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_645_ _314_ _310_ _313_ _316_ _317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_576_ counter\[6\] _255_ counter\[4\] _251_ _261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_1_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__707__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_430_ m_clkdiv\[0\] _146_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_361_ _085_ _086_ _087_ _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_23_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_628_ _152_ _302_ _303_ _304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_13_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_559_ counter\[3\] _246_ _247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__495__A2 _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_413_ _137_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_344_ r_counter\[0\] _071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5__f_wb_clk_i clknet_0_wb_clk_i clknet_3_5__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__395__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_592_ _270_ _257_ _272_ _273_ _274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_730_ _056_ clknet_3_0__leaf_wb_clk_i clkdiv\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_661_ _081_ _089_ _326_ _329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_41_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__522__A1 _196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput9 net9 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput11 net11 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_644_ _109_ _316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_575_ _256_ _252_ _259_ _260_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_713_ _039_ clknet_3_1__leaf_wb_clk_i counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_360_ m_clkdiv\[3\] m_clkdiv\[2\] m_clkdiv\[5\] m_clkdiv\[4\] _087_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_23_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_558_ _236_ _246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_627_ counter\[15\] _229_ _299_ _303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_489_ lfsr\[4\] _186_ _193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__601__B _281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_4__f_wb_clk_i clknet_0_wb_clk_i clknet_3_4__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_412_ _125_ _129_ _136_ _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_343_ r_counter\[2\] lfsr\[2\] _069_ _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_36_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__692__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_660_ _328_ _058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_591_ _230_ _177_ _273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__480__I _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_712_ _038_ clknet_3_0__leaf_wb_clk_i counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__730__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__475__I _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_0__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_574_ _145_ _260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_643_ _314_ _310_ _315_ _260_ _054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_26_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_3__f_wb_clk_i clknet_0_wb_clk_i clknet_3_3__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__509__B _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_488_ _178_ _192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_557_ _242_ _245_ _146_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_626_ _277_ _298_ _301_ _302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_411_ net2 _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_342_ _065_ _067_ _068_ _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_609_ counter\[12\] _288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_590_ _270_ _265_ _266_ _272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_output10_I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_2__f_wb_clk_i clknet_0_wb_clk_i clknet_3_2__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__682__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__530__B _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_642_ _314_ _310_ _313_ _315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_711_ _037_ clknet_3_0__leaf_wb_clk_i counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_573_ _255_ _257_ _248_ _258_ _259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_625_ counter\[15\] _301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_487_ _190_ _179_ _191_ _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_556_ _239_ _243_ _244_ _245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_14_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input1_I io_in vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__720__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_410_ _017_ _130_ _019_ _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_341_ _066_ lfsr\[1\] _068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_608_ _286_ _287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_19_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_539_ _225_ _226_ net1 _230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_49_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__552__A1 _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__517__C _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_3_1__f_wb_clk_i clknet_0_wb_clk_i clknet_3_1__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__494__I _196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__618__B _281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_45_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_572_ _255_ _250_ _251_ _258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_710_ _036_ clknet_3_1__leaf_wb_clk_i counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_641_ _112_ _314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_624_ _296_ _297_ _299_ _300_ _157_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_555_ _111_ _235_ _224_ _244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_486_ lfsr\[2\] _182_ _183_ _191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_340_ _066_ lfsr\[1\] _067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__695__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_607_ counter\[11\] _275_ _266_ _285_ _286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_538_ _228_ _229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_469_ lfsr\[1\] _176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_0__f_wb_clk_i clknet_0_wb_clk_i clknet_3_0__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__710__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__733__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__454__B _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_571_ _236_ _257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_640_ _311_ _313_ _281_ _053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__539__B net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__673__A1 _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__655__A1 _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_485_ net11 _190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_623_ counter\[14\] _246_ _300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_554_ _094_ _100_ _104_ _243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__628__A1 _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_606_ _270_ counter\[8\] _285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_468_ _173_ _175_ _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_537_ _088_ _227_ _228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_399_ _123_ _124_ _125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__685__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__700__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__723__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_570_ _255_ _256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_699_ _025_ clknet_3_7__leaf_wb_clk_i lfsr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__664__A2 _196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_622_ _273_ _298_ _299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_484_ _176_ _185_ _187_ _189_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_553_ _111_ _237_ _242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__591__A1 _230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_605_ _282_ _284_ _281_ _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_398_ _118_ _124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_467_ m_clkdiv\[9\] _174_ _175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_536_ _089_ _225_ _226_ _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_42_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_33_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__537__A1 _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_519_ lfsr\[11\] _209_ _188_ _215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__675__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__698__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_698_ _024_ clknet_3_7__leaf_wb_clk_i lfsr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_621_ counter\[14\] _292_ counter\[12\] _286_ _298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_552_ _173_ _241_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_483_ _188_ _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__713__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__736__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_36_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_604_ _275_ _276_ _283_ _284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_535_ _081_ _098_ _099_ _079_ _226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_397_ bcd\[1\] _123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_466_ m_clkdiv\[8\] _171_ _174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_5__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_518_ lfsr\[12\] _214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_449_ _151_ _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_697_ _023_ clknet_3_7__leaf_wb_clk_i net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__672__B net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_620_ _292_ _288_ _287_ _297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_551_ _235_ _237_ _239_ _240_ _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_482_ _150_ _188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__511__I _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__688__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_603_ counter\[11\] _277_ _283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_465_ _157_ _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_27_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_534_ _109_ _103_ _082_ _083_ _225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_396_ _122_ _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__703__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_517_ _208_ _197_ _212_ _213_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_448_ m_clkdiv\[4\] _158_ _161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_379_ _103_ _104_ counter\[0\] _105_ _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__726__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__484__C _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__659__C _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_696_ _022_ clknet_3_7__leaf_wb_clk_i lfsr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_481_ lfsr\[2\] _186_ _187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_550_ _235_ _224_ _240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_679_ _004_ clknet_3_6__leaf_wb_clk_i net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_602_ _246_ _278_ counter\[11\] _282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_464_ m_clkdiv\[8\] _171_ _172_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_533_ counter\[0\] _224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_27_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_395_ net2 _119_ _121_ _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_49_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_378_ clkdiv\[0\] _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_447_ _160_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_516_ _145_ _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__678__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__716__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_695_ _021_ clknet_3_7__leaf_wb_clk_i lfsr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_480_ _181_ _186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__435__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_678_ _003_ clknet_3_6__leaf_wb_clk_i net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_601_ _279_ _280_ _281_ _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_4_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_394_ _120_ _118_ _121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_39_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__593__C _260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_463_ m_clkdiv\[8\] _171_ _168_ _172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_27_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_532_ _218_ _185_ _223_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_515_ _196_ _211_ _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_446_ _156_ _159_ _160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_377_ counter\[2\] _104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__443__I _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_429_ _145_ _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput1 io_in net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_694_ _020_ clknet_3_7__leaf_wb_clk_i lfsr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__706__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_677_ _002_ clknet_3_6__leaf_wb_clk_i net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__729__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_600_ _157_ _281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_531_ lfsr\[15\] _209_ _188_ _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_393_ bcd\[0\] _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_462_ _147_ _170_ _171_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_27_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_3_2__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_729_ _055_ clknet_3_2__leaf_wb_clk_i clkdiv\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_514_ _180_ lfsr\[11\] _211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_376_ clkdiv\[2\] _103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_445_ _157_ _158_ _159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_428_ _136_ _145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_359_ m_clkdiv\[1\] m_clkdiv\[0\] _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput2 rst_n net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__603__A2 _277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__521__A1 _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_693_ _019_ clknet_3_2__leaf_wb_clk_i bcd\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_676_ _001_ clknet_3_3__leaf_wb_clk_i net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_461_ m_clkdiv\[7\] _167_ _164_ _171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_530_ _221_ _222_ _146_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_27_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_392_ _073_ _074_ _077_ _118_ _119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_10_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_31_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_728_ _054_ clknet_3_2__leaf_wb_clk_i clkdiv\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_659_ _098_ _325_ _327_ _152_ _328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_45_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__547__I _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_513_ _208_ _179_ _210_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_444_ _155_ _153_ _158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__457__I _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__719__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_375_ _098_ _093_ counter\[5\] _099_ _101_ _102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_46_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_427_ _144_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_43_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_358_ m_clkdiv\[7\] m_clkdiv\[6\] m_clkdiv\[9\] m_clkdiv\[8\] _085_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__691__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__470__I _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_692_ _018_ clknet_3_2__leaf_wb_clk_i bcd\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__465__I _157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__497__A1 _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_675_ _000_ clknet_3_2__leaf_wb_clk_i net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_460_ _167_ _165_ m_clkdiv\[7\] _170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_391_ _090_ _097_ _102_ _117_ _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_10_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_727_ _053_ clknet_3_2__leaf_wb_clk_i clkdiv\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_589_ _270_ _271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_658_ _312_ _326_ _233_ _327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_512_ lfsr\[9\] _209_ _183_ _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_374_ _099_ counter\[5\] _100_ _083_ _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_443_ _136_ _157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__558__I _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_426_ _135_ _140_ _144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_43_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_357_ _081_ clkdiv\[6\] _082_ _083_ _084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_11_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__709__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_409_ _134_ _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__610__B _277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__571__I _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_691_ _017_ clknet_3_2__leaf_wb_clk_i bcd\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__681__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__605__B _281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__430__A2 _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_674_ _005_ clknet_3_3__leaf_wb_clk_i net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__476__I _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_390_ _106_ _110_ _113_ _116_ _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_35_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_726_ _052_ clknet_3_3__leaf_wb_clk_i clkdiv\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_657_ _098_ clkdiv\[5\] _320_ _326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_588_ counter\[9\] _270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_18_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_511_ _181_ _209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_442_ _155_ _153_ _156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_373_ counter\[0\] _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_709_ _035_ clknet_3_7__leaf_wb_clk_i lfsr\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_425_ _122_ _138_ _018_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__417__C _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_356_ clkdiv\[0\] _083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__515__A1 _196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_408_ net2 _132_ _133_ _134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_339_ r_counter\[1\] _066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__506__A1 _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_690_ _016_ clknet_3_4__leaf_wb_clk_i m_clkdiv\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_48_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_673_ _197_ _227_ _336_ _194_ _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_21_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_656_ clkdiv\[5\] _232_ _320_ _325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_587_ _268_ _269_ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_725_ _051_ clknet_3_4__leaf_wb_clk_i counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__694__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_510_ lfsr\[10\] _208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_441_ m_clkdiv\[3\] _155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_35_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_372_ _078_ _099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_708_ _034_ clknet_3_6__leaf_wb_clk_i lfsr\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_639_ _312_ _181_ _313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__523__C _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_424_ _143_ _142_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_43_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_355_ clkdiv\[1\] _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__732__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_407_ bcd\[2\] _118_ _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_338_ r_counter\[0\] lfsr\[0\] _065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_22_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__433__A1 _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__672__A1 _230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__663__A1 _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_672_ _230_ _203_ net10 _336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__632__B _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_35_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_724_ _050_ clknet_3_4__leaf_wb_clk_i counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_655_ _194_ _323_ _324_ _057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_586_ _265_ _266_ _162_ _269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_371_ clkdiv\[6\] _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_440_ _149_ _154_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_707_ _033_ clknet_3_5__leaf_wb_clk_i lfsr\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_638_ net1 _312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_569_ counter\[5\] _255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__684__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_423_ _138_ _018_ _143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_43_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_354_ clkdiv\[7\] _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_23_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__624__C _157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__640__B _281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_3_7__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_337_ r_counter\[1\] lfsr\[1\] _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_406_ _124_ _128_ _131_ _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_22_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__722__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_16_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_671_ _213_ _335_ _062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_723_ _049_ clknet_3_4__leaf_wb_clk_i counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_654_ _099_ _089_ _233_ _320_ _324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_585_ _265_ _237_ _239_ _267_ _268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_370_ _091_ _092_ _096_ _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_23_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_706_ _032_ clknet_3_5__leaf_wb_clk_i lfsr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_637_ _082_ _306_ _310_ _311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_499_ lfsr\[5\] _182_ _183_ _201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_568_ _253_ _254_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__463__B _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__527__A1 _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_422_ _017_ _130_ _142_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_353_ _078_ _079_ clkdiv\[3\] clkdiv\[2\] _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__458__B _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_405_ _070_ _076_ _131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__674__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__697__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_670_ r_counter\[2\] _333_ _335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__712__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_653_ _305_ _321_ clkdiv\[5\] _323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_722_ _048_ clknet_3_4__leaf_wb_clk_i counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_584_ _265_ _266_ _267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__735__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__643__C _260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_567_ _250_ _251_ _162_ _254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_705_ _031_ clknet_3_7__leaf_wb_clk_i lfsr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_636_ _309_ _310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_498_ lfsr\[6\] _200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_39_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_421_ _134_ _140_ _142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_352_ clkdiv\[4\] _079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_619_ counter\[14\] _296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__445__A1 _157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_404_ _125_ _129_ _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__651__C _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_26_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__411__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__687__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_721_ _047_ clknet_3_4__leaf_wb_clk_i counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__567__B _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_583_ _107_ _261_ _266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_652_ _322_ _056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_32_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_13_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_704_ _030_ clknet_3_7__leaf_wb_clk_i lfsr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_566_ _250_ _237_ _239_ _252_ _253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_635_ _232_ _308_ _309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_497_ _194_ _198_ _199_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_26_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__702__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_420_ _017_ _141_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_351_ clkdiv\[5\] _078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__725__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_618_ _293_ _295_ _281_ _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_549_ _238_ _239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_40_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_403_ _124_ _126_ _128_ _129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_28_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_1_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__639__A2 _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_720_ _046_ clknet_3_1__leaf_wb_clk_i counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_582_ counter\[8\] _265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_651_ _079_ _319_ _321_ _305_ _168_ _322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_703_ _029_ clknet_3_7__leaf_wb_clk_i lfsr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_634_ _115_ _105_ _308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_46_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_496_ lfsr\[5\] _192_ _199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_565_ _250_ _251_ _252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__677__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_350_ _075_ _076_ _077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_617_ _294_ _288_ _273_ _287_ _295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_clkbuf_3_4__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_479_ _178_ _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_548_ _195_ _231_ _238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__490__C _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__575__C _260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_402_ _070_ _127_ _128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__715__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__586__B _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__648__A3 _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__673__C _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_650_ _312_ _320_ _321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_581_ _107_ _261_ _263_ _264_ _147_ _043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_633_ _306_ _307_ _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_702_ _028_ clknet_3_6__leaf_wb_clk_i lfsr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__578__C _260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_495_ lfsr\[4\] _197_ _198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_564_ counter\[3\] _111_ _235_ counter\[0\] _251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_26_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__439__A1 _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__611__A1 _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_616_ _292_ _294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_547_ _236_ _237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_478_ _176_ _179_ _184_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_401_ _064_ _072_ _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__428__I _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__597__B _277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__705__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__728__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_580_ _107_ _261_ _248_ _264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__436__I _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__484__A2 _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_632_ _083_ _124_ _168_ _307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_701_ _027_ clknet_3_7__leaf_wb_clk_i lfsr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_563_ counter\[4\] _250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_494_ _196_ _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_42_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_615_ _292_ _290_ _293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_546_ _177_ _227_ _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_477_ _180_ _182_ _183_ _184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_400_ _077_ _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_529_ lfsr\[15\] _186_ _222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_47_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__542__I _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__362__I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_700_ _026_ clknet_3_7__leaf_wb_clk_i lfsr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_631_ _105_ _305_ _306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_562_ _108_ _244_ _247_ _249_ _147_ _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_493_ _195_ _196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__718__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_476_ _150_ _183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_614_ counter\[13\] _292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_545_ counter\[1\] _235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__690__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_459_ _167_ _165_ _169_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_528_ lfsr\[14\] _203_ _221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__520__A2 _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_630_ _229_ _231_ _305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_561_ _108_ _244_ _248_ _249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_492_ _085_ _086_ _087_ _195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_1_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__412__B _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__638__I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_3_1__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_613_ _173_ _291_ _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_475_ _181_ _182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_544_ _224_ _229_ _233_ _234_ _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_26_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_527_ _185_ _219_ _220_ _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__708__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_458_ _167_ _165_ _168_ _169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_389_ _114_ counter\[3\] counter\[1\] _115_ _116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_10_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__680__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_12_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__502__C _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_560_ _238_ _248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_491_ _151_ _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_689_ _015_ clknet_3_5__leaf_wb_clk_i m_clkdiv\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_612_ _287_ _289_ _290_ _288_ _291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_543_ _224_ _229_ _151_ _234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_474_ _088_ _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__474__I _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__514__A1 _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_526_ lfsr\[13\] _209_ _188_ _220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_388_ clkdiv\[1\] _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_457_ _150_ _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_509_ _206_ _207_ _146_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__482__I _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_3_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_26_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__693__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_490_ _190_ _192_ _193_ _189_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_688_ _014_ clknet_3_4__leaf_wb_clk_i m_clkdiv\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_473_ lfsr\[0\] _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_611_ _236_ _289_ _290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_542_ _232_ _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__532__A2 _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__523__A2 _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__731__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_456_ m_clkdiv\[6\] _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_525_ _218_ lfsr\[14\] _219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_387_ _109_ _114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__671__A1 _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_508_ lfsr\[9\] _186_ _207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_439_ _152_ _153_ _154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__635__A1 _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_26_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__626__A1 _277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_31_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_687_ _013_ clknet_3_5__leaf_wb_clk_i m_clkdiv\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_610_ _288_ _287_ _277_ _289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_472_ _178_ _179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_541_ _228_ _231_ _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__683__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__540__B _230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_455_ _165_ _166_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_386_ _081_ counter\[7\] _111_ _112_ _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_524_ _180_ _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__450__B _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_507_ lfsr\[8\] _203_ _206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__721__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_438_ m_clkdiv\[1\] m_clkdiv\[0\] m_clkdiv\[2\] _153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_23_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_369_ clkdiv\[6\] _093_ _094_ _082_ _095_ _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_686_ _012_ clknet_3_5__leaf_wb_clk_i m_clkdiv\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__363__B _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_540_ _097_ _102_ _117_ _230_ _231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_471_ _177_ _178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_669_ _332_ _334_ _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_523_ _214_ _197_ _217_ _213_ _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_385_ clkdiv\[2\] _112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_454_ m_clkdiv\[5\] _161_ _162_ _166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_18_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_506_ _194_ _204_ _205_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_437_ _151_ _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_368_ clkdiv\[4\] counter\[4\] _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__696__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__711__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__617__A3 _273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__734__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_685_ _011_ clknet_3_5__leaf_wb_clk_i m_clkdiv\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__462__A1 _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__517__A2 _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_470_ _088_ _177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_668_ _152_ _333_ _334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_599_ _276_ _278_ _280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_737_ _063_ clknet_3_6__leaf_wb_clk_i net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_453_ _164_ _165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_522_ _196_ _216_ _217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_384_ counter\[2\] _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__665__A1 _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__408__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_505_ lfsr\[8\] _192_ _205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_436_ _150_ _151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_367_ counter\[1\] _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_clkbuf_3_6__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_419_ _130_ _138_ _141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__647__B _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__557__B _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__686__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_684_ _010_ clknet_3_5__leaf_wb_clk_i m_clkdiv\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__701__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_736_ _062_ clknet_3_6__leaf_wb_clk_i r_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_667_ _066_ _071_ _177_ _333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_598_ _246_ _278_ _275_ _279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__724__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_16_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_452_ m_clkdiv\[5\] _161_ _164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_383_ clkdiv\[7\] _107_ _108_ _109_ _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_521_ _180_ lfsr\[13\] _216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput3 net3 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_719_ _045_ clknet_3_1__leaf_wb_clk_i counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_18_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__656__A2 _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_435_ net2 _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_504_ lfsr\[7\] _203_ _204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__592__B2 _273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_366_ counter\[6\] _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_2_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__562__C _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_418_ _135_ _140_ _139_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_349_ _065_ _064_ _076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_46_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_683_ _009_ clknet_3_5__leaf_wb_clk_i m_clkdiv\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__676__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_735_ _061_ clknet_3_6__leaf_wb_clk_i r_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_666_ _071_ _178_ _066_ _332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_597_ _275_ _276_ _277_ _278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__699__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_520_ _214_ _185_ _215_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_382_ clkdiv\[3\] _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_451_ _161_ _163_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_33_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput4 net4 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__600__I _157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_718_ _044_ clknet_3_0__leaf_wb_clk_i counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_649_ _079_ _316_ _103_ _308_ _320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__714__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_503_ _195_ _203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_365_ counter\[15\] counter\[14\] counter\[13\] counter\[12\] _092_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_434_ m_clkdiv\[2\] _148_ _149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__737__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_417_ _119_ _121_ _125_ _129_ _136_ _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_348_ _072_ _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_682_ _008_ clknet_3_4__leaf_wb_clk_i m_clkdiv\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_734_ _060_ clknet_3_6__leaf_wb_clk_i r_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_665_ _213_ _331_ _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_596_ _090_ _277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__668__A1 _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_450_ m_clkdiv\[4\] _158_ _162_ _163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_381_ counter\[3\] _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xoutput5 net5 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__581__C _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_717_ _043_ clknet_3_1__leaf_wb_clk_i counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_648_ _316_ _103_ _232_ _308_ _319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_41_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_579_ counter\[7\] _257_ _263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_502_ _200_ _192_ _202_ _189_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_433_ _147_ _086_ _148_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_364_ counter\[11\] counter\[10\] counter\[9\] counter\[8\] _091_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__689__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_416_ _135_ _139_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_347_ _070_ _072_ _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_11_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__704__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__727__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_681_ _007_ clknet_3_5__leaf_wb_clk_i m_clkdiv\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_664_ _071_ _196_ _331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_595_ _271_ _267_ _276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_733_ _059_ clknet_3_3__leaf_wb_clk_i clkdiv\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__524__I _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_380_ counter\[7\] _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xoutput6 net6 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_716_ _042_ clknet_3_0__leaf_wb_clk_i counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_647_ _317_ _318_ _173_ _055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_578_ _093_ _258_ _262_ _260_ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
.ends

