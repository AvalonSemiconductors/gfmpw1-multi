magic
tech gf180mcuD
magscale 1 5
timestamp 1702247549
<< obsm1 >>
rect 672 1538 24304 28545
<< metal2 >>
rect 1792 29600 1848 30000
rect 2576 29600 2632 30000
rect 3360 29600 3416 30000
rect 4144 29600 4200 30000
rect 4928 29600 4984 30000
rect 5712 29600 5768 30000
rect 6496 29600 6552 30000
rect 7280 29600 7336 30000
rect 8064 29600 8120 30000
rect 8848 29600 8904 30000
rect 9632 29600 9688 30000
rect 10416 29600 10472 30000
rect 11200 29600 11256 30000
rect 11984 29600 12040 30000
rect 12768 29600 12824 30000
rect 13552 29600 13608 30000
rect 14336 29600 14392 30000
rect 15120 29600 15176 30000
rect 15904 29600 15960 30000
rect 16688 29600 16744 30000
rect 17472 29600 17528 30000
rect 18256 29600 18312 30000
rect 19040 29600 19096 30000
rect 19824 29600 19880 30000
rect 20608 29600 20664 30000
rect 21392 29600 21448 30000
rect 22176 29600 22232 30000
rect 22960 29600 23016 30000
<< obsm2 >>
rect 742 29570 1762 29666
rect 1878 29570 2546 29666
rect 2662 29570 3330 29666
rect 3446 29570 4114 29666
rect 4230 29570 4898 29666
rect 5014 29570 5682 29666
rect 5798 29570 6466 29666
rect 6582 29570 7250 29666
rect 7366 29570 8034 29666
rect 8150 29570 8818 29666
rect 8934 29570 9602 29666
rect 9718 29570 10386 29666
rect 10502 29570 11170 29666
rect 11286 29570 11954 29666
rect 12070 29570 12738 29666
rect 12854 29570 13522 29666
rect 13638 29570 14306 29666
rect 14422 29570 15090 29666
rect 15206 29570 15874 29666
rect 15990 29570 16658 29666
rect 16774 29570 17442 29666
rect 17558 29570 18226 29666
rect 18342 29570 19010 29666
rect 19126 29570 19794 29666
rect 19910 29570 20578 29666
rect 20694 29570 21362 29666
rect 21478 29570 22146 29666
rect 22262 29570 22930 29666
rect 23046 29570 24234 29666
rect 742 1549 24234 29570
<< metal3 >>
rect 24600 28000 25000 28056
rect 24600 25088 25000 25144
rect 0 24864 400 24920
rect 24600 22176 25000 22232
rect 24600 19264 25000 19320
rect 24600 16352 25000 16408
rect 0 14896 400 14952
rect 24600 13440 25000 13496
rect 24600 10528 25000 10584
rect 24600 7616 25000 7672
rect 0 4928 400 4984
rect 24600 4704 25000 4760
rect 24600 1792 25000 1848
<< obsm3 >>
rect 400 28086 24600 28546
rect 400 27970 24570 28086
rect 400 25174 24600 27970
rect 400 25058 24570 25174
rect 400 24950 24600 25058
rect 430 24834 24600 24950
rect 400 22262 24600 24834
rect 400 22146 24570 22262
rect 400 19350 24600 22146
rect 400 19234 24570 19350
rect 400 16438 24600 19234
rect 400 16322 24570 16438
rect 400 14982 24600 16322
rect 430 14866 24600 14982
rect 400 13526 24600 14866
rect 400 13410 24570 13526
rect 400 10614 24600 13410
rect 400 10498 24570 10614
rect 400 7702 24600 10498
rect 400 7586 24570 7702
rect 400 5014 24600 7586
rect 430 4898 24600 5014
rect 400 4790 24600 4898
rect 400 4674 24570 4790
rect 400 1878 24600 4674
rect 400 1762 24570 1878
rect 400 1554 24600 1762
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
<< obsm4 >>
rect 4382 2585 9874 27543
rect 10094 2585 17554 27543
rect 17774 2585 22218 27543
<< labels >>
rlabel metal3 s 24600 25088 25000 25144 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 24600 28000 25000 28056 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 24600 1792 25000 1848 6 io_in_1[0]
port 3 nsew signal input
rlabel metal3 s 24600 4704 25000 4760 6 io_in_1[1]
port 4 nsew signal input
rlabel metal3 s 24600 7616 25000 7672 6 io_in_1[2]
port 5 nsew signal input
rlabel metal3 s 24600 10528 25000 10584 6 io_in_1[3]
port 6 nsew signal input
rlabel metal3 s 24600 13440 25000 13496 6 io_in_1[4]
port 7 nsew signal input
rlabel metal3 s 24600 16352 25000 16408 6 io_in_1[5]
port 8 nsew signal input
rlabel metal3 s 24600 19264 25000 19320 6 io_in_1[6]
port 9 nsew signal input
rlabel metal3 s 24600 22176 25000 22232 6 io_in_1[7]
port 10 nsew signal input
rlabel metal3 s 0 24864 400 24920 6 io_in_2
port 11 nsew signal input
rlabel metal2 s 1792 29600 1848 30000 6 io_out[0]
port 12 nsew signal output
rlabel metal2 s 9632 29600 9688 30000 6 io_out[10]
port 13 nsew signal output
rlabel metal2 s 10416 29600 10472 30000 6 io_out[11]
port 14 nsew signal output
rlabel metal2 s 11200 29600 11256 30000 6 io_out[12]
port 15 nsew signal output
rlabel metal2 s 11984 29600 12040 30000 6 io_out[13]
port 16 nsew signal output
rlabel metal2 s 12768 29600 12824 30000 6 io_out[14]
port 17 nsew signal output
rlabel metal2 s 13552 29600 13608 30000 6 io_out[15]
port 18 nsew signal output
rlabel metal2 s 14336 29600 14392 30000 6 io_out[16]
port 19 nsew signal output
rlabel metal2 s 15120 29600 15176 30000 6 io_out[17]
port 20 nsew signal output
rlabel metal2 s 15904 29600 15960 30000 6 io_out[18]
port 21 nsew signal output
rlabel metal2 s 16688 29600 16744 30000 6 io_out[19]
port 22 nsew signal output
rlabel metal2 s 2576 29600 2632 30000 6 io_out[1]
port 23 nsew signal output
rlabel metal2 s 17472 29600 17528 30000 6 io_out[20]
port 24 nsew signal output
rlabel metal2 s 18256 29600 18312 30000 6 io_out[21]
port 25 nsew signal output
rlabel metal2 s 19040 29600 19096 30000 6 io_out[22]
port 26 nsew signal output
rlabel metal2 s 19824 29600 19880 30000 6 io_out[23]
port 27 nsew signal output
rlabel metal2 s 20608 29600 20664 30000 6 io_out[24]
port 28 nsew signal output
rlabel metal2 s 21392 29600 21448 30000 6 io_out[25]
port 29 nsew signal output
rlabel metal2 s 22176 29600 22232 30000 6 io_out[26]
port 30 nsew signal output
rlabel metal2 s 22960 29600 23016 30000 6 io_out[27]
port 31 nsew signal output
rlabel metal2 s 3360 29600 3416 30000 6 io_out[2]
port 32 nsew signal output
rlabel metal2 s 4144 29600 4200 30000 6 io_out[3]
port 33 nsew signal output
rlabel metal2 s 4928 29600 4984 30000 6 io_out[4]
port 34 nsew signal output
rlabel metal2 s 5712 29600 5768 30000 6 io_out[5]
port 35 nsew signal output
rlabel metal2 s 6496 29600 6552 30000 6 io_out[6]
port 36 nsew signal output
rlabel metal2 s 7280 29600 7336 30000 6 io_out[7]
port 37 nsew signal output
rlabel metal2 s 8064 29600 8120 30000 6 io_out[8]
port 38 nsew signal output
rlabel metal2 s 8848 29600 8904 30000 6 io_out[9]
port 39 nsew signal output
rlabel metal3 s 0 14896 400 14952 6 rst_n
port 40 nsew signal input
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 42 nsew ground bidirectional
rlabel metal3 s 0 4928 400 4984 6 wb_clk_i
port 43 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 25000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2748630
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_sn76489/runs/23_12_10_23_29/results/signoff/wrapped_sn76489.magic.gds
string GDS_START 402272
<< end >>

