magic
tech gf180mcuD
magscale 1 5
timestamp 1753965646
<< nwell >>
rect 629 1525 19363 18467
<< obsm1 >>
rect 672 1538 19400 18454
<< metal2 >>
rect 1568 19600 1624 20000
rect 2128 19600 2184 20000
rect 2688 19600 2744 20000
rect 3248 19600 3304 20000
rect 3808 19600 3864 20000
rect 4368 19600 4424 20000
rect 4928 19600 4984 20000
rect 5488 19600 5544 20000
rect 6048 19600 6104 20000
rect 6608 19600 6664 20000
rect 7168 19600 7224 20000
rect 7728 19600 7784 20000
rect 8288 19600 8344 20000
rect 8848 19600 8904 20000
rect 9408 19600 9464 20000
rect 9968 19600 10024 20000
rect 10528 19600 10584 20000
rect 11088 19600 11144 20000
rect 11648 19600 11704 20000
rect 12208 19600 12264 20000
rect 12768 19600 12824 20000
rect 13328 19600 13384 20000
rect 13888 19600 13944 20000
rect 14448 19600 14504 20000
rect 15008 19600 15064 20000
rect 15568 19600 15624 20000
rect 16128 19600 16184 20000
rect 16688 19600 16744 20000
rect 17248 19600 17304 20000
rect 17808 19600 17864 20000
rect 18368 19600 18424 20000
rect 560 0 616 400
rect 1456 0 1512 400
rect 2352 0 2408 400
rect 3248 0 3304 400
rect 4144 0 4200 400
rect 5040 0 5096 400
rect 5936 0 5992 400
rect 6832 0 6888 400
rect 7728 0 7784 400
rect 8624 0 8680 400
rect 9520 0 9576 400
rect 10416 0 10472 400
rect 11312 0 11368 400
rect 12208 0 12264 400
rect 13104 0 13160 400
rect 14000 0 14056 400
rect 14896 0 14952 400
rect 15792 0 15848 400
rect 16688 0 16744 400
rect 17584 0 17640 400
rect 18480 0 18536 400
rect 19376 0 19432 400
<< obsm2 >>
rect 574 19570 1538 19642
rect 1654 19570 2098 19642
rect 2214 19570 2658 19642
rect 2774 19570 3218 19642
rect 3334 19570 3778 19642
rect 3894 19570 4338 19642
rect 4454 19570 4898 19642
rect 5014 19570 5458 19642
rect 5574 19570 6018 19642
rect 6134 19570 6578 19642
rect 6694 19570 7138 19642
rect 7254 19570 7698 19642
rect 7814 19570 8258 19642
rect 8374 19570 8818 19642
rect 8934 19570 9378 19642
rect 9494 19570 9938 19642
rect 10054 19570 10498 19642
rect 10614 19570 11058 19642
rect 11174 19570 11618 19642
rect 11734 19570 12178 19642
rect 12294 19570 12738 19642
rect 12854 19570 13298 19642
rect 13414 19570 13858 19642
rect 13974 19570 14418 19642
rect 14534 19570 14978 19642
rect 15094 19570 15538 19642
rect 15654 19570 16098 19642
rect 16214 19570 16658 19642
rect 16774 19570 17218 19642
rect 17334 19570 17778 19642
rect 17894 19570 18338 19642
rect 18454 19570 19530 19642
rect 574 430 19530 19570
rect 646 400 1426 430
rect 1542 400 2322 430
rect 2438 400 3218 430
rect 3334 400 4114 430
rect 4230 400 5010 430
rect 5126 400 5906 430
rect 6022 400 6802 430
rect 6918 400 7698 430
rect 7814 400 8594 430
rect 8710 400 9490 430
rect 9606 400 10386 430
rect 10502 400 11282 430
rect 11398 400 12178 430
rect 12294 400 13074 430
rect 13190 400 13970 430
rect 14086 400 14866 430
rect 14982 400 15762 430
rect 15878 400 16658 430
rect 16774 400 17554 430
rect 17670 400 18450 430
rect 18566 400 19346 430
rect 19462 400 19530 430
<< metal3 >>
rect 19600 18704 20000 18760
rect 19600 17248 20000 17304
rect 19600 15792 20000 15848
rect 19600 14336 20000 14392
rect 19600 12880 20000 12936
rect 19600 11424 20000 11480
rect 19600 9968 20000 10024
rect 19600 8512 20000 8568
rect 19600 7056 20000 7112
rect 19600 5600 20000 5656
rect 19600 4144 20000 4200
rect 19600 2688 20000 2744
rect 19600 1232 20000 1288
<< obsm3 >>
rect 569 18674 19570 18746
rect 569 17334 19642 18674
rect 569 17218 19570 17334
rect 569 15878 19642 17218
rect 569 15762 19570 15878
rect 569 14422 19642 15762
rect 569 14306 19570 14422
rect 569 12966 19642 14306
rect 569 12850 19570 12966
rect 569 11510 19642 12850
rect 569 11394 19570 11510
rect 569 10054 19642 11394
rect 569 9938 19570 10054
rect 569 8598 19642 9938
rect 569 8482 19570 8598
rect 569 7142 19642 8482
rect 569 7026 19570 7142
rect 569 5686 19642 7026
rect 569 5570 19570 5686
rect 569 4230 19642 5570
rect 569 4114 19570 4230
rect 569 2774 19642 4114
rect 569 2658 19570 2774
rect 569 1318 19642 2658
rect 569 1202 19570 1318
rect 569 406 19642 1202
<< metal4 >>
rect 2923 1538 3083 18454
rect 5254 1538 5414 18454
rect 7585 1538 7745 18454
rect 9916 1538 10076 18454
rect 12247 1538 12407 18454
rect 14578 1538 14738 18454
rect 16909 1538 17069 18454
rect 19240 1538 19400 18454
<< obsm4 >>
rect 5446 6337 7555 17687
rect 7775 6337 9886 17687
rect 10106 6337 12217 17687
rect 12437 6337 14548 17687
rect 14768 6337 16879 17687
rect 17099 6337 18858 17687
<< labels >>
rlabel metal3 s 19600 15792 20000 15848 6 SDI
port 1 nsew signal input
rlabel metal3 s 19600 1232 20000 1288 6 clk_i
port 2 nsew signal input
rlabel metal3 s 19600 18704 20000 18760 6 custom_setting
port 3 nsew signal input
rlabel metal3 s 19600 4144 20000 4200 6 io_in[0]
port 4 nsew signal input
rlabel metal3 s 19600 5600 20000 5656 6 io_in[1]
port 5 nsew signal input
rlabel metal3 s 19600 7056 20000 7112 6 io_in[2]
port 6 nsew signal input
rlabel metal3 s 19600 8512 20000 8568 6 io_in[3]
port 7 nsew signal input
rlabel metal3 s 19600 9968 20000 10024 6 io_in[4]
port 8 nsew signal input
rlabel metal3 s 19600 11424 20000 11480 6 io_in[5]
port 9 nsew signal input
rlabel metal3 s 19600 12880 20000 12936 6 io_in[6]
port 10 nsew signal input
rlabel metal3 s 19600 14336 20000 14392 6 io_in[7]
port 11 nsew signal input
rlabel metal2 s 1568 19600 1624 20000 6 io_out[0]
port 12 nsew signal output
rlabel metal2 s 7168 19600 7224 20000 6 io_out[10]
port 13 nsew signal output
rlabel metal2 s 7728 19600 7784 20000 6 io_out[11]
port 14 nsew signal output
rlabel metal2 s 8288 19600 8344 20000 6 io_out[12]
port 15 nsew signal output
rlabel metal2 s 8848 19600 8904 20000 6 io_out[13]
port 16 nsew signal output
rlabel metal2 s 9408 19600 9464 20000 6 io_out[14]
port 17 nsew signal output
rlabel metal2 s 9968 19600 10024 20000 6 io_out[15]
port 18 nsew signal output
rlabel metal2 s 10528 19600 10584 20000 6 io_out[16]
port 19 nsew signal output
rlabel metal2 s 11088 19600 11144 20000 6 io_out[17]
port 20 nsew signal output
rlabel metal2 s 11648 19600 11704 20000 6 io_out[18]
port 21 nsew signal output
rlabel metal2 s 12208 19600 12264 20000 6 io_out[19]
port 22 nsew signal output
rlabel metal2 s 2128 19600 2184 20000 6 io_out[1]
port 23 nsew signal output
rlabel metal2 s 12768 19600 12824 20000 6 io_out[20]
port 24 nsew signal output
rlabel metal2 s 13328 19600 13384 20000 6 io_out[21]
port 25 nsew signal output
rlabel metal2 s 13888 19600 13944 20000 6 io_out[22]
port 26 nsew signal output
rlabel metal2 s 14448 19600 14504 20000 6 io_out[23]
port 27 nsew signal output
rlabel metal2 s 15008 19600 15064 20000 6 io_out[24]
port 28 nsew signal output
rlabel metal2 s 15568 19600 15624 20000 6 io_out[25]
port 29 nsew signal output
rlabel metal2 s 16128 19600 16184 20000 6 io_out[26]
port 30 nsew signal output
rlabel metal2 s 16688 19600 16744 20000 6 io_out[27]
port 31 nsew signal output
rlabel metal2 s 17248 19600 17304 20000 6 io_out[28]
port 32 nsew signal output
rlabel metal2 s 17808 19600 17864 20000 6 io_out[29]
port 33 nsew signal output
rlabel metal2 s 2688 19600 2744 20000 6 io_out[2]
port 34 nsew signal output
rlabel metal2 s 18368 19600 18424 20000 6 io_out[30]
port 35 nsew signal output
rlabel metal2 s 3248 19600 3304 20000 6 io_out[3]
port 36 nsew signal output
rlabel metal2 s 3808 19600 3864 20000 6 io_out[4]
port 37 nsew signal output
rlabel metal2 s 4368 19600 4424 20000 6 io_out[5]
port 38 nsew signal output
rlabel metal2 s 4928 19600 4984 20000 6 io_out[6]
port 39 nsew signal output
rlabel metal2 s 5488 19600 5544 20000 6 io_out[7]
port 40 nsew signal output
rlabel metal2 s 6048 19600 6104 20000 6 io_out[8]
port 41 nsew signal output
rlabel metal2 s 6608 19600 6664 20000 6 io_out[9]
port 42 nsew signal output
rlabel metal3 s 19600 2688 20000 2744 6 rst_n
port 43 nsew signal input
rlabel metal2 s 560 0 616 400 6 sram_addr[0]
port 44 nsew signal output
rlabel metal2 s 1456 0 1512 400 6 sram_addr[1]
port 45 nsew signal output
rlabel metal2 s 2352 0 2408 400 6 sram_addr[2]
port 46 nsew signal output
rlabel metal2 s 3248 0 3304 400 6 sram_addr[3]
port 47 nsew signal output
rlabel metal2 s 4144 0 4200 400 6 sram_addr[4]
port 48 nsew signal output
rlabel metal2 s 5040 0 5096 400 6 sram_addr[5]
port 49 nsew signal output
rlabel metal3 s 19600 17248 20000 17304 6 sram_gwe
port 50 nsew signal output
rlabel metal2 s 5936 0 5992 400 6 sram_in[0]
port 51 nsew signal output
rlabel metal2 s 6832 0 6888 400 6 sram_in[1]
port 52 nsew signal output
rlabel metal2 s 7728 0 7784 400 6 sram_in[2]
port 53 nsew signal output
rlabel metal2 s 8624 0 8680 400 6 sram_in[3]
port 54 nsew signal output
rlabel metal2 s 9520 0 9576 400 6 sram_in[4]
port 55 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 sram_in[5]
port 56 nsew signal output
rlabel metal2 s 11312 0 11368 400 6 sram_in[6]
port 57 nsew signal output
rlabel metal2 s 12208 0 12264 400 6 sram_in[7]
port 58 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 sram_out[0]
port 59 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 sram_out[1]
port 60 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 sram_out[2]
port 61 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 sram_out[3]
port 62 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 sram_out[4]
port 63 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 sram_out[5]
port 64 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 sram_out[6]
port 65 nsew signal input
rlabel metal2 s 19376 0 19432 400 6 sram_out[7]
port 66 nsew signal input
rlabel metal4 s 2923 1538 3083 18454 6 vdd
port 67 nsew power bidirectional
rlabel metal4 s 7585 1538 7745 18454 6 vdd
port 67 nsew power bidirectional
rlabel metal4 s 12247 1538 12407 18454 6 vdd
port 67 nsew power bidirectional
rlabel metal4 s 16909 1538 17069 18454 6 vdd
port 67 nsew power bidirectional
rlabel metal4 s 5254 1538 5414 18454 6 vss
port 68 nsew ground bidirectional
rlabel metal4 s 9916 1538 10076 18454 6 vss
port 68 nsew ground bidirectional
rlabel metal4 s 14578 1538 14738 18454 6 vss
port 68 nsew ground bidirectional
rlabel metal4 s 19240 1538 19400 18454 6 vss
port 68 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1391206
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/wrapped_mc14500/runs/25_07_31_14_39/results/signoff/wrapped_mc14500.magic.gds
string GDS_START 198350
<< end >>

