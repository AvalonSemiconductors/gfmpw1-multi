module ue1 (clk,
    io_oeb,
    rst_n,
    vdd,
    vss,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst_n;
 inout vdd;
 inout vss;
 input [4:0] io_in;
 output [9:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire \main.CAR ;
 wire \main.GATES_1.input1 ;
 wire \main.GATES_100.input1 ;
 wire \main.GATES_100.input2 ;
 wire \main.GATES_102.input1 ;
 wire \main.GATES_102.input2 ;
 wire \main.GATES_102.input3 ;
 wire \main.GATES_103.input2 ;
 wire \main.GATES_105.input3 ;
 wire \main.GATES_106.input2 ;
 wire \main.GATES_107.input2 ;
 wire \main.GATES_108.input1 ;
 wire \main.GATES_109.input1 ;
 wire \main.GATES_109.input2 ;
 wire \main.GATES_11.input2 ;
 wire \main.GATES_110.input1 ;
 wire \main.GATES_111.input2 ;
 wire \main.GATES_113.input1 ;
 wire \main.GATES_114.input2 ;
 wire \main.GATES_115.input2 ;
 wire \main.GATES_116.input1 ;
 wire \main.GATES_116.input3 ;
 wire \main.GATES_119.result ;
 wire \main.GATES_124.input2 ;
 wire \main.GATES_125.input2 ;
 wire \main.GATES_127.result ;
 wire \main.GATES_132.input1 ;
 wire \main.GATES_15.input3 ;
 wire \main.GATES_16.input1 ;
 wire \main.GATES_18.result ;
 wire \main.GATES_19.input1 ;
 wire \main.GATES_20.result ;
 wire \main.GATES_26.input3 ;
 wire \main.GATES_29.input3 ;
 wire \main.GATES_46.input3 ;
 wire \main.GATES_65.result ;
 wire \main.GATES_8.result ;
 wire \main.NOPF ;
 wire \main.WRITE ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__110__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clk));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__111__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_094_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__123__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clk));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__127__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_002_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__139__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_010_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__146__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_002_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__158__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\main.GATES_1.input1 ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__164__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_010_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__171__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\main.GATES_1.input1 ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__175__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\main.GATES_1.input1 ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__191__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\main.GATES_1.input1 ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__194__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_058_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__194__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_094_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__219__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_002_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__223__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_010_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__226__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_058_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__227__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_094_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__231__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_002_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__231__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_058_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__238__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_094_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__241__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_058_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__244__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\main.GATES_1.input1 ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input1_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in[0]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input2_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in[1]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input3_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in[2]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input4_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in[3]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input5_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in[4]));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input6_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(rst_n));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_11_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_11_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_14_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_14_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_1_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_20_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_145 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_20_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_20_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_71 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_4_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_4_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_7_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_7_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_7_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_7_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Left_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Left_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Left_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Left_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Left_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Left_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Left_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Left_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Left_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Left_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Left_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Left_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Left_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Left_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Left_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Left_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Left_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Left_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Left_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Left_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Left_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Left_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _102_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net6),
    .Y(_088_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _103_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_089_),
    .A(_088_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _104_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_089_),
    .Y(_090_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _105_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_091_),
    .B(\main.GATES_109.input2 ),
    .A(\main.GATES_109.input1 ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _106_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_090_),
    .B(\main.GATES_106.input2 ),
    .C(_091_),
    .Y(_092_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _107_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_092_),
    .Y(\main.GATES_109.input1 ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _108_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_090_),
    .B(\main.GATES_107.input2 ),
    .C(\main.GATES_115.input2 ),
    .Y(_093_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _109_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_093_),
    .Y(\main.GATES_102.input2 ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _110_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_094_),
    .B(net6),
    .A(clk));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _111_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_094_),
    .Y(_095_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _112_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\main.GATES_15.input3 ),
    .A(\main.GATES_127.result ),
    .Y(_096_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _113_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_097_),
    .B(_096_),
    .A(_095_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _114_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_102.input1 ),
    .B(_097_),
    .A(\main.GATES_116.input1 ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _115_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_102.input3 ),
    .Y(_098_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _116_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_090_),
    .B(_098_),
    .C(\main.GATES_20.result ),
    .Y(_099_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _117_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_099_),
    .Y(\main.GATES_116.input3 ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _118_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_100_),
    .A(\main.GATES_11.input2 ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _119_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_101_),
    .A(\main.GATES_124.input2 ));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _120_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net6),
    .B(_100_),
    .C(_101_),
    .Y(_000_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _121_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_000_),
    .Y(_001_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _122_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_001_),
    .Y(_002_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _123_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(net6),
    .A(clk),
    .Y(_003_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _124_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_003_),
    .Y(_004_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _125_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_005_),
    .B(\main.GATES_26.input3 ),
    .A(\main.GATES_124.input2 ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _126_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_006_),
    .B(_005_),
    .A(_004_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _127_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_006_),
    .A(_002_),
    .Y(_007_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _128_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_007_),
    .Y(\main.GATES_11.input2 ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _129_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_089_),
    .B(\main.GATES_102.input1 ),
    .C(\main.GATES_127.result ),
    .Y(_008_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _130_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_008_),
    .Y(\main.GATES_116.input1 ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _131_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_100_),
    .Y(_009_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _132_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_003_),
    .A(_009_),
    .Y(_010_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _133_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\main.GATES_102.input2 ),
    .A(\main.GATES_102.input1 ),
    .Y(_011_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _134_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_012_),
    .B(_011_),
    .A(\main.GATES_116.input3 ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _135_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_116.input3 ),
    .Y(_013_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _136_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_013_),
    .B(\main.GATES_102.input2 ),
    .C(\main.GATES_116.input1 ),
    .Y(_014_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _137_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_014_),
    .A(_012_),
    .Y(_015_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _138_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_015_),
    .A(\main.GATES_109.input1 ),
    .Y(_016_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _139_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(net7),
    .B(_016_),
    .A(_010_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _140_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.WRITE ),
    .A(net7));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _141_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\main.GATES_29.input3 ),
    .A(\main.GATES_115.input2 ),
    .Y(_017_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _142_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_018_),
    .B(_017_),
    .A(_095_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _143_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_107.input2 ),
    .B(_018_),
    .A(\main.GATES_102.input2 ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _144_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\main.GATES_107.input2 ),
    .A(\main.GATES_102.input1 ),
    .Y(_019_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _145_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_020_),
    .B(_019_),
    .A(_013_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _146_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_020_),
    .A(_002_),
    .Y(_021_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _147_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_021_),
    .Y(\main.GATES_114.input2 ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _148_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_088_),
    .Y(_022_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _149_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_100.input1 ),
    .Y(_023_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _150_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_024_),
    .A(_022_),
    .B(net2),
    .C(_023_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _151_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_15.input3 ),
    .B(_024_),
    .A(_097_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _152_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_096_),
    .A(_004_),
    .Y(_025_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _153_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_025_),
    .Y(\main.GATES_127.result ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _154_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_1.input1 ),
    .B(\main.GATES_108.input1 ),
    .A(\main.GATES_119.result ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _155_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_108.input1 ),
    .B(_004_),
    .A(\main.GATES_113.input1 ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _156_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_026_),
    .A(\main.GATES_108.input1 ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _157_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_095_),
    .Y(_027_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _158_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_119.result ),
    .C(\main.GATES_1.input1 ),
    .B(_027_),
    .A(_026_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _159_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_102.input3 ),
    .B(\main.GATES_19.input1 ),
    .A(_013_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _160_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_098_),
    .B(\main.GATES_11.input2 ),
    .C(_019_),
    .Y(_028_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _161_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_028_),
    .Y(\main.GATES_100.input2 ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _162_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\main.GATES_116.input1 ),
    .A(\main.GATES_107.input2 ),
    .Y(_029_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _163_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_030_),
    .B(_029_),
    .A(_013_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _164_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_030_),
    .A(_010_),
    .Y(_031_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _165_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_032_),
    .B(\main.GATES_105.input3 ),
    .A(\main.GATES_103.input2 ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _166_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_033_),
    .B(_032_),
    .A(_031_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _167_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_034_),
    .B(\main.GATES_111.input2 ),
    .A(\main.GATES_103.input2 ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _168_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_111.input2 ),
    .C(_090_),
    .B(_034_),
    .A(_033_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _169_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\main.GATES_119.result ),
    .A(_009_),
    .Y(_035_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _170_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_088_),
    .B(net1),
    .C(_012_),
    .D(_035_),
    .Y(_036_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _171_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_009_),
    .B(\main.GATES_1.input1 ),
    .C(_014_),
    .Y(_037_),
    .D(_036_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _172_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_110.input1 ),
    .B(_037_),
    .A(\main.GATES_111.input2 ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _173_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_000_),
    .Y(_038_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _174_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_039_),
    .C(\main.GATES_114.input2 ),
    .B(_030_),
    .A(_038_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _175_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_040_),
    .A(\main.GATES_1.input1 ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _176_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_041_),
    .C(_040_),
    .B(_012_),
    .A(_001_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _177_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_042_),
    .B(_041_),
    .A(_039_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _178_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_043_),
    .A(\main.GATES_110.input1 ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _179_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_011_),
    .A(\main.GATES_102.input3 ),
    .Y(_044_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _180_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_045_),
    .B(_000_),
    .A(_044_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _181_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_046_),
    .B(_029_),
    .A(_098_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _182_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\main.GATES_119.result ),
    .A(_043_),
    .Y(_047_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _183_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_048_),
    .C(_047_),
    .B(_046_),
    .A(_038_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _184_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_048_),
    .A(_040_),
    .B(_043_),
    .C(_045_),
    .Y(_049_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _185_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_098_),
    .A(_011_),
    .B(_019_),
    .C(_029_),
    .Y(_050_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _186_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_051_),
    .B(_050_),
    .A(_038_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _187_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_051_),
    .B(_049_),
    .A(_042_),
    .Y(_052_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _188_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_053_),
    .A(_001_),
    .B(_030_),
    .C(\main.GATES_114.input2 ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _189_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_054_),
    .A(\main.CAR ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _190_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\main.GATES_114.input2 ),
    .A(\main.GATES_110.input1 ),
    .Y(_055_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _191_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_055_),
    .A(\main.GATES_1.input1 ),
    .Y(_056_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _192_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_056_),
    .A(_054_),
    .Y(_057_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _193_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_102.input3 ),
    .B(\main.GATES_102.input2 ),
    .C(\main.GATES_116.input1 ),
    .Y(_058_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _194_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_059_),
    .A(_000_),
    .B(_058_),
    .C(_094_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _195_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_059_),
    .A(\main.GATES_110.input1 ),
    .B(_001_),
    .C(_012_),
    .Y(_060_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _196_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_061_),
    .C(_060_),
    .B(_057_),
    .A(_053_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _197_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_113.input1 ),
    .A(_022_),
    .B(\main.GATES_108.input1 ),
    .C(_052_),
    .D(_061_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _198_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_017_),
    .A(_004_),
    .Y(_062_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _199_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_062_),
    .Y(\main.GATES_115.input2 ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _200_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_063_),
    .A(_088_),
    .B(net3),
    .C(\main.GATES_100.input1 ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _201_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_29.input3 ),
    .B(_063_),
    .A(_018_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _202_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_064_),
    .A(\main.GATES_18.result ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _203_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_18.result ),
    .B(\main.GATES_46.input3 ),
    .C(_095_),
    .Y(_065_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _204_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_065_),
    .A(_022_),
    .B(_064_),
    .C(_023_),
    .Y(_066_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _205_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_066_),
    .Y(\main.GATES_100.input1 ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _206_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_067_),
    .A(\main.GATES_46.input3 ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _207_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_18.result ),
    .C(_027_),
    .B(_067_),
    .A(_064_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _208_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_068_),
    .A(_023_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _209_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_125.input2 ),
    .B(_044_),
    .A(\main.GATES_11.input2 ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _210_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_069_),
    .A(_035_),
    .B(_046_),
    .C(\main.GATES_125.input2 ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _211_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_46.input3 ),
    .C(_065_),
    .B(_069_),
    .A(_068_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _212_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_070_),
    .C(_023_),
    .B(net5),
    .A(_022_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _213_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_070_),
    .A(_006_),
    .Y(_071_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _214_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_071_),
    .Y(\main.GATES_26.input3 ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _215_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_124.input2 ),
    .B(_005_),
    .A(_027_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _216_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_037_),
    .A(_033_),
    .Y(_072_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _217_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_072_),
    .Y(\main.GATES_105.input3 ));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _218_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_103.input2 ),
    .B(_032_),
    .A(_031_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _219_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_014_),
    .A(_002_),
    .Y(_073_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _220_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_073_),
    .Y(\main.GATES_65.result ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _221_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_074_),
    .A(\main.GATES_109.input2 ));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _222_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_075_),
    .A(_074_),
    .B(_037_),
    .C(\main.GATES_106.input2 ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _223_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_076_),
    .B(_020_),
    .A(_010_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _224_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_106.input2 ),
    .B(_076_),
    .A(_075_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _225_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_109.input2 ),
    .B(_076_),
    .A(_075_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _226_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_077_),
    .B(_058_),
    .A(_038_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _227_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_078_),
    .C(_094_),
    .B(_077_),
    .A(_039_));
 gf180mcu_as_sc_mcu7t3v3__mux2_2 _228_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .S(_078_),
    .B(\main.CAR ),
    .A(\main.GATES_132.input1 ),
    .Y(_079_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _229_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_079_),
    .Y(\main.CAR ));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _230_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_080_),
    .A(_040_),
    .B(_054_),
    .C(_055_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _231_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_081_),
    .A(_002_),
    .B(_058_),
    .C(_080_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _232_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_089_),
    .B(\main.GATES_132.input1 ),
    .C(_078_),
    .Y(_082_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _233_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_132.input1 ),
    .C(_082_),
    .B(_081_),
    .A(_078_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _234_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\main.GATES_16.input1 ),
    .A(\main.GATES_100.input1 ),
    .Y(_083_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _235_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_083_),
    .A(\main.GATES_100.input2 ),
    .Y(_084_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _236_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_084_),
    .Y(\main.GATES_16.input1 ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _237_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net4),
    .B(\main.GATES_100.input1 ),
    .C(\main.GATES_19.input1 ),
    .Y(_085_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _238_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_20.result ),
    .B(_094_),
    .C(_085_),
    .Y(_086_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _239_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_086_),
    .Y(\main.GATES_19.input1 ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _240_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.GATES_20.result ),
    .B(\main.GATES_19.input1 ),
    .A(_027_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _241_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_058_),
    .A(_009_),
    .Y(_087_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _242_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_087_),
    .Y(\main.GATES_8.result ));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _243_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(\main.NOPF ),
    .B(\main.GATES_16.input1 ),
    .A(\main.GATES_100.input2 ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _244_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_1.input1 ),
    .Y(net8));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _245_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.WRITE ),
    .Y(net9));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _246_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.CAR ),
    .Y(net10));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _247_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_111.input2 ),
    .Y(net11));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _248_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_8.result ),
    .Y(net12));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _249_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.NOPF ),
    .Y(net13));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _250_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_65.result ),
    .Y(net14));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _251_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_109.input1 ),
    .Y(net15));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _252_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_125.input2 ),
    .Y(net16));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _253_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\main.GATES_100.input1 ),
    .Y(net17));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input1 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in[0]),
    .Y(net1));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in[1]),
    .Y(net2));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input3 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in[2]),
    .Y(net3));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in[3]),
    .Y(net4));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in[4]),
    .Y(net5));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(rst_n),
    .Y(net6));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net10),
    .Y(io_out[2]));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net11),
    .Y(io_out[3]));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net12),
    .Y(io_out[4]));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net13),
    .Y(io_out[5]));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net14),
    .Y(io_out[6]));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net15),
    .Y(io_out[7]));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net16),
    .Y(io_out[8]));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net17),
    .Y(io_out[9]));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net7),
    .Y(io_oeb));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net8),
    .Y(io_out[0]));
 gf180mcu_as_sc_mcu7t3v3__buff_2 output9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net9),
    .Y(io_out[1]));
endmodule
