magic
tech gf180mcuD
magscale 1 10
timestamp 1753967821
<< metal1 >>
rect 1344 42362 44576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 44576 42362
rect 1344 42276 44576 42310
rect 41694 42194 41746 42206
rect 41694 42130 41746 42142
rect 32286 42008 32338 42020
rect 31266 41933 31278 41985
rect 31330 41933 31342 41985
rect 31602 41918 31614 41970
rect 31666 41918 31678 41970
rect 32846 41970 32898 41982
rect 32286 41944 32338 41956
rect 32610 41918 32622 41970
rect 32674 41918 32686 41970
rect 36878 41970 36930 41982
rect 32846 41906 32898 41918
rect 33014 41914 33066 41926
rect 36878 41906 36930 41918
rect 37102 41970 37154 41982
rect 43026 41945 43038 41997
rect 43090 41945 43102 41997
rect 37102 41906 37154 41918
rect 31154 41806 31166 41858
rect 31218 41806 31230 41858
rect 33014 41850 33066 41862
rect 33618 41694 33630 41746
rect 33682 41743 33694 41746
rect 34626 41743 34638 41746
rect 33682 41697 34638 41743
rect 33682 41694 33694 41697
rect 34626 41694 34638 41697
rect 34690 41694 34702 41746
rect 36586 41694 36598 41746
rect 36650 41694 36662 41746
rect 37426 41694 37438 41746
rect 37490 41743 37502 41746
rect 38322 41743 38334 41746
rect 37490 41697 38334 41743
rect 37490 41694 37502 41697
rect 38322 41694 38334 41697
rect 38386 41694 38398 41746
rect 1344 41578 44576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 44576 41578
rect 1344 41492 44576 41526
rect 35422 41410 35474 41422
rect 35422 41346 35474 41358
rect 22978 41246 22990 41298
rect 23042 41246 23054 41298
rect 26450 41246 26462 41298
rect 26514 41246 26526 41298
rect 30930 41246 30942 41298
rect 30994 41246 31006 41298
rect 33282 41246 33294 41298
rect 33346 41246 33358 41298
rect 35970 41246 35982 41298
rect 36034 41246 36046 41298
rect 37426 41246 37438 41298
rect 37490 41246 37502 41298
rect 22542 41186 22594 41198
rect 22542 41122 22594 41134
rect 22654 41186 22706 41198
rect 26014 41186 26066 41198
rect 22654 41122 22706 41134
rect 23090 41090 23102 41142
rect 23154 41090 23166 41142
rect 23314 41134 23326 41186
rect 23378 41134 23390 41186
rect 26014 41122 26066 41134
rect 26238 41186 26290 41198
rect 30158 41186 30210 41198
rect 35758 41186 35810 41198
rect 37662 41186 37714 41198
rect 26238 41122 26290 41134
rect 26562 41090 26574 41142
rect 26626 41090 26638 41142
rect 26898 41134 26910 41186
rect 26962 41134 26974 41186
rect 30158 41122 30210 41134
rect 33394 41119 33406 41171
rect 33458 41119 33470 41171
rect 33618 41134 33630 41186
rect 33682 41134 33694 41186
rect 35758 41122 35810 41134
rect 36082 41119 36094 41171
rect 36146 41119 36158 41171
rect 36418 41134 36430 41186
rect 36482 41134 36494 41186
rect 36978 41134 36990 41186
rect 37042 41134 37054 41186
rect 37314 41119 37326 41171
rect 37378 41119 37390 41171
rect 37662 41122 37714 41134
rect 41358 41130 41410 41142
rect 32846 41074 32898 41086
rect 22250 41022 22262 41074
rect 22314 41022 22326 41074
rect 25722 41022 25734 41074
rect 25786 41022 25798 41074
rect 32846 41010 32898 41022
rect 40518 41074 40570 41086
rect 40786 41078 40798 41130
rect 40850 41078 40862 41130
rect 41010 41078 41022 41130
rect 41074 41078 41086 41130
rect 41234 41078 41246 41130
rect 41298 41078 41310 41130
rect 42018 41106 42030 41158
rect 42082 41106 42094 41158
rect 41358 41066 41410 41078
rect 40518 41010 40570 41022
rect 37998 40962 38050 40974
rect 37998 40898 38050 40910
rect 43374 40962 43426 40974
rect 43374 40898 43426 40910
rect 1344 40794 44576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 44576 40794
rect 1344 40708 44576 40742
rect 23942 40570 23994 40582
rect 23942 40506 23994 40518
rect 32398 40514 32450 40526
rect 28634 40462 28646 40514
rect 28698 40462 28710 40514
rect 32398 40450 32450 40462
rect 33182 40514 33234 40526
rect 33182 40450 33234 40462
rect 37774 40514 37826 40526
rect 20750 40402 20802 40414
rect 20750 40338 20802 40350
rect 23438 40402 23490 40414
rect 24782 40402 24834 40414
rect 23762 40350 23774 40402
rect 23826 40350 23838 40402
rect 23438 40338 23490 40350
rect 24782 40338 24834 40350
rect 25118 40402 25170 40414
rect 25118 40338 25170 40350
rect 27806 40402 27858 40414
rect 27806 40338 27858 40350
rect 28142 40402 28194 40414
rect 28142 40338 28194 40350
rect 28366 40402 28418 40414
rect 28366 40338 28418 40350
rect 29710 40402 29762 40414
rect 33413 40406 33425 40458
rect 33477 40406 33489 40458
rect 37774 40450 37826 40462
rect 29710 40338 29762 40350
rect 34302 40402 34354 40414
rect 34302 40338 34354 40350
rect 35086 40402 35138 40414
rect 38110 40402 38162 40414
rect 35858 40350 35870 40402
rect 35922 40350 35934 40402
rect 35086 40338 35138 40350
rect 38110 40338 38162 40350
rect 38334 40402 38386 40414
rect 39790 40402 39842 40414
rect 38602 40350 38614 40402
rect 38666 40350 38678 40402
rect 38334 40338 38386 40350
rect 39790 40338 39842 40350
rect 40462 40402 40514 40414
rect 40462 40338 40514 40350
rect 40798 40402 40850 40414
rect 40798 40338 40850 40350
rect 43486 40402 43538 40414
rect 43486 40338 43538 40350
rect 24446 40290 24498 40302
rect 29206 40290 29258 40302
rect 40126 40290 40178 40302
rect 21522 40238 21534 40290
rect 21586 40238 21598 40290
rect 25890 40238 25902 40290
rect 25954 40238 25966 40290
rect 30482 40238 30494 40290
rect 30546 40238 30558 40290
rect 41570 40238 41582 40290
rect 41634 40238 41646 40290
rect 24446 40226 24498 40238
rect 29206 40226 29258 40238
rect 40126 40226 40178 40238
rect 39454 40178 39506 40190
rect 39454 40114 39506 40126
rect 1344 40010 44576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 44576 40010
rect 1344 39924 44576 39958
rect 40294 39842 40346 39854
rect 21870 39786 21922 39798
rect 23090 39734 23102 39786
rect 23154 39734 23166 39786
rect 21870 39722 21922 39734
rect 28646 39730 28698 39742
rect 34290 39734 34302 39786
rect 34354 39734 34366 39786
rect 40294 39778 40346 39790
rect 43934 39842 43986 39854
rect 43934 39778 43986 39790
rect 27346 39678 27358 39730
rect 27410 39678 27422 39730
rect 41346 39678 41358 39730
rect 41410 39678 41422 39730
rect 28646 39666 28698 39678
rect 24110 39618 24162 39630
rect 27918 39618 27970 39630
rect 21970 39566 21982 39618
rect 22034 39566 22046 39618
rect 22306 39566 22318 39618
rect 22370 39566 22382 39618
rect 22638 39528 22650 39580
rect 22702 39528 22714 39580
rect 23314 39566 23326 39618
rect 23378 39566 23390 39618
rect 24882 39566 24894 39618
rect 24946 39566 24958 39618
rect 27234 39566 27246 39618
rect 27298 39566 27310 39618
rect 24110 39554 24162 39566
rect 26798 39506 26850 39518
rect 27682 39510 27694 39562
rect 27746 39510 27758 39562
rect 27918 39554 27970 39566
rect 30270 39618 30322 39630
rect 33742 39618 33794 39630
rect 31042 39566 31054 39618
rect 31106 39566 31118 39618
rect 30270 39554 30322 39566
rect 33742 39554 33794 39566
rect 33854 39618 33906 39630
rect 35758 39618 35810 39630
rect 37662 39618 37714 39630
rect 34178 39566 34190 39618
rect 34242 39566 34254 39618
rect 34514 39566 34526 39618
rect 34578 39566 34590 39618
rect 33854 39554 33906 39566
rect 35758 39554 35810 39566
rect 35982 39579 36034 39591
rect 36306 39566 36318 39618
rect 36370 39566 36382 39618
rect 36978 39566 36990 39618
rect 37042 39566 37054 39618
rect 37438 39579 37490 39591
rect 26798 39442 26850 39454
rect 32958 39506 33010 39518
rect 35982 39515 36034 39527
rect 40574 39618 40626 39630
rect 39566 39590 39618 39602
rect 37662 39554 37714 39566
rect 39454 39562 39506 39574
rect 37438 39515 37490 39527
rect 39566 39526 39618 39538
rect 39790 39590 39842 39602
rect 39790 39526 39842 39538
rect 40014 39590 40066 39602
rect 40574 39554 40626 39566
rect 43598 39618 43650 39630
rect 43598 39554 43650 39566
rect 40014 39526 40066 39538
rect 33450 39454 33462 39506
rect 33514 39454 33526 39506
rect 39454 39498 39506 39510
rect 43262 39506 43314 39518
rect 32958 39442 33010 39454
rect 35634 39398 35646 39450
rect 35698 39398 35710 39450
rect 37538 39398 37550 39450
rect 37602 39398 37614 39450
rect 43262 39442 43314 39454
rect 1344 39226 44576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 44576 39226
rect 1344 39140 44576 39174
rect 32398 39058 32450 39070
rect 32398 38994 32450 39006
rect 34974 39058 35026 39070
rect 34974 38994 35026 39006
rect 22430 38946 22482 38958
rect 22990 38946 23042 38958
rect 38110 38946 38162 38958
rect 22430 38882 22482 38894
rect 22822 38890 22874 38902
rect 19742 38834 19794 38846
rect 24602 38894 24614 38946
rect 24666 38894 24678 38946
rect 22990 38882 23042 38894
rect 38110 38882 38162 38894
rect 39454 38869 39506 38881
rect 22822 38826 22874 38838
rect 23202 38782 23214 38834
rect 23266 38782 23278 38834
rect 23426 38810 23438 38862
rect 23490 38810 23502 38862
rect 24110 38834 24162 38846
rect 19742 38770 19794 38782
rect 24110 38770 24162 38782
rect 24334 38834 24386 38846
rect 24334 38770 24386 38782
rect 25118 38834 25170 38846
rect 28702 38834 28754 38846
rect 25890 38782 25902 38834
rect 25954 38782 25966 38834
rect 30370 38809 30382 38861
rect 30434 38809 30446 38861
rect 31726 38834 31778 38846
rect 25118 38770 25170 38782
rect 28702 38770 28754 38782
rect 31726 38770 31778 38782
rect 31950 38834 32002 38846
rect 31950 38770 32002 38782
rect 32062 38834 32114 38846
rect 33406 38834 33458 38846
rect 33114 38782 33126 38834
rect 33178 38782 33190 38834
rect 32062 38770 32114 38782
rect 33406 38770 33458 38782
rect 33630 38834 33682 38846
rect 33630 38770 33682 38782
rect 35310 38834 35362 38846
rect 35310 38770 35362 38782
rect 35422 38834 35474 38846
rect 36194 38782 36206 38834
rect 36258 38782 36270 38834
rect 39554 38838 39566 38890
rect 39618 38838 39630 38890
rect 39790 38862 39842 38874
rect 39454 38805 39506 38817
rect 39790 38798 39842 38810
rect 40014 38862 40066 38874
rect 40014 38798 40066 38810
rect 43710 38834 43762 38846
rect 35422 38770 35474 38782
rect 43710 38770 43762 38782
rect 20514 38670 20526 38722
rect 20578 38670 20590 38722
rect 27794 38670 27806 38722
rect 27858 38670 27870 38722
rect 31434 38670 31446 38722
rect 31498 38670 31510 38722
rect 41010 38670 41022 38722
rect 41074 38670 41086 38722
rect 42914 38670 42926 38722
rect 42978 38670 42990 38722
rect 40294 38610 40346 38622
rect 40294 38546 40346 38558
rect 1344 38442 44576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 44576 38442
rect 1344 38356 44576 38390
rect 43710 38274 43762 38286
rect 21870 38218 21922 38230
rect 29530 38222 29542 38274
rect 29594 38222 29606 38274
rect 31322 38222 31334 38274
rect 31386 38222 31398 38274
rect 34190 38218 34242 38230
rect 24882 38166 24894 38218
rect 24946 38166 24958 38218
rect 26226 38166 26238 38218
rect 26290 38166 26302 38218
rect 20290 38110 20302 38162
rect 20354 38110 20366 38162
rect 21870 38154 21922 38166
rect 31838 38162 31890 38174
rect 43710 38210 43762 38222
rect 34190 38154 34242 38166
rect 40562 38110 40574 38162
rect 40626 38110 40638 38162
rect 31838 38098 31890 38110
rect 22990 38050 23042 38062
rect 20402 37954 20414 38006
rect 20466 37954 20478 38006
rect 20738 37998 20750 38050
rect 20802 37998 20814 38050
rect 21970 37998 21982 38050
rect 22034 37998 22046 38050
rect 22306 37998 22318 38050
rect 22370 37998 22382 38050
rect 22990 37986 23042 37998
rect 23102 38050 23154 38062
rect 23102 37986 23154 37998
rect 23326 38050 23378 38062
rect 23326 37986 23378 37998
rect 23550 38050 23602 38062
rect 24110 38050 24162 38062
rect 23818 37998 23830 38050
rect 23882 37998 23894 38050
rect 23550 37986 23602 37998
rect 24110 37986 24162 37998
rect 24446 38050 24498 38062
rect 25678 38050 25730 38062
rect 27246 38050 27298 38062
rect 24994 37998 25006 38050
rect 25058 37998 25070 38050
rect 26226 37998 26238 38050
rect 26290 37998 26302 38050
rect 26450 37998 26462 38050
rect 26514 37998 26526 38050
rect 26954 37998 26966 38050
rect 27018 37998 27030 38050
rect 24446 37986 24498 37998
rect 25678 37986 25730 37998
rect 27246 37986 27298 37998
rect 27470 38050 27522 38062
rect 27470 37986 27522 37998
rect 27582 38050 27634 38062
rect 27582 37986 27634 37998
rect 29038 38050 29090 38062
rect 29038 37986 29090 37998
rect 29262 38050 29314 38062
rect 29262 37986 29314 37998
rect 30830 38050 30882 38062
rect 30830 37986 30882 37998
rect 31054 38050 31106 38062
rect 31054 37986 31106 37998
rect 32174 38050 32226 38062
rect 37438 38050 37490 38062
rect 34290 37998 34302 38050
rect 34354 37998 34366 38050
rect 34626 37998 34638 38050
rect 34690 37998 34702 38050
rect 36530 37998 36542 38050
rect 36594 37998 36606 38050
rect 32174 37986 32226 37998
rect 37438 37986 37490 37998
rect 38670 38050 38722 38062
rect 38670 37986 38722 37998
rect 41358 38050 41410 38062
rect 42422 38050 42474 38062
rect 41358 37986 41410 37998
rect 41582 38015 41634 38027
rect 41918 38022 41970 38034
rect 41582 37951 41634 37963
rect 37102 37938 37154 37950
rect 41682 37942 41694 37994
rect 41746 37942 41758 37994
rect 41918 37958 41970 37970
rect 42130 37942 42142 37994
rect 42194 37942 42206 37994
rect 42422 37986 42474 37998
rect 42702 38050 42754 38062
rect 42702 37986 42754 37998
rect 43374 38050 43426 38062
rect 43374 37986 43426 37998
rect 22698 37886 22710 37938
rect 22762 37886 22774 37938
rect 37102 37874 37154 37886
rect 36374 37826 36426 37838
rect 36374 37762 36426 37774
rect 43038 37826 43090 37838
rect 43038 37762 43090 37774
rect 1344 37658 44576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 44576 37658
rect 1344 37572 44576 37606
rect 34862 37490 34914 37502
rect 34862 37426 34914 37438
rect 39566 37490 39618 37502
rect 39566 37426 39618 37438
rect 40238 37490 40290 37502
rect 40238 37426 40290 37438
rect 30718 37378 30770 37390
rect 23930 37326 23942 37378
rect 23994 37326 24006 37378
rect 30718 37314 30770 37326
rect 19630 37266 19682 37278
rect 19630 37202 19682 37214
rect 22318 37266 22370 37278
rect 22318 37202 22370 37214
rect 22654 37266 22706 37278
rect 22654 37202 22706 37214
rect 22878 37266 22930 37278
rect 22878 37202 22930 37214
rect 23438 37266 23490 37278
rect 23438 37202 23490 37214
rect 23662 37266 23714 37278
rect 23662 37202 23714 37214
rect 27134 37266 27186 37278
rect 27414 37266 27466 37278
rect 27234 37214 27246 37266
rect 27298 37214 27310 37266
rect 27134 37202 27186 37214
rect 27414 37202 27466 37214
rect 27582 37266 27634 37278
rect 27582 37202 27634 37214
rect 28030 37266 28082 37278
rect 28030 37202 28082 37214
rect 31502 37266 31554 37278
rect 31502 37202 31554 37214
rect 31614 37266 31666 37278
rect 31614 37202 31666 37214
rect 31838 37266 31890 37278
rect 31838 37202 31890 37214
rect 32062 37266 32114 37278
rect 34526 37266 34578 37278
rect 33170 37214 33182 37266
rect 33234 37214 33246 37266
rect 33506 37214 33518 37266
rect 33570 37214 33582 37266
rect 33842 37214 33854 37266
rect 33906 37214 33918 37266
rect 34178 37214 34190 37266
rect 34242 37214 34254 37266
rect 35858 37214 35870 37266
rect 35922 37214 35934 37266
rect 36082 37229 36094 37281
rect 36146 37229 36158 37281
rect 36642 37229 36654 37281
rect 36706 37229 36718 37281
rect 37214 37266 37266 37278
rect 36978 37214 36990 37266
rect 37042 37214 37054 37266
rect 32062 37202 32114 37214
rect 34526 37202 34578 37214
rect 37214 37202 37266 37214
rect 37886 37266 37938 37278
rect 37886 37202 37938 37214
rect 39230 37266 39282 37278
rect 39230 37202 39282 37214
rect 39902 37266 39954 37278
rect 39902 37202 39954 37214
rect 40910 37266 40962 37278
rect 41682 37214 41694 37266
rect 41746 37214 41758 37266
rect 40910 37202 40962 37214
rect 20402 37102 20414 37154
rect 20466 37102 20478 37154
rect 28802 37102 28814 37154
rect 28866 37102 28878 37154
rect 33070 37098 33122 37110
rect 26854 37042 26906 37054
rect 23146 36990 23158 37042
rect 23210 36990 23222 37042
rect 31210 36990 31222 37042
rect 31274 36990 31286 37042
rect 32330 36990 32342 37042
rect 32394 36990 32406 37042
rect 33070 37034 33122 37046
rect 34302 37098 34354 37110
rect 36194 37102 36206 37154
rect 36258 37102 36270 37154
rect 36530 37102 36542 37154
rect 36594 37102 36606 37154
rect 43586 37102 43598 37154
rect 43650 37102 43662 37154
rect 34302 37034 34354 37046
rect 37550 37042 37602 37054
rect 26854 36978 26906 36990
rect 37550 36978 37602 36990
rect 38222 37042 38274 37054
rect 38222 36978 38274 36990
rect 1344 36874 44576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 44576 36874
rect 1344 36788 44576 36822
rect 29934 36706 29986 36718
rect 21758 36650 21810 36662
rect 29934 36642 29986 36654
rect 33730 36598 33742 36650
rect 33794 36598 33806 36650
rect 20290 36542 20302 36594
rect 20354 36542 20366 36594
rect 21758 36586 21810 36598
rect 22138 36542 22150 36594
rect 22202 36542 22214 36594
rect 37986 36542 37998 36594
rect 38050 36542 38062 36594
rect 43138 36542 43150 36594
rect 43202 36542 43214 36594
rect 12126 36482 12178 36494
rect 22430 36482 22482 36494
rect 12126 36418 12178 36430
rect 20402 36415 20414 36467
rect 20466 36415 20478 36467
rect 20626 36430 20638 36482
rect 20690 36430 20702 36482
rect 21410 36430 21422 36482
rect 21474 36430 21486 36482
rect 21634 36430 21646 36482
rect 21698 36430 21710 36482
rect 22430 36418 22482 36430
rect 22654 36482 22706 36494
rect 22654 36418 22706 36430
rect 22766 36482 22818 36494
rect 22766 36418 22818 36430
rect 22990 36482 23042 36494
rect 22990 36418 23042 36430
rect 26910 36482 26962 36494
rect 26910 36418 26962 36430
rect 29038 36482 29090 36494
rect 27774 36374 27786 36426
rect 27838 36374 27850 36426
rect 29038 36418 29090 36430
rect 30270 36482 30322 36494
rect 30830 36482 30882 36494
rect 30538 36430 30550 36482
rect 30602 36430 30614 36482
rect 30270 36418 30322 36430
rect 30830 36418 30882 36430
rect 31054 36482 31106 36494
rect 31950 36482 32002 36494
rect 31658 36430 31670 36482
rect 31722 36430 31734 36482
rect 31054 36418 31106 36430
rect 31950 36418 32002 36430
rect 32174 36482 32226 36494
rect 32174 36418 32226 36430
rect 32958 36482 33010 36494
rect 34134 36482 34186 36494
rect 33506 36430 33518 36482
rect 33570 36430 33582 36482
rect 32958 36418 33010 36430
rect 34134 36418 34186 36430
rect 34414 36482 34466 36494
rect 34862 36482 34914 36494
rect 34514 36430 34526 36482
rect 34578 36430 34590 36482
rect 41022 36454 41074 36466
rect 34414 36418 34466 36430
rect 28030 36370 28082 36382
rect 34682 36374 34694 36426
rect 34746 36374 34758 36426
rect 34862 36418 34914 36430
rect 37202 36402 37214 36454
rect 37266 36402 37278 36454
rect 23258 36318 23270 36370
rect 23322 36318 23334 36370
rect 28030 36306 28082 36318
rect 40518 36370 40570 36382
rect 40786 36374 40798 36426
rect 40850 36374 40862 36426
rect 41022 36390 41074 36402
rect 41246 36454 41298 36466
rect 41246 36390 41298 36402
rect 41358 36426 41410 36438
rect 43810 36402 43822 36454
rect 43874 36402 43886 36454
rect 41358 36362 41410 36374
rect 40518 36306 40570 36318
rect 11790 36258 11842 36270
rect 29374 36258 29426 36270
rect 15362 36206 15374 36258
rect 15426 36255 15438 36258
rect 16650 36255 16662 36258
rect 15426 36209 16662 36255
rect 15426 36206 15438 36209
rect 16650 36206 16662 36209
rect 16714 36206 16726 36258
rect 11790 36194 11842 36206
rect 29374 36194 29426 36206
rect 1344 36090 44576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 44576 36090
rect 1344 36004 44576 36038
rect 30718 35922 30770 35934
rect 30718 35858 30770 35870
rect 20190 35810 20242 35822
rect 29598 35810 29650 35822
rect 16650 35758 16662 35810
rect 16714 35758 16726 35810
rect 26618 35758 26630 35810
rect 26682 35758 26694 35810
rect 20190 35746 20242 35758
rect 29598 35746 29650 35758
rect 34302 35810 34354 35822
rect 34302 35746 34354 35758
rect 34694 35810 34746 35822
rect 34694 35746 34746 35758
rect 37886 35754 37938 35766
rect 37326 35726 37378 35738
rect 9550 35698 9602 35710
rect 12574 35698 12626 35710
rect 10414 35646 10426 35698
rect 10478 35646 10490 35698
rect 11685 35646 11697 35698
rect 11749 35646 11761 35698
rect 9550 35634 9602 35646
rect 12574 35634 12626 35646
rect 13134 35698 13186 35710
rect 13134 35634 13186 35646
rect 15822 35698 15874 35710
rect 15822 35634 15874 35646
rect 16158 35698 16210 35710
rect 16158 35634 16210 35646
rect 16382 35698 16434 35710
rect 16382 35634 16434 35646
rect 17278 35698 17330 35710
rect 17278 35634 17330 35646
rect 22878 35698 22930 35710
rect 22878 35634 22930 35646
rect 26126 35698 26178 35710
rect 26126 35634 26178 35646
rect 26350 35698 26402 35710
rect 26350 35634 26402 35646
rect 26910 35698 26962 35710
rect 31054 35698 31106 35710
rect 27682 35646 27694 35698
rect 27746 35646 27758 35698
rect 26910 35634 26962 35646
rect 31054 35634 31106 35646
rect 31838 35698 31890 35710
rect 33070 35698 33122 35710
rect 32050 35646 32062 35698
rect 32114 35646 32126 35698
rect 32386 35646 32398 35698
rect 32450 35646 32462 35698
rect 31838 35634 31890 35646
rect 33070 35634 33122 35646
rect 33182 35698 33234 35710
rect 33182 35634 33234 35646
rect 33966 35698 34018 35710
rect 34414 35698 34466 35710
rect 33966 35634 34018 35646
rect 34134 35642 34186 35654
rect 23270 35586 23322 35598
rect 13906 35534 13918 35586
rect 13970 35534 13982 35586
rect 22082 35534 22094 35586
rect 22146 35534 22158 35586
rect 23270 35522 23322 35534
rect 25958 35586 26010 35598
rect 25958 35522 26010 35534
rect 31502 35586 31554 35598
rect 34414 35634 34466 35646
rect 34974 35698 35026 35710
rect 34974 35634 35026 35646
rect 35198 35698 35250 35710
rect 35466 35646 35478 35698
rect 35530 35646 35542 35698
rect 37538 35702 37550 35754
rect 37602 35702 37614 35754
rect 37762 35702 37774 35754
rect 37826 35702 37838 35754
rect 37886 35690 37938 35702
rect 39790 35698 39842 35710
rect 37326 35662 37378 35674
rect 35198 35634 35250 35646
rect 39790 35634 39842 35646
rect 39902 35698 39954 35710
rect 39902 35634 39954 35646
rect 40798 35698 40850 35710
rect 40798 35634 40850 35646
rect 31502 35522 31554 35534
rect 32510 35530 32562 35542
rect 33450 35534 33462 35586
rect 33514 35534 33526 35586
rect 34134 35578 34186 35590
rect 39454 35586 39506 35598
rect 41570 35534 41582 35586
rect 41634 35534 41646 35586
rect 43474 35534 43486 35586
rect 43538 35534 43550 35586
rect 10670 35474 10722 35486
rect 10670 35410 10722 35422
rect 11454 35474 11506 35486
rect 11454 35410 11506 35422
rect 17614 35474 17666 35486
rect 39454 35522 39506 35534
rect 32510 35466 32562 35478
rect 37046 35474 37098 35486
rect 17614 35410 17666 35422
rect 37046 35410 37098 35422
rect 40238 35474 40290 35486
rect 40238 35410 40290 35422
rect 1344 35306 44576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 44576 35306
rect 1344 35220 44576 35254
rect 21422 35138 21474 35150
rect 21422 35074 21474 35086
rect 31614 35138 31666 35150
rect 31614 35074 31666 35086
rect 43150 35138 43202 35150
rect 43150 35074 43202 35086
rect 27974 35026 28026 35038
rect 36318 35026 36370 35038
rect 10322 34974 10334 35026
rect 10386 34974 10398 35026
rect 32386 34974 32398 35026
rect 32450 34974 32462 35026
rect 37090 34974 37102 35026
rect 37154 34974 37166 35026
rect 40674 34974 40686 35026
rect 40738 34974 40750 35026
rect 27974 34962 28026 34974
rect 36318 34962 36370 34974
rect 13022 34914 13074 34926
rect 12226 34862 12238 34914
rect 12290 34862 12302 34914
rect 13022 34850 13074 34862
rect 13358 34914 13410 34926
rect 13358 34850 13410 34862
rect 15150 34914 15202 34926
rect 18174 34914 18226 34926
rect 17378 34862 17390 34914
rect 17442 34862 17454 34914
rect 15150 34850 15202 34862
rect 18174 34850 18226 34862
rect 18286 34914 18338 34926
rect 18286 34850 18338 34862
rect 18622 34914 18674 34926
rect 18622 34850 18674 34862
rect 21758 34914 21810 34926
rect 21758 34850 21810 34862
rect 25678 34914 25730 34926
rect 25678 34850 25730 34862
rect 31950 34914 32002 34926
rect 35086 34914 35138 34926
rect 34290 34862 34302 34914
rect 34354 34862 34366 34914
rect 31950 34850 32002 34862
rect 35086 34850 35138 34862
rect 35646 34914 35698 34926
rect 35926 34914 35978 34926
rect 39790 34914 39842 34926
rect 35746 34862 35758 34914
rect 35810 34862 35822 34914
rect 38994 34862 39006 34914
rect 39058 34862 39070 34914
rect 35646 34850 35698 34862
rect 35926 34850 35978 34862
rect 39790 34850 39842 34862
rect 39902 34914 39954 34926
rect 39902 34850 39954 34862
rect 43486 34914 43538 34926
rect 43486 34850 43538 34862
rect 15486 34802 15538 34814
rect 15486 34738 15538 34750
rect 42590 34802 42642 34814
rect 42590 34738 42642 34750
rect 13694 34690 13746 34702
rect 13694 34626 13746 34638
rect 14814 34690 14866 34702
rect 14814 34626 14866 34638
rect 31222 34690 31274 34702
rect 31222 34626 31274 34638
rect 1344 34522 44576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 44576 34522
rect 1344 34436 44576 34470
rect 26910 34354 26962 34366
rect 26910 34290 26962 34302
rect 13694 34242 13746 34254
rect 13694 34178 13746 34190
rect 33070 34242 33122 34254
rect 33070 34178 33122 34190
rect 37326 34186 37378 34198
rect 9102 34130 9154 34142
rect 10782 34130 10834 34142
rect 9893 34078 9905 34130
rect 9957 34078 9969 34130
rect 9102 34066 9154 34078
rect 10782 34066 10834 34078
rect 11006 34130 11058 34142
rect 14030 34130 14082 34142
rect 17278 34130 17330 34142
rect 24558 34130 24610 34142
rect 11778 34078 11790 34130
rect 11842 34078 11854 34130
rect 14802 34078 14814 34130
rect 14866 34078 14878 34130
rect 18050 34078 18062 34130
rect 18114 34078 18126 34130
rect 11006 34066 11058 34078
rect 14030 34066 14082 34078
rect 17278 34066 17330 34078
rect 24558 34066 24610 34078
rect 24782 34130 24834 34142
rect 25442 34078 25454 34130
rect 25506 34078 25518 34130
rect 28242 34105 28254 34157
rect 28306 34105 28318 34157
rect 31938 34078 31950 34130
rect 32002 34078 32014 34130
rect 32274 34078 32286 34130
rect 32338 34078 32350 34130
rect 33196 34118 33208 34170
rect 33260 34118 33272 34170
rect 33506 34111 33518 34163
rect 33570 34111 33582 34163
rect 33842 34114 33854 34166
rect 33906 34114 33918 34166
rect 34178 34134 34190 34186
rect 34242 34134 34254 34186
rect 36766 34158 36818 34170
rect 35310 34130 35362 34142
rect 34738 34078 34750 34130
rect 34802 34078 34814 34130
rect 35074 34078 35086 34130
rect 35138 34078 35150 34130
rect 36978 34134 36990 34186
rect 37042 34134 37054 34186
rect 37214 34158 37266 34170
rect 36766 34094 36818 34106
rect 37326 34122 37378 34134
rect 37214 34094 37266 34106
rect 37874 34105 37886 34157
rect 37938 34105 37950 34157
rect 40798 34130 40850 34142
rect 24782 34066 24834 34078
rect 35310 34066 35362 34078
rect 41570 34078 41582 34130
rect 41634 34078 41646 34130
rect 40798 34066 40850 34078
rect 16706 33966 16718 34018
rect 16770 33966 16782 34018
rect 19954 33966 19966 34018
rect 20018 33966 20030 34018
rect 32398 33962 32450 33974
rect 8766 33906 8818 33918
rect 8766 33842 8818 33854
rect 9662 33906 9714 33918
rect 25286 33906 25338 33918
rect 24266 33854 24278 33906
rect 24330 33854 24342 33906
rect 32398 33898 32450 33910
rect 34638 33962 34690 33974
rect 43474 33966 43486 34018
rect 43538 33966 43550 34018
rect 34638 33898 34690 33910
rect 35646 33906 35698 33918
rect 9662 33842 9714 33854
rect 25286 33842 25338 33854
rect 35646 33842 35698 33854
rect 36486 33906 36538 33918
rect 36486 33842 36538 33854
rect 38894 33906 38946 33918
rect 38894 33842 38946 33854
rect 1344 33738 44576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 44576 33738
rect 1344 33652 44576 33686
rect 12294 33570 12346 33582
rect 12294 33506 12346 33518
rect 15822 33570 15874 33582
rect 27694 33570 27746 33582
rect 16762 33518 16774 33570
rect 16826 33518 16838 33570
rect 17546 33518 17558 33570
rect 17610 33518 17622 33570
rect 42814 33570 42866 33582
rect 15822 33506 15874 33518
rect 27694 33506 27746 33518
rect 28590 33514 28642 33526
rect 42814 33506 42866 33518
rect 8754 33406 8766 33458
rect 8818 33406 8830 33458
rect 9874 33406 9886 33458
rect 9938 33406 9950 33458
rect 11778 33406 11790 33458
rect 11842 33406 11854 33458
rect 24210 33406 24222 33458
rect 24274 33406 24286 33458
rect 26114 33406 26126 33458
rect 26178 33406 26190 33458
rect 28590 33450 28642 33462
rect 31602 33406 31614 33458
rect 31666 33406 31678 33458
rect 6078 33346 6130 33358
rect 9102 33346 9154 33358
rect 16158 33346 16210 33358
rect 6850 33294 6862 33346
rect 6914 33294 6926 33346
rect 12450 33294 12462 33346
rect 12514 33294 12526 33346
rect 6078 33282 6130 33294
rect 9102 33282 9154 33294
rect 16158 33282 16210 33294
rect 16382 33346 16434 33358
rect 16382 33282 16434 33294
rect 16494 33346 16546 33358
rect 16494 33282 16546 33294
rect 17054 33346 17106 33358
rect 17054 33282 17106 33294
rect 17278 33346 17330 33358
rect 20862 33346 20914 33358
rect 23438 33346 23490 33358
rect 20066 33294 20078 33346
rect 20130 33294 20142 33346
rect 22978 33294 22990 33346
rect 23042 33294 23054 33346
rect 17278 33282 17330 33294
rect 20862 33282 20914 33294
rect 23438 33282 23490 33294
rect 26574 33346 26626 33358
rect 30046 33346 30098 33358
rect 34862 33346 34914 33358
rect 27438 33294 27450 33346
rect 27502 33294 27514 33346
rect 28130 33294 28142 33346
rect 28194 33294 28206 33346
rect 28466 33294 28478 33346
rect 28530 33294 28542 33346
rect 26574 33282 26626 33294
rect 29094 33290 29146 33302
rect 18174 33234 18226 33246
rect 29250 33238 29262 33290
rect 29314 33238 29326 33290
rect 29474 33255 29486 33307
rect 29538 33255 29550 33307
rect 31266 33294 31278 33346
rect 31330 33294 31342 33346
rect 30046 33282 30098 33294
rect 31490 33279 31502 33331
rect 31554 33279 31566 33331
rect 32162 33294 32174 33346
rect 32226 33294 32238 33346
rect 34402 33266 34414 33318
rect 34466 33266 34478 33318
rect 34862 33282 34914 33294
rect 35534 33346 35586 33358
rect 39454 33346 39506 33358
rect 42478 33346 42530 33358
rect 35534 33282 35586 33294
rect 37326 33318 37378 33330
rect 37326 33254 37378 33266
rect 37550 33318 37602 33330
rect 37550 33254 37602 33266
rect 37718 33311 37770 33323
rect 37718 33247 37770 33259
rect 37886 33290 37938 33302
rect 38098 33294 38110 33346
rect 38162 33294 38174 33346
rect 40226 33294 40238 33346
rect 40290 33294 40302 33346
rect 29094 33226 29146 33238
rect 37046 33234 37098 33246
rect 18174 33170 18226 33182
rect 23158 33178 23210 33190
rect 39454 33282 39506 33294
rect 42478 33282 42530 33294
rect 43710 33346 43762 33358
rect 43710 33282 43762 33294
rect 37886 33226 37938 33238
rect 42142 33234 42194 33246
rect 37046 33170 37098 33182
rect 42142 33170 42194 33182
rect 23158 33114 23210 33126
rect 35198 33122 35250 33134
rect 35198 33058 35250 33070
rect 35870 33122 35922 33134
rect 35870 33058 35922 33070
rect 36486 33122 36538 33134
rect 36486 33058 36538 33070
rect 43374 33122 43426 33134
rect 43374 33058 43426 33070
rect 1344 32954 44576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 44576 32954
rect 1344 32868 44576 32902
rect 20078 32786 20130 32798
rect 38334 32786 38386 32798
rect 20078 32722 20130 32734
rect 25398 32730 25450 32742
rect 6414 32674 6466 32686
rect 6414 32610 6466 32622
rect 12238 32674 12290 32686
rect 38334 32722 38386 32734
rect 38838 32786 38890 32798
rect 38838 32722 38890 32734
rect 19114 32622 19126 32674
rect 19178 32622 19190 32674
rect 25398 32666 25450 32678
rect 34022 32674 34074 32686
rect 37662 32674 37714 32686
rect 12238 32610 12290 32622
rect 30904 32599 30956 32611
rect 9102 32562 9154 32574
rect 9102 32498 9154 32510
rect 9550 32562 9602 32574
rect 17726 32562 17778 32574
rect 10322 32510 10334 32562
rect 10386 32510 10398 32562
rect 9550 32498 9602 32510
rect 17726 32498 17778 32510
rect 17950 32562 18002 32574
rect 17950 32498 18002 32510
rect 19406 32562 19458 32574
rect 19406 32498 19458 32510
rect 19630 32562 19682 32574
rect 19630 32498 19682 32510
rect 19742 32562 19794 32574
rect 19742 32498 19794 32510
rect 20862 32562 20914 32574
rect 25678 32562 25730 32574
rect 21634 32510 21646 32562
rect 21698 32510 21710 32562
rect 24322 32510 24334 32562
rect 24386 32510 24398 32562
rect 24546 32510 24558 32562
rect 24610 32510 24622 32562
rect 25218 32510 25230 32562
rect 25282 32510 25294 32562
rect 20862 32498 20914 32510
rect 25678 32498 25730 32510
rect 28366 32562 28418 32574
rect 30606 32562 30658 32574
rect 29026 32510 29038 32562
rect 29090 32510 29102 32562
rect 30706 32510 30718 32562
rect 30770 32510 30782 32562
rect 31984 32599 32036 32611
rect 34022 32610 34074 32622
rect 34750 32618 34802 32630
rect 30904 32535 30956 32547
rect 31726 32562 31778 32574
rect 31826 32510 31838 32562
rect 31890 32510 31902 32562
rect 34302 32562 34354 32574
rect 34570 32566 34582 32618
rect 34634 32566 34646 32618
rect 37662 32610 37714 32622
rect 39510 32674 39562 32686
rect 39510 32610 39562 32622
rect 40350 32618 40402 32630
rect 31984 32535 32036 32547
rect 33394 32510 33406 32562
rect 33458 32510 33470 32562
rect 34402 32510 34414 32562
rect 34466 32510 34478 32562
rect 34750 32554 34802 32566
rect 34974 32562 35026 32574
rect 37998 32562 38050 32574
rect 39778 32566 39790 32618
rect 39842 32566 39854 32618
rect 40014 32590 40066 32602
rect 35746 32510 35758 32562
rect 35810 32510 35822 32562
rect 38658 32510 38670 32562
rect 38722 32510 38734 32562
rect 40014 32526 40066 32538
rect 40182 32597 40234 32609
rect 40350 32554 40402 32566
rect 40182 32533 40234 32545
rect 43810 32537 43822 32589
rect 43874 32537 43886 32589
rect 28366 32498 28418 32510
rect 30606 32498 30658 32510
rect 31726 32498 31778 32510
rect 34302 32498 34354 32510
rect 34974 32498 35026 32510
rect 37998 32498 38050 32510
rect 8306 32398 8318 32450
rect 8370 32398 8382 32450
rect 23538 32398 23550 32450
rect 23602 32398 23614 32450
rect 24670 32394 24722 32406
rect 26450 32398 26462 32450
rect 26514 32398 26526 32450
rect 17434 32286 17446 32338
rect 17498 32286 17510 32338
rect 24670 32330 24722 32342
rect 28870 32394 28922 32406
rect 43138 32398 43150 32450
rect 43202 32398 43214 32450
rect 28870 32330 28922 32342
rect 31278 32338 31330 32350
rect 31278 32274 31330 32286
rect 32398 32338 32450 32350
rect 32398 32274 32450 32286
rect 33574 32338 33626 32350
rect 33574 32274 33626 32286
rect 1344 32170 44576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 44576 32170
rect 1344 32084 44576 32118
rect 34078 32002 34130 32014
rect 29654 31946 29706 31958
rect 18062 31890 18114 31902
rect 18062 31826 18114 31838
rect 18846 31890 18898 31902
rect 24726 31890 24778 31902
rect 34078 31938 34130 31950
rect 34582 32002 34634 32014
rect 34582 31938 34634 31950
rect 23874 31838 23886 31890
rect 23938 31838 23950 31890
rect 27906 31838 27918 31890
rect 27970 31838 27982 31890
rect 29654 31882 29706 31894
rect 33182 31890 33234 31902
rect 18846 31826 18898 31838
rect 24726 31826 24778 31838
rect 33182 31826 33234 31838
rect 35142 31834 35194 31846
rect 42242 31838 42254 31890
rect 42306 31838 42318 31890
rect 15038 31778 15090 31790
rect 15038 31714 15090 31726
rect 15598 31778 15650 31790
rect 15598 31714 15650 31726
rect 15710 31778 15762 31790
rect 15710 31714 15762 31726
rect 16830 31778 16882 31790
rect 16830 31714 16882 31726
rect 17726 31778 17778 31790
rect 17726 31714 17778 31726
rect 18398 31778 18450 31790
rect 18398 31714 18450 31726
rect 18510 31778 18562 31790
rect 18510 31714 18562 31726
rect 21198 31778 21250 31790
rect 28702 31778 28754 31790
rect 30270 31778 30322 31790
rect 21970 31726 21982 31778
rect 22034 31726 22046 31778
rect 25454 31750 25506 31762
rect 21198 31714 21250 31726
rect 24994 31670 25006 31722
rect 25058 31670 25070 31722
rect 25218 31670 25230 31722
rect 25282 31670 25294 31722
rect 25610 31710 25622 31762
rect 25674 31710 25686 31762
rect 29026 31726 29038 31778
rect 29090 31726 29102 31778
rect 29474 31726 29486 31778
rect 29538 31726 29550 31778
rect 28702 31714 28754 31726
rect 30270 31714 30322 31726
rect 31390 31778 31442 31790
rect 33406 31778 33458 31790
rect 34862 31778 34914 31790
rect 31826 31726 31838 31778
rect 31890 31726 31902 31778
rect 32162 31726 32174 31778
rect 32226 31726 32238 31778
rect 32722 31726 32734 31778
rect 32786 31726 32798 31778
rect 32946 31726 32958 31778
rect 33010 31726 33022 31778
rect 33506 31726 33518 31778
rect 33570 31726 33582 31778
rect 34962 31726 34974 31778
rect 35026 31726 35038 31778
rect 35142 31770 35194 31782
rect 35310 31778 35362 31790
rect 25454 31686 25506 31698
rect 26014 31666 26066 31678
rect 31134 31670 31146 31722
rect 31198 31670 31210 31722
rect 31390 31714 31442 31726
rect 33406 31714 33458 31726
rect 33674 31670 33686 31722
rect 33738 31670 33750 31722
rect 34862 31714 34914 31726
rect 35310 31714 35362 31726
rect 35534 31778 35586 31790
rect 35534 31714 35586 31726
rect 35758 31778 35810 31790
rect 35758 31714 35810 31726
rect 39566 31778 39618 31790
rect 40338 31726 40350 31778
rect 40402 31726 40414 31778
rect 39566 31714 39618 31726
rect 15306 31614 15318 31666
rect 15370 31614 15382 31666
rect 36026 31614 36038 31666
rect 36090 31614 36102 31666
rect 26014 31602 26066 31614
rect 14702 31554 14754 31566
rect 14702 31490 14754 31502
rect 16494 31554 16546 31566
rect 16494 31490 16546 31502
rect 17390 31554 17442 31566
rect 17390 31490 17442 31502
rect 29206 31554 29258 31566
rect 29206 31490 29258 31502
rect 42870 31554 42922 31566
rect 42870 31490 42922 31502
rect 1344 31386 44576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 44576 31386
rect 1344 31300 44576 31334
rect 18398 31218 18450 31230
rect 18398 31154 18450 31166
rect 30326 31218 30378 31230
rect 30326 31154 30378 31166
rect 15374 31106 15426 31118
rect 29598 31106 29650 31118
rect 17434 31054 17446 31106
rect 17498 31054 17510 31106
rect 28970 31054 28982 31106
rect 29034 31054 29046 31106
rect 37662 31106 37714 31118
rect 15374 31042 15426 31054
rect 27246 31033 27298 31045
rect 29598 31042 29650 31054
rect 31614 31050 31666 31062
rect 20078 31014 20130 31026
rect 12686 30994 12738 31006
rect 16270 30994 16322 31006
rect 13458 30942 13470 30994
rect 13522 30942 13534 30994
rect 12686 30930 12738 30942
rect 16270 30930 16322 30942
rect 16494 30994 16546 31006
rect 16494 30930 16546 30942
rect 17726 30994 17778 31006
rect 17726 30930 17778 30942
rect 17838 30994 17890 31006
rect 17838 30930 17890 30942
rect 18062 30994 18114 31006
rect 20078 30950 20130 30962
rect 20190 30994 20242 31006
rect 22878 30994 22930 31006
rect 18062 30930 18114 30942
rect 20962 30942 20974 30994
rect 21026 30942 21038 30994
rect 20190 30930 20242 30942
rect 22878 30930 22930 30942
rect 25454 30994 25506 31006
rect 25454 30930 25506 30942
rect 25790 30994 25842 31006
rect 26114 30969 26126 31021
rect 26178 30969 26190 31021
rect 26450 30942 26462 30994
rect 26514 30942 26526 30994
rect 26786 30942 26798 30994
rect 26850 30942 26862 30994
rect 27246 30969 27298 30981
rect 27470 30994 27522 31006
rect 25790 30930 25842 30942
rect 27470 30930 27522 30942
rect 27806 30994 27858 31006
rect 27806 30930 27858 30942
rect 28478 30994 28530 31006
rect 28478 30930 28530 30942
rect 28702 30994 28754 31006
rect 28702 30930 28754 30942
rect 29262 30994 29314 31006
rect 30606 30994 30658 31006
rect 30146 30942 30158 30994
rect 30210 30942 30222 30994
rect 29262 30930 29314 30942
rect 30606 30930 30658 30942
rect 30830 30994 30882 31006
rect 31714 30998 31726 31050
rect 31778 30998 31790 31050
rect 31938 30998 31950 31050
rect 32002 30998 32014 31050
rect 37662 31042 37714 31054
rect 32174 31022 32226 31034
rect 31098 30942 31110 30994
rect 31162 30942 31174 30994
rect 31614 30986 31666 30998
rect 32174 30958 32226 30970
rect 33070 30994 33122 31006
rect 33350 30994 33402 31006
rect 34974 30994 35026 31006
rect 42366 30994 42418 31006
rect 33170 30942 33182 30994
rect 33234 30942 33246 30994
rect 34178 30942 34190 30994
rect 34242 30942 34254 30994
rect 34514 30942 34526 30994
rect 34578 30942 34590 30994
rect 35746 30942 35758 30994
rect 35810 30942 35822 30994
rect 41458 30942 41470 30994
rect 41522 30942 41534 30994
rect 30830 30930 30882 30942
rect 33070 30930 33122 30942
rect 33350 30930 33402 30942
rect 34974 30930 35026 30942
rect 42366 30930 42418 30942
rect 27134 30882 27186 30894
rect 26226 30830 26238 30882
rect 26290 30830 26302 30882
rect 27134 30818 27186 30830
rect 19910 30770 19962 30782
rect 16762 30718 16774 30770
rect 16826 30718 16838 30770
rect 19910 30706 19962 30718
rect 32454 30770 32506 30782
rect 32454 30706 32506 30718
rect 33742 30770 33794 30782
rect 34402 30774 34414 30826
rect 34466 30774 34478 30826
rect 33742 30706 33794 30718
rect 41302 30770 41354 30782
rect 41302 30706 41354 30718
rect 42702 30770 42754 30782
rect 42702 30706 42754 30718
rect 1344 30602 44576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 44576 30602
rect 1344 30516 44576 30550
rect 20638 30434 20690 30446
rect 20638 30370 20690 30382
rect 28086 30434 28138 30446
rect 28086 30370 28138 30382
rect 32734 30434 32786 30446
rect 32734 30370 32786 30382
rect 33854 30434 33906 30446
rect 33854 30370 33906 30382
rect 17826 30270 17838 30322
rect 17890 30270 17902 30322
rect 19730 30270 19742 30322
rect 19794 30270 19806 30322
rect 21970 30270 21982 30322
rect 22034 30270 22046 30322
rect 40450 30270 40462 30322
rect 40514 30270 40526 30322
rect 13918 30210 13970 30222
rect 13918 30146 13970 30158
rect 14030 30210 14082 30222
rect 16718 30210 16770 30222
rect 14802 30158 14814 30210
rect 14866 30158 14878 30210
rect 14030 30146 14082 30158
rect 16718 30146 16770 30158
rect 17054 30210 17106 30222
rect 17054 30146 17106 30158
rect 20302 30210 20354 30222
rect 20302 30146 20354 30158
rect 21198 30210 21250 30222
rect 21198 30146 21250 30158
rect 23886 30210 23938 30222
rect 23886 30146 23938 30158
rect 24222 30210 24274 30222
rect 24222 30146 24274 30158
rect 25006 30210 25058 30222
rect 25006 30146 25058 30158
rect 25230 30210 25282 30222
rect 26350 30210 26402 30222
rect 25498 30158 25510 30210
rect 25562 30158 25574 30210
rect 31614 30210 31666 30222
rect 25230 30146 25282 30158
rect 26350 30146 26402 30158
rect 27246 30175 27298 30187
rect 27246 30111 27298 30123
rect 27414 30175 27466 30187
rect 27414 30111 27466 30123
rect 27638 30175 27690 30187
rect 27638 30111 27690 30123
rect 27862 30175 27914 30187
rect 31614 30146 31666 30158
rect 33182 30210 33234 30222
rect 33462 30210 33514 30222
rect 33282 30158 33294 30210
rect 33346 30158 33358 30210
rect 27862 30111 27914 30123
rect 32478 30102 32490 30154
rect 32542 30102 32554 30154
rect 33182 30146 33234 30158
rect 33462 30146 33514 30158
rect 37774 30210 37826 30222
rect 37774 30146 37826 30158
rect 38110 30210 38162 30222
rect 38110 30146 38162 30158
rect 38558 30210 38610 30222
rect 38558 30146 38610 30158
rect 39678 30210 39730 30222
rect 39678 30146 39730 30158
rect 42366 30210 42418 30222
rect 42366 30146 42418 30158
rect 13582 29986 13634 29998
rect 13582 29922 13634 29934
rect 24558 29986 24610 29998
rect 24558 29922 24610 29934
rect 26686 29986 26738 29998
rect 26686 29922 26738 29934
rect 37606 29986 37658 29998
rect 37606 29922 37658 29934
rect 38894 29986 38946 29998
rect 38894 29922 38946 29934
rect 39510 29986 39562 29998
rect 39510 29922 39562 29934
rect 42982 29986 43034 29998
rect 42982 29922 43034 29934
rect 1344 29818 44576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 44576 29818
rect 1344 29732 44576 29766
rect 18622 29650 18674 29662
rect 18622 29586 18674 29598
rect 25902 29650 25954 29662
rect 43374 29650 43426 29662
rect 26674 29598 26686 29650
rect 26738 29647 26750 29650
rect 27234 29647 27246 29650
rect 26738 29601 27246 29647
rect 26738 29598 26750 29601
rect 27234 29598 27246 29601
rect 27298 29598 27310 29650
rect 25902 29586 25954 29598
rect 43374 29586 43426 29598
rect 16158 29538 16210 29550
rect 19742 29538 19794 29550
rect 18106 29486 18118 29538
rect 18170 29486 18182 29538
rect 16158 29474 16210 29486
rect 19742 29474 19794 29486
rect 32398 29538 32450 29550
rect 32398 29474 32450 29486
rect 13470 29426 13522 29438
rect 17726 29426 17778 29438
rect 14242 29374 14254 29426
rect 14306 29374 14318 29426
rect 13470 29362 13522 29374
rect 17726 29362 17778 29374
rect 17838 29426 17890 29438
rect 17838 29362 17890 29374
rect 18958 29426 19010 29438
rect 22430 29426 22482 29438
rect 21634 29374 21646 29426
rect 21698 29374 21710 29426
rect 18958 29362 19010 29374
rect 22430 29362 22482 29374
rect 22822 29426 22874 29438
rect 22822 29362 22874 29374
rect 23550 29426 23602 29438
rect 23550 29362 23602 29374
rect 24222 29426 24274 29438
rect 24222 29362 24274 29374
rect 25566 29426 25618 29438
rect 25566 29362 25618 29374
rect 31278 29426 31330 29438
rect 32142 29374 32154 29426
rect 32206 29374 32218 29426
rect 36306 29374 36318 29426
rect 36370 29374 36382 29426
rect 36866 29374 36878 29426
rect 36930 29374 36942 29426
rect 37202 29374 37214 29426
rect 37266 29374 37278 29426
rect 37426 29389 37438 29441
rect 37490 29389 37502 29441
rect 40002 29401 40014 29453
rect 40066 29401 40078 29453
rect 40898 29374 40910 29426
rect 40962 29374 40974 29426
rect 41234 29389 41246 29441
rect 41298 29389 41310 29441
rect 41906 29401 41918 29453
rect 41970 29401 41982 29453
rect 31278 29362 31330 29374
rect 37538 29262 37550 29314
rect 37602 29262 37614 29314
rect 39330 29262 39342 29314
rect 39394 29262 39406 29314
rect 41346 29262 41358 29314
rect 41410 29262 41422 29314
rect 23214 29202 23266 29214
rect 23214 29138 23266 29150
rect 23886 29202 23938 29214
rect 23886 29138 23938 29150
rect 36150 29202 36202 29214
rect 36150 29138 36202 29150
rect 36710 29202 36762 29214
rect 36710 29138 36762 29150
rect 1344 29034 44576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 44576 29034
rect 1344 28948 44576 28982
rect 25902 28866 25954 28878
rect 31882 28814 31894 28866
rect 31946 28814 31958 28866
rect 25902 28802 25954 28814
rect 31042 28758 31054 28810
rect 31106 28758 31118 28810
rect 15922 28702 15934 28754
rect 15986 28702 15998 28754
rect 17826 28702 17838 28754
rect 17890 28702 17902 28754
rect 35858 28702 35870 28754
rect 35922 28702 35934 28754
rect 36978 28702 36990 28754
rect 37042 28702 37054 28754
rect 38658 28702 38670 28754
rect 38722 28702 38734 28754
rect 43586 28702 43598 28754
rect 43650 28702 43662 28754
rect 15150 28642 15202 28654
rect 15150 28578 15202 28590
rect 20862 28642 20914 28654
rect 20862 28578 20914 28590
rect 21310 28642 21362 28654
rect 24110 28642 24162 28654
rect 22174 28590 22186 28642
rect 22238 28590 22250 28642
rect 21310 28578 21362 28590
rect 24110 28578 24162 28590
rect 24222 28642 24274 28654
rect 24222 28578 24274 28590
rect 24558 28642 24610 28654
rect 24558 28578 24610 28590
rect 25566 28642 25618 28654
rect 25566 28578 25618 28590
rect 26238 28642 26290 28654
rect 31390 28642 31442 28654
rect 26450 28590 26462 28642
rect 26514 28590 26526 28642
rect 26238 28578 26290 28590
rect 26786 28575 26798 28627
rect 26850 28575 26862 28627
rect 27234 28590 27246 28642
rect 27298 28590 27310 28642
rect 27570 28575 27582 28627
rect 27634 28575 27646 28627
rect 30818 28590 30830 28642
rect 30882 28590 30894 28642
rect 31042 28590 31054 28642
rect 31106 28590 31118 28642
rect 31390 28578 31442 28590
rect 31614 28642 31666 28654
rect 37886 28642 37938 28654
rect 31614 28578 31666 28590
rect 34738 28562 34750 28614
rect 34802 28562 34814 28614
rect 35410 28590 35422 28642
rect 35474 28590 35486 28642
rect 35746 28546 35758 28598
rect 35810 28546 35822 28598
rect 36418 28590 36430 28642
rect 36482 28590 36494 28642
rect 37090 28546 37102 28598
rect 37154 28546 37166 28598
rect 37314 28590 37326 28642
rect 37378 28590 37390 28642
rect 37886 28578 37938 28590
rect 40910 28642 40962 28654
rect 41682 28590 41694 28642
rect 41746 28590 41758 28642
rect 40910 28578 40962 28590
rect 22430 28530 22482 28542
rect 22430 28466 22482 28478
rect 40574 28530 40626 28542
rect 20526 28418 20578 28430
rect 20526 28354 20578 28366
rect 23774 28418 23826 28430
rect 23774 28354 23826 28366
rect 25230 28418 25282 28430
rect 26562 28422 26574 28474
rect 26626 28422 26638 28474
rect 27346 28422 27358 28474
rect 27410 28422 27422 28474
rect 40574 28466 40626 28478
rect 25230 28354 25282 28366
rect 33742 28418 33794 28430
rect 33742 28354 33794 28366
rect 36262 28418 36314 28430
rect 36262 28354 36314 28366
rect 44214 28418 44266 28430
rect 44214 28354 44266 28366
rect 1344 28250 44576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 44576 28250
rect 1344 28164 44576 28198
rect 16494 28082 16546 28094
rect 16494 28018 16546 28030
rect 31166 28082 31218 28094
rect 31166 28018 31218 28030
rect 24110 27970 24162 27982
rect 24110 27906 24162 27918
rect 28254 27970 28306 27982
rect 33954 27974 33966 28026
rect 34018 27974 34030 28026
rect 28254 27906 28306 27918
rect 34526 27970 34578 27982
rect 34526 27906 34578 27918
rect 16830 27858 16882 27870
rect 11778 27806 11790 27858
rect 11842 27806 11854 27858
rect 16830 27794 16882 27806
rect 21422 27858 21474 27870
rect 24726 27858 24778 27870
rect 22194 27806 22206 27858
rect 22258 27806 22270 27858
rect 21422 27794 21474 27806
rect 24726 27794 24778 27806
rect 25566 27858 25618 27870
rect 26338 27806 26350 27858
rect 26402 27806 26414 27858
rect 28802 27850 28814 27902
rect 28866 27850 28878 27902
rect 29138 27806 29150 27858
rect 29202 27806 29214 27858
rect 29810 27806 29822 27858
rect 29874 27806 29886 27858
rect 32498 27833 32510 27885
rect 32562 27833 32574 27885
rect 33730 27850 33742 27902
rect 33794 27850 33806 27902
rect 37214 27858 37266 27870
rect 40462 27858 40514 27870
rect 34066 27806 34078 27858
rect 34130 27806 34142 27858
rect 36418 27806 36430 27858
rect 36482 27806 36494 27858
rect 39666 27806 39678 27858
rect 39730 27806 39742 27858
rect 25566 27794 25618 27806
rect 37214 27794 37266 27806
rect 40462 27794 40514 27806
rect 41134 27858 41186 27870
rect 41134 27794 41186 27806
rect 28690 27694 28702 27746
rect 28754 27694 28766 27746
rect 37762 27694 37774 27746
rect 37826 27694 37838 27746
rect 41906 27694 41918 27746
rect 41970 27694 41982 27746
rect 43810 27694 43822 27746
rect 43874 27694 43886 27746
rect 11622 27634 11674 27646
rect 11622 27570 11674 27582
rect 29654 27634 29706 27646
rect 29654 27570 29706 27582
rect 1344 27466 44576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 44576 27466
rect 1344 27380 44576 27414
rect 14142 27298 14194 27310
rect 14142 27234 14194 27246
rect 20526 27298 20578 27310
rect 20526 27234 20578 27246
rect 21422 27298 21474 27310
rect 37998 27298 38050 27310
rect 22586 27246 22598 27298
rect 22650 27246 22662 27298
rect 21422 27234 21474 27246
rect 27794 27190 27806 27242
rect 27858 27190 27870 27242
rect 37998 27234 38050 27246
rect 40854 27298 40906 27310
rect 40854 27234 40906 27246
rect 12786 27134 12798 27186
rect 12850 27134 12862 27186
rect 15586 27134 15598 27186
rect 15650 27134 15662 27186
rect 23650 27134 23662 27186
rect 23714 27134 23726 27186
rect 25554 27134 25566 27186
rect 25618 27134 25630 27186
rect 30258 27134 30270 27186
rect 30322 27134 30334 27186
rect 32162 27134 32174 27186
rect 32226 27134 32238 27186
rect 33394 27134 33406 27186
rect 33458 27134 33470 27186
rect 34402 27134 34414 27186
rect 34466 27134 34478 27186
rect 36306 27134 36318 27186
rect 36370 27134 36382 27186
rect 10110 27074 10162 27086
rect 14478 27074 14530 27086
rect 19462 27074 19514 27086
rect 10882 27022 10894 27074
rect 10946 27022 10958 27074
rect 16034 27022 16046 27074
rect 16098 27022 16110 27074
rect 16594 27022 16606 27074
rect 16658 27022 16670 27074
rect 10110 27010 10162 27022
rect 14478 27010 14530 27022
rect 15754 26966 15766 27018
rect 15818 26966 15830 27018
rect 19462 27010 19514 27022
rect 19854 27074 19906 27086
rect 19854 27010 19906 27022
rect 20190 27074 20242 27086
rect 20190 27010 20242 27022
rect 20862 27074 20914 27086
rect 20862 27010 20914 27022
rect 21758 27074 21810 27086
rect 21758 27010 21810 27022
rect 22878 27074 22930 27086
rect 22878 27010 22930 27022
rect 23102 27074 23154 27086
rect 23102 27010 23154 27022
rect 26350 27074 26402 27086
rect 27246 27074 27298 27086
rect 28590 27074 28642 27086
rect 26562 27022 26574 27074
rect 26626 27022 26638 27074
rect 28018 27022 28030 27074
rect 28082 27022 28094 27074
rect 26350 27010 26402 27022
rect 22150 26962 22202 26974
rect 26898 26966 26910 27018
rect 26962 26966 26974 27018
rect 27246 27010 27298 27022
rect 28590 27010 28642 27022
rect 29486 27074 29538 27086
rect 33630 27074 33682 27086
rect 32946 27022 32958 27074
rect 33010 27022 33022 27074
rect 29486 27010 29538 27022
rect 33282 27007 33294 27059
rect 33346 27007 33358 27059
rect 39678 27074 39730 27086
rect 41134 27074 41186 27086
rect 33630 27010 33682 27022
rect 36978 26994 36990 27046
rect 37042 26994 37054 27046
rect 40674 27022 40686 27074
rect 40738 27022 40750 27074
rect 41906 27022 41918 27074
rect 41970 27022 41982 27074
rect 39678 27010 39730 27022
rect 41134 27010 41186 27022
rect 16774 26906 16826 26918
rect 22150 26898 22202 26910
rect 43822 26962 43874 26974
rect 16774 26842 16826 26854
rect 18566 26850 18618 26862
rect 26674 26854 26686 26906
rect 26738 26854 26750 26906
rect 43822 26898 43874 26910
rect 18566 26786 18618 26798
rect 1344 26682 44576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 44576 26682
rect 1344 26596 44576 26630
rect 9718 26514 9770 26526
rect 9718 26450 9770 26462
rect 22318 26514 22370 26526
rect 33238 26514 33290 26526
rect 22318 26450 22370 26462
rect 26238 26458 26290 26470
rect 16494 26402 16546 26414
rect 33238 26450 33290 26462
rect 40182 26514 40234 26526
rect 40182 26450 40234 26462
rect 42254 26514 42306 26526
rect 42254 26450 42306 26462
rect 26238 26394 26290 26406
rect 29710 26402 29762 26414
rect 16494 26338 16546 26350
rect 9874 26238 9886 26290
rect 9938 26238 9950 26290
rect 10210 26238 10222 26290
rect 10274 26238 10286 26290
rect 10434 26282 10446 26334
rect 10498 26282 10510 26334
rect 18118 26319 18170 26331
rect 10782 26290 10834 26302
rect 10782 26226 10834 26238
rect 13806 26290 13858 26302
rect 14578 26238 14590 26290
rect 14642 26238 14654 26290
rect 17266 26238 17278 26290
rect 17330 26238 17342 26290
rect 17826 26238 17838 26290
rect 17890 26238 17902 26290
rect 18118 26255 18170 26267
rect 18734 26290 18786 26302
rect 13806 26226 13858 26238
rect 18734 26226 18786 26238
rect 19070 26290 19122 26302
rect 19070 26226 19122 26238
rect 19742 26290 19794 26302
rect 20066 26238 20078 26290
rect 20130 26238 20142 26290
rect 20402 26282 20414 26334
rect 20466 26282 20478 26334
rect 26350 26329 26402 26341
rect 29710 26338 29762 26350
rect 37774 26402 37826 26414
rect 37774 26338 37826 26350
rect 20782 26276 20794 26328
rect 20846 26276 20858 26328
rect 22654 26290 22706 26302
rect 25118 26290 25170 26302
rect 21522 26238 21534 26290
rect 21586 26238 21598 26290
rect 23090 26238 23102 26290
rect 23154 26238 23166 26290
rect 19742 26226 19794 26238
rect 22654 26226 22706 26238
rect 25118 26226 25170 26238
rect 25454 26290 25506 26302
rect 26002 26238 26014 26290
rect 26066 26238 26078 26290
rect 26350 26265 26402 26277
rect 26574 26290 26626 26302
rect 25454 26226 25506 26238
rect 26574 26226 26626 26238
rect 27022 26290 27074 26302
rect 27022 26226 27074 26238
rect 30942 26290 30994 26302
rect 32162 26282 32174 26334
rect 32226 26282 32238 26334
rect 33630 26290 33682 26302
rect 35086 26290 35138 26302
rect 38558 26290 38610 26302
rect 32498 26238 32510 26290
rect 32562 26238 32574 26290
rect 33058 26238 33070 26290
rect 33122 26238 33134 26290
rect 34494 26238 34506 26290
rect 34558 26238 34570 26290
rect 35858 26238 35870 26290
rect 35922 26238 35934 26290
rect 39422 26238 39434 26290
rect 39486 26238 39498 26290
rect 40338 26238 40350 26290
rect 40402 26238 40414 26290
rect 41234 26265 41246 26317
rect 41298 26265 41310 26317
rect 43866 26294 43878 26346
rect 43930 26294 43942 26346
rect 44034 26294 44046 26346
rect 44098 26294 44110 26346
rect 30942 26226 30994 26238
rect 33630 26226 33682 26238
rect 35086 26226 35138 26238
rect 38558 26226 38610 26238
rect 10546 26126 10558 26178
rect 10610 26126 10622 26178
rect 11554 26126 11566 26178
rect 11618 26126 11630 26178
rect 13458 26126 13470 26178
rect 13522 26126 13534 26178
rect 18274 26126 18286 26178
rect 18338 26126 18350 26178
rect 20514 26126 20526 26178
rect 20578 26126 20590 26178
rect 21646 26122 21698 26134
rect 27794 26126 27806 26178
rect 27858 26126 27870 26178
rect 32050 26126 32062 26178
rect 32114 26126 32126 26178
rect 43698 26126 43710 26178
rect 43762 26126 43774 26178
rect 17446 26066 17498 26078
rect 17446 26002 17498 26014
rect 19406 26066 19458 26078
rect 21646 26058 21698 26070
rect 22934 26066 22986 26078
rect 19406 26002 19458 26014
rect 22934 26002 22986 26014
rect 30606 26066 30658 26078
rect 30606 26002 30658 26014
rect 34750 26066 34802 26078
rect 34750 26002 34802 26014
rect 39678 26066 39730 26078
rect 39678 26002 39730 26014
rect 1344 25898 44576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 44576 25898
rect 1344 25812 44576 25846
rect 28142 25730 28194 25742
rect 14086 25674 14138 25686
rect 28142 25666 28194 25678
rect 36206 25730 36258 25742
rect 36206 25666 36258 25678
rect 14086 25610 14138 25622
rect 17042 25566 17054 25618
rect 17106 25566 17118 25618
rect 18162 25566 18174 25618
rect 18226 25566 18238 25618
rect 21970 25566 21982 25618
rect 22034 25566 22046 25618
rect 23874 25566 23886 25618
rect 23938 25566 23950 25618
rect 30706 25566 30718 25618
rect 30770 25566 30782 25618
rect 32610 25566 32622 25618
rect 32674 25566 32686 25618
rect 37986 25566 37998 25618
rect 38050 25566 38062 25618
rect 40786 25566 40798 25618
rect 40850 25566 40862 25618
rect 13022 25506 13074 25518
rect 14366 25506 14418 25518
rect 21198 25506 21250 25518
rect 26126 25506 26178 25518
rect 27358 25506 27410 25518
rect 12226 25454 12238 25506
rect 12290 25454 12302 25506
rect 13794 25454 13806 25506
rect 13858 25454 13870 25506
rect 13022 25442 13074 25454
rect 14254 25450 14306 25462
rect 10334 25394 10386 25406
rect 15138 25454 15150 25506
rect 15202 25454 15214 25506
rect 17434 25454 17446 25506
rect 17498 25454 17510 25506
rect 20850 25454 20862 25506
rect 20914 25454 20926 25506
rect 25554 25454 25566 25506
rect 25618 25454 25630 25506
rect 26674 25454 26686 25506
rect 26738 25454 26750 25506
rect 14366 25442 14418 25454
rect 21198 25442 21250 25454
rect 14254 25386 14306 25398
rect 20078 25394 20130 25406
rect 25890 25398 25902 25450
rect 25954 25398 25966 25450
rect 26126 25442 26178 25454
rect 27010 25398 27022 25450
rect 27074 25398 27086 25450
rect 27358 25442 27410 25454
rect 27806 25506 27858 25518
rect 27806 25442 27858 25454
rect 29934 25506 29986 25518
rect 36542 25506 36594 25518
rect 29934 25442 29986 25454
rect 33282 25426 33294 25478
rect 33346 25426 33358 25478
rect 43822 25506 43874 25518
rect 36542 25442 36594 25454
rect 36978 25426 36990 25478
rect 37042 25426 37054 25478
rect 39778 25426 39790 25478
rect 39842 25426 39854 25478
rect 10334 25330 10386 25342
rect 20078 25330 20130 25342
rect 29766 25394 29818 25406
rect 42702 25394 42754 25406
rect 42933 25398 42945 25450
rect 42997 25398 43009 25450
rect 43822 25442 43874 25454
rect 34962 25342 34974 25394
rect 35026 25342 35038 25394
rect 13638 25282 13690 25294
rect 13638 25218 13690 25230
rect 20694 25282 20746 25294
rect 25554 25286 25566 25338
rect 25618 25286 25630 25338
rect 27458 25286 27470 25338
rect 27522 25286 27534 25338
rect 29766 25330 29818 25342
rect 42702 25330 42754 25342
rect 20694 25218 20746 25230
rect 1344 25114 44576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 44576 25114
rect 1344 25028 44576 25062
rect 13526 24946 13578 24958
rect 13526 24882 13578 24894
rect 37438 24946 37490 24958
rect 37438 24882 37490 24894
rect 42366 24946 42418 24958
rect 42366 24882 42418 24894
rect 19966 24834 20018 24846
rect 28634 24782 28646 24834
rect 28698 24782 28710 24834
rect 19966 24770 20018 24782
rect 13010 24697 13022 24749
rect 13074 24697 13086 24749
rect 14030 24722 14082 24734
rect 13346 24670 13358 24722
rect 13410 24670 13422 24722
rect 14030 24658 14082 24670
rect 17278 24722 17330 24734
rect 23762 24697 23774 24749
rect 23826 24697 23838 24749
rect 24782 24722 24834 24734
rect 17278 24658 17330 24670
rect 25442 24697 25454 24749
rect 25506 24697 25518 24749
rect 28142 24722 28194 24734
rect 24782 24658 24834 24670
rect 28142 24658 28194 24670
rect 28366 24722 28418 24734
rect 28366 24658 28418 24670
rect 29262 24722 29314 24734
rect 29262 24658 29314 24670
rect 29374 24722 29426 24734
rect 32498 24697 32510 24749
rect 32562 24697 32574 24749
rect 32958 24722 33010 24734
rect 29374 24658 29426 24670
rect 33730 24670 33742 24722
rect 33794 24670 33806 24722
rect 36082 24697 36094 24749
rect 36146 24697 36158 24749
rect 39118 24722 39170 24734
rect 39982 24670 39994 24722
rect 40046 24670 40058 24722
rect 41010 24697 41022 24749
rect 41074 24697 41086 24749
rect 44270 24722 44322 24734
rect 32958 24658 33010 24670
rect 39118 24658 39170 24670
rect 44270 24658 44322 24670
rect 14802 24558 14814 24610
rect 14866 24558 14878 24610
rect 16706 24558 16718 24610
rect 16770 24558 16782 24610
rect 18050 24558 18062 24610
rect 18114 24558 18126 24610
rect 35634 24558 35646 24610
rect 35698 24558 35710 24610
rect 11678 24498 11730 24510
rect 11678 24434 11730 24446
rect 22206 24498 22258 24510
rect 22206 24434 22258 24446
rect 24446 24498 24498 24510
rect 24446 24434 24498 24446
rect 26462 24498 26514 24510
rect 31502 24498 31554 24510
rect 29642 24446 29654 24498
rect 29706 24446 29718 24498
rect 26462 24434 26514 24446
rect 31502 24434 31554 24446
rect 40238 24498 40290 24510
rect 40238 24434 40290 24446
rect 43934 24498 43986 24510
rect 43934 24434 43986 24446
rect 1344 24330 44576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 44576 24330
rect 1344 24244 44576 24278
rect 11062 24162 11114 24174
rect 11062 24098 11114 24110
rect 19518 24162 19570 24174
rect 19518 24098 19570 24110
rect 10278 24050 10330 24062
rect 41022 24050 41074 24062
rect 11442 23998 11454 24050
rect 11506 23998 11518 24050
rect 12226 23998 12238 24050
rect 12290 23998 12302 24050
rect 15586 23998 15598 24050
rect 15650 23998 15662 24050
rect 16818 23998 16830 24050
rect 16882 23998 16894 24050
rect 18610 23998 18622 24050
rect 18674 23998 18686 24050
rect 21970 23998 21982 24050
rect 22034 23998 22046 24050
rect 23874 23998 23886 24050
rect 23938 23998 23950 24050
rect 25330 23998 25342 24050
rect 25394 23998 25406 24050
rect 30146 23998 30158 24050
rect 30210 23998 30222 24050
rect 33618 23998 33630 24050
rect 33682 23998 33694 24050
rect 35970 23998 35982 24050
rect 36034 23998 36046 24050
rect 10278 23986 10330 23998
rect 41022 23986 41074 23998
rect 19854 23938 19906 23950
rect 10782 23882 10834 23894
rect 10882 23886 10894 23938
rect 10946 23886 10958 23938
rect 11554 23842 11566 23894
rect 11618 23842 11630 23894
rect 11890 23886 11902 23938
rect 11954 23886 11966 23938
rect 12338 23871 12350 23923
rect 12402 23871 12414 23923
rect 12674 23886 12686 23938
rect 12738 23886 12750 23938
rect 15698 23871 15710 23923
rect 15762 23871 15774 23923
rect 16034 23886 16046 23938
rect 16098 23886 16110 23938
rect 16930 23871 16942 23923
rect 16994 23871 17006 23923
rect 17154 23886 17166 23938
rect 17218 23886 17230 23938
rect 18790 23908 18842 23920
rect 18946 23886 18958 23938
rect 19010 23886 19022 23938
rect 19854 23874 19906 23886
rect 21198 23938 21250 23950
rect 21198 23874 21250 23886
rect 24558 23938 24610 23950
rect 24558 23874 24610 23886
rect 28702 23938 28754 23950
rect 31838 23938 31890 23950
rect 28702 23874 28754 23886
rect 29138 23858 29150 23910
rect 29202 23858 29214 23910
rect 31838 23874 31890 23886
rect 32846 23938 32898 23950
rect 32846 23874 32898 23886
rect 35534 23938 35586 23950
rect 37550 23938 37602 23950
rect 39790 23938 39842 23950
rect 35534 23874 35586 23886
rect 36150 23908 36202 23920
rect 18790 23844 18842 23856
rect 36306 23886 36318 23938
rect 36370 23886 36382 23938
rect 38210 23886 38222 23938
rect 38274 23886 38286 23938
rect 37550 23874 37602 23886
rect 36150 23844 36202 23856
rect 10782 23818 10834 23830
rect 27246 23826 27298 23838
rect 37930 23830 37942 23882
rect 37994 23830 38006 23882
rect 27246 23762 27298 23774
rect 38670 23826 38722 23838
rect 38901 23830 38913 23882
rect 38965 23830 38977 23882
rect 39790 23874 39842 23886
rect 40350 23938 40402 23950
rect 40350 23874 40402 23886
rect 40686 23938 40738 23950
rect 40686 23874 40738 23886
rect 40910 23899 40962 23911
rect 41234 23886 41246 23938
rect 41298 23886 41310 23938
rect 41682 23858 41694 23910
rect 41746 23858 41758 23910
rect 40910 23835 40962 23847
rect 10614 23714 10666 23726
rect 10614 23650 10666 23662
rect 32174 23714 32226 23726
rect 37650 23718 37662 23770
rect 37714 23718 37726 23770
rect 38670 23762 38722 23774
rect 32174 23650 32226 23662
rect 43374 23714 43426 23726
rect 43374 23650 43426 23662
rect 1344 23546 44576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 44576 23546
rect 1344 23460 44576 23494
rect 32398 23378 32450 23390
rect 32398 23314 32450 23326
rect 33126 23378 33178 23390
rect 33126 23314 33178 23326
rect 33574 23378 33626 23390
rect 33574 23314 33626 23326
rect 27806 23266 27858 23278
rect 20582 23210 20634 23222
rect 21198 23210 21250 23222
rect 9650 23102 9662 23154
rect 9714 23102 9726 23154
rect 9874 23146 9886 23198
rect 9938 23146 9950 23198
rect 10546 23146 10558 23198
rect 10610 23146 10622 23198
rect 10882 23102 10894 23154
rect 10946 23102 10958 23154
rect 13682 23129 13694 23181
rect 13746 23129 13758 23181
rect 14478 23154 14530 23166
rect 14478 23090 14530 23102
rect 15710 23154 15762 23166
rect 15710 23090 15762 23102
rect 16830 23154 16882 23166
rect 20582 23146 20634 23158
rect 20862 23182 20914 23194
rect 21074 23158 21086 23210
rect 21138 23158 21150 23210
rect 31054 23266 31106 23278
rect 27806 23202 27858 23214
rect 28702 23210 28754 23222
rect 21198 23146 21250 23158
rect 20862 23118 20914 23130
rect 21746 23102 21758 23154
rect 21810 23102 21822 23154
rect 23986 23129 23998 23181
rect 24050 23129 24062 23181
rect 25118 23154 25170 23166
rect 28130 23102 28142 23154
rect 28194 23102 28206 23154
rect 28702 23146 28754 23158
rect 28814 23182 28866 23194
rect 28814 23118 28866 23130
rect 29038 23182 29090 23194
rect 29250 23158 29262 23210
rect 29314 23158 29326 23210
rect 31054 23202 31106 23214
rect 29038 23118 29090 23130
rect 29934 23154 29986 23166
rect 31390 23154 31442 23166
rect 30798 23102 30810 23154
rect 30862 23102 30874 23154
rect 16830 23090 16882 23102
rect 25118 23090 25170 23102
rect 29934 23090 29986 23102
rect 31390 23090 31442 23102
rect 32062 23154 32114 23166
rect 34862 23154 34914 23166
rect 36430 23154 36482 23166
rect 37550 23154 37602 23166
rect 33282 23102 33294 23154
rect 33346 23102 33358 23154
rect 33730 23102 33742 23154
rect 33794 23102 33806 23154
rect 35726 23102 35738 23154
rect 35790 23102 35802 23154
rect 37294 23102 37306 23154
rect 37358 23102 37370 23154
rect 37986 23102 37998 23154
rect 38050 23102 38062 23154
rect 38322 23129 38334 23181
rect 38386 23129 38398 23181
rect 38670 23154 38722 23166
rect 32062 23090 32114 23102
rect 34862 23090 34914 23102
rect 36430 23090 36482 23102
rect 37550 23090 37602 23102
rect 38670 23090 38722 23102
rect 39006 23154 39058 23166
rect 39006 23090 39058 23102
rect 39454 23154 39506 23166
rect 40450 23102 40462 23154
rect 40514 23102 40526 23154
rect 41010 23102 41022 23154
rect 41074 23102 41086 23154
rect 41346 23117 41358 23169
rect 41410 23117 41422 23169
rect 43038 23154 43090 23166
rect 42149 23102 42161 23154
rect 42213 23102 42225 23154
rect 43474 23146 43486 23198
rect 43538 23146 43550 23198
rect 43810 23102 43822 23154
rect 43874 23102 43886 23154
rect 39454 23090 39506 23102
rect 43038 23090 43090 23102
rect 9986 22990 9998 23042
rect 10050 22990 10062 23042
rect 10434 22990 10446 23042
rect 10498 22990 10510 23042
rect 25890 22990 25902 23042
rect 25954 22990 25966 23042
rect 28310 22986 28362 22998
rect 38098 22990 38110 23042
rect 38162 22990 38174 23042
rect 41458 22990 41470 23042
rect 41522 22990 41534 23042
rect 43362 22990 43374 23042
rect 43426 22990 43438 23042
rect 12686 22930 12738 22942
rect 12686 22866 12738 22878
rect 14142 22930 14194 22942
rect 14142 22866 14194 22878
rect 15374 22930 15426 22942
rect 15374 22866 15426 22878
rect 16494 22930 16546 22942
rect 20358 22930 20410 22942
rect 17490 22878 17502 22930
rect 17554 22927 17566 22930
rect 18274 22927 18286 22930
rect 17554 22881 18286 22927
rect 17554 22878 17566 22881
rect 18274 22878 18286 22881
rect 18338 22878 18350 22930
rect 28310 22922 28362 22934
rect 29542 22930 29594 22942
rect 16494 22866 16546 22878
rect 20358 22866 20410 22878
rect 29542 22866 29594 22878
rect 31726 22930 31778 22942
rect 31726 22866 31778 22878
rect 35982 22930 36034 22942
rect 35982 22866 36034 22878
rect 39790 22930 39842 22942
rect 39790 22866 39842 22878
rect 40294 22930 40346 22942
rect 40294 22866 40346 22878
rect 41918 22930 41970 22942
rect 41918 22866 41970 22878
rect 1344 22762 44576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 44576 22762
rect 1344 22676 44576 22710
rect 16158 22594 16210 22606
rect 16158 22530 16210 22542
rect 19630 22594 19682 22606
rect 19630 22530 19682 22542
rect 22654 22594 22706 22606
rect 22654 22530 22706 22542
rect 24446 22594 24498 22606
rect 24446 22530 24498 22542
rect 36206 22594 36258 22606
rect 36206 22530 36258 22542
rect 38110 22594 38162 22606
rect 38110 22530 38162 22542
rect 42926 22594 42978 22606
rect 42926 22530 42978 22542
rect 10882 22430 10894 22482
rect 10946 22430 10958 22482
rect 12786 22430 12798 22482
rect 12850 22430 12862 22482
rect 26226 22430 26238 22482
rect 26290 22430 26302 22482
rect 27682 22430 27694 22482
rect 27746 22430 27758 22482
rect 29138 22430 29150 22482
rect 29202 22430 29214 22482
rect 38658 22430 38670 22482
rect 38722 22430 38734 22482
rect 10110 22370 10162 22382
rect 9762 22290 9774 22342
rect 9826 22290 9838 22342
rect 10110 22306 10162 22318
rect 13582 22370 13634 22382
rect 20750 22370 20802 22382
rect 13582 22306 13634 22318
rect 14446 22262 14458 22314
rect 14510 22262 14522 22314
rect 15138 22290 15150 22342
rect 15202 22290 15214 22342
rect 19861 22318 19873 22370
rect 19925 22318 19937 22370
rect 20750 22306 20802 22318
rect 22318 22370 22370 22382
rect 27470 22370 27522 22382
rect 29934 22370 29986 22382
rect 31950 22370 32002 22382
rect 22318 22306 22370 22318
rect 23538 22290 23550 22342
rect 23602 22290 23614 22342
rect 26338 22274 26350 22326
rect 26402 22274 26414 22326
rect 26674 22318 26686 22370
rect 26738 22318 26750 22370
rect 27470 22306 27522 22318
rect 27750 22340 27802 22352
rect 28018 22318 28030 22370
rect 28082 22318 28094 22370
rect 27750 22276 27802 22288
rect 29250 22274 29262 22326
rect 29314 22274 29326 22326
rect 29586 22318 29598 22370
rect 29650 22318 29662 22370
rect 30798 22318 30810 22370
rect 30862 22318 30874 22370
rect 29934 22306 29986 22318
rect 31950 22306 32002 22318
rect 34190 22370 34242 22382
rect 34190 22306 34242 22318
rect 35086 22370 35138 22382
rect 35086 22306 35138 22318
rect 36990 22370 37042 22382
rect 39230 22370 39282 22382
rect 38546 22318 38558 22370
rect 38610 22318 38622 22370
rect 14702 22258 14754 22270
rect 14702 22194 14754 22206
rect 31054 22258 31106 22270
rect 35950 22262 35962 22314
rect 36014 22262 36026 22314
rect 36990 22306 37042 22318
rect 37854 22262 37866 22314
rect 37918 22262 37930 22314
rect 38826 22262 38838 22314
rect 38890 22262 38902 22314
rect 39230 22306 39282 22318
rect 39678 22370 39730 22382
rect 44046 22370 44098 22382
rect 40450 22318 40462 22370
rect 40514 22318 40526 22370
rect 39678 22306 39730 22318
rect 31054 22194 31106 22206
rect 42366 22258 42418 22270
rect 43157 22262 43169 22314
rect 43221 22262 43233 22314
rect 44046 22306 44098 22318
rect 42366 22194 42418 22206
rect 8430 22146 8482 22158
rect 8430 22082 8482 22094
rect 27134 22146 27186 22158
rect 27134 22082 27186 22094
rect 28646 22146 28698 22158
rect 28646 22082 28698 22094
rect 31614 22146 31666 22158
rect 31614 22082 31666 22094
rect 32342 22146 32394 22158
rect 32342 22082 32394 22094
rect 33854 22146 33906 22158
rect 33854 22082 33906 22094
rect 1344 21978 44576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 44576 21978
rect 1344 21892 44576 21926
rect 17950 21810 18002 21822
rect 17950 21746 18002 21758
rect 19294 21810 19346 21822
rect 19294 21746 19346 21758
rect 32006 21810 32058 21822
rect 28466 21702 28478 21754
rect 28530 21702 28542 21754
rect 32006 21746 32058 21758
rect 29206 21698 29258 21710
rect 29206 21634 29258 21646
rect 37774 21698 37826 21710
rect 8542 21586 8594 21598
rect 8082 21534 8094 21586
rect 8146 21534 8158 21586
rect 8542 21522 8594 21534
rect 9438 21586 9490 21598
rect 12574 21586 12626 21598
rect 16942 21586 16994 21598
rect 10210 21534 10222 21586
rect 10274 21534 10286 21586
rect 13438 21534 13450 21586
rect 13502 21534 13514 21586
rect 16146 21534 16158 21586
rect 16210 21534 16222 21586
rect 9438 21522 9490 21534
rect 12574 21522 12626 21534
rect 16942 21522 16994 21534
rect 17614 21586 17666 21598
rect 17614 21522 17666 21534
rect 18398 21586 18450 21598
rect 18398 21522 18450 21534
rect 19630 21586 19682 21598
rect 21086 21586 21138 21598
rect 20197 21534 20209 21586
rect 20261 21534 20273 21586
rect 19630 21522 19682 21534
rect 21086 21522 21138 21534
rect 24110 21586 24162 21598
rect 24110 21522 24162 21534
rect 24334 21586 24386 21598
rect 25442 21561 25454 21613
rect 25506 21561 25518 21613
rect 28354 21578 28366 21630
rect 28418 21578 28430 21630
rect 29486 21586 29538 21598
rect 29754 21590 29766 21642
rect 29818 21590 29830 21642
rect 37774 21634 37826 21646
rect 43822 21698 43874 21710
rect 43822 21634 43874 21646
rect 29934 21586 29986 21598
rect 28690 21534 28702 21586
rect 28754 21534 28766 21586
rect 29586 21534 29598 21586
rect 29650 21534 29662 21586
rect 30370 21534 30382 21586
rect 30434 21534 30446 21586
rect 31110 21572 31122 21624
rect 31174 21572 31186 21624
rect 32958 21586 33010 21598
rect 40462 21586 40514 21598
rect 39666 21534 39678 21586
rect 39730 21534 39742 21586
rect 24334 21522 24386 21534
rect 29486 21522 29538 21534
rect 29934 21522 29986 21534
rect 32958 21522 33010 21534
rect 40462 21522 40514 21534
rect 41134 21586 41186 21598
rect 41134 21522 41186 21534
rect 31558 21474 31610 21486
rect 8262 21418 8314 21430
rect 12114 21422 12126 21474
rect 12178 21422 12190 21474
rect 14242 21422 14254 21474
rect 14306 21422 14318 21474
rect 26450 21422 26462 21474
rect 26514 21422 26526 21474
rect 33730 21422 33742 21474
rect 33794 21422 33806 21474
rect 35634 21422 35646 21474
rect 35698 21422 35710 21474
rect 41906 21422 41918 21474
rect 41970 21422 41982 21474
rect 8262 21354 8314 21366
rect 8878 21362 8930 21374
rect 8878 21298 8930 21310
rect 13694 21362 13746 21374
rect 13694 21298 13746 21310
rect 18734 21362 18786 21374
rect 18734 21298 18786 21310
rect 19966 21362 20018 21374
rect 30594 21366 30606 21418
rect 30658 21366 30670 21418
rect 31558 21410 31610 21422
rect 23818 21310 23830 21362
rect 23882 21310 23894 21362
rect 19966 21298 20018 21310
rect 1344 21194 44576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 44576 21194
rect 1344 21108 44576 21142
rect 18268 21026 18320 21038
rect 18268 20962 18320 20974
rect 25398 21026 25450 21038
rect 25398 20962 25450 20974
rect 29374 21026 29426 21038
rect 29374 20962 29426 20974
rect 32062 21026 32114 21038
rect 21404 20914 21456 20926
rect 12226 20862 12238 20914
rect 12290 20862 12302 20914
rect 19014 20858 19066 20870
rect 8990 20802 9042 20814
rect 8194 20750 8206 20802
rect 8258 20750 8270 20802
rect 8990 20738 9042 20750
rect 9102 20802 9154 20814
rect 13582 20802 13634 20814
rect 17950 20802 18002 20814
rect 9874 20750 9886 20802
rect 9938 20750 9950 20802
rect 9102 20738 9154 20750
rect 12338 20706 12350 20758
rect 12402 20706 12414 20758
rect 12562 20750 12574 20802
rect 12626 20750 12638 20802
rect 14446 20750 14458 20802
rect 14510 20750 14522 20802
rect 17154 20750 17166 20802
rect 17218 20750 17230 20802
rect 13582 20738 13634 20750
rect 17950 20738 18002 20750
rect 18510 20802 18562 20814
rect 22822 20914 22874 20926
rect 30706 20918 30718 20970
rect 30770 20918 30782 20970
rect 32062 20962 32114 20974
rect 42254 21026 42306 21038
rect 42254 20962 42306 20974
rect 39360 20914 39412 20926
rect 21404 20850 21456 20862
rect 22150 20858 22202 20870
rect 19014 20794 19066 20806
rect 20862 20802 20914 20814
rect 18510 20738 18562 20750
rect 20862 20738 20914 20750
rect 21646 20802 21698 20814
rect 22822 20850 22874 20862
rect 24838 20858 24890 20870
rect 26898 20862 26910 20914
rect 26962 20862 26974 20914
rect 28130 20862 28142 20914
rect 28194 20862 28206 20914
rect 33282 20862 33294 20914
rect 33346 20862 33358 20914
rect 35186 20862 35198 20914
rect 35250 20862 35262 20914
rect 22150 20794 22202 20806
rect 24670 20802 24722 20814
rect 21646 20738 21698 20750
rect 38614 20858 38666 20870
rect 24838 20794 24890 20806
rect 25118 20802 25170 20814
rect 24670 20738 24722 20750
rect 25118 20738 25170 20750
rect 26574 20802 26626 20814
rect 29710 20802 29762 20814
rect 26574 20738 26626 20750
rect 27010 20706 27022 20758
rect 27074 20706 27086 20758
rect 27234 20750 27246 20802
rect 27298 20750 27310 20802
rect 27682 20750 27694 20802
rect 27746 20750 27758 20802
rect 28018 20706 28030 20758
rect 28082 20706 28094 20758
rect 29710 20738 29762 20750
rect 29934 20802 29986 20814
rect 32398 20802 32450 20814
rect 30482 20750 30494 20802
rect 30546 20750 30558 20802
rect 29934 20738 29986 20750
rect 32398 20738 32450 20750
rect 32510 20802 32562 20814
rect 39360 20850 39412 20862
rect 40630 20858 40682 20870
rect 38614 20794 38666 20806
rect 39118 20802 39170 20814
rect 32510 20738 32562 20750
rect 39118 20738 39170 20750
rect 40126 20802 40178 20814
rect 43654 20858 43706 20870
rect 40630 20794 40682 20806
rect 41302 20802 41354 20814
rect 40126 20738 40178 20750
rect 41302 20738 41354 20750
rect 42590 20802 42642 20814
rect 42590 20738 42642 20750
rect 42908 20802 42960 20814
rect 42908 20738 42960 20750
rect 43150 20802 43202 20814
rect 43654 20794 43706 20806
rect 43150 20738 43202 20750
rect 6302 20690 6354 20702
rect 6302 20626 6354 20638
rect 11790 20690 11842 20702
rect 11790 20626 11842 20638
rect 14702 20690 14754 20702
rect 14702 20626 14754 20638
rect 15262 20690 15314 20702
rect 15262 20626 15314 20638
rect 19182 20690 19234 20702
rect 19182 20626 19234 20638
rect 22318 20690 22370 20702
rect 22318 20626 22370 20638
rect 25006 20690 25058 20702
rect 25006 20626 25058 20638
rect 39884 20690 39936 20702
rect 19686 20578 19738 20590
rect 19686 20514 19738 20526
rect 20526 20578 20578 20590
rect 20526 20514 20578 20526
rect 28646 20578 28698 20590
rect 28646 20514 28698 20526
rect 31334 20578 31386 20590
rect 31334 20514 31386 20526
rect 35814 20578 35866 20590
rect 38770 20582 38782 20634
rect 38834 20582 38846 20634
rect 39884 20626 39936 20638
rect 40798 20690 40850 20702
rect 40798 20626 40850 20638
rect 35814 20514 35866 20526
rect 41862 20578 41914 20590
rect 43586 20582 43598 20634
rect 43650 20582 43662 20634
rect 41862 20514 41914 20526
rect 1344 20410 44576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 44576 20410
rect 1344 20324 44576 20358
rect 13358 20242 13410 20254
rect 13358 20178 13410 20190
rect 17614 20242 17666 20254
rect 17614 20178 17666 20190
rect 25342 20242 25394 20254
rect 25342 20178 25394 20190
rect 12126 20130 12178 20142
rect 12126 20066 12178 20078
rect 15822 20130 15874 20142
rect 15822 20066 15874 20078
rect 21870 20130 21922 20142
rect 28354 20134 28366 20186
rect 28418 20134 28430 20186
rect 29934 20130 29986 20142
rect 26842 20078 26854 20130
rect 26906 20078 26918 20130
rect 21870 20066 21922 20078
rect 28702 20057 28754 20069
rect 29934 20066 29986 20078
rect 33164 20130 33216 20142
rect 33164 20066 33216 20078
rect 34508 20130 34560 20142
rect 35074 20134 35086 20186
rect 35138 20134 35150 20186
rect 8418 19981 8430 20033
rect 8482 19981 8494 20033
rect 9438 20018 9490 20030
rect 8754 19966 8766 20018
rect 8818 19966 8830 20018
rect 10210 19966 10222 20018
rect 10274 19966 10286 20018
rect 14690 19993 14702 20045
rect 14754 19993 14766 20045
rect 16494 20018 16546 20030
rect 9438 19954 9490 19966
rect 15990 19962 16042 19974
rect 8038 19906 8090 19918
rect 16494 19954 16546 19966
rect 16736 20018 16788 20030
rect 16736 19954 16788 19966
rect 17278 20018 17330 20030
rect 17278 19954 17330 19966
rect 19182 20018 19234 20030
rect 22206 20018 22258 20030
rect 19954 19966 19966 20018
rect 20018 19966 20030 20018
rect 19182 19954 19234 19966
rect 22206 19954 22258 19966
rect 24278 20018 24330 20030
rect 24278 19954 24330 19966
rect 25678 20018 25730 20030
rect 25678 19954 25730 19966
rect 26350 20018 26402 20030
rect 26350 19954 26402 19966
rect 27134 20018 27186 20030
rect 27134 19954 27186 19966
rect 27358 20018 27410 20030
rect 27458 19966 27470 20018
rect 27522 19966 27534 20018
rect 28242 19966 28254 20018
rect 28306 19966 28318 20018
rect 28702 19993 28754 20005
rect 28926 20018 28978 20030
rect 27358 19954 27410 19966
rect 28926 19954 28978 19966
rect 30270 20018 30322 20030
rect 33406 20018 33458 20030
rect 33898 20022 33910 20074
rect 33962 20022 33974 20074
rect 34508 20066 34560 20078
rect 40238 20130 40290 20142
rect 30706 19966 30718 20018
rect 30770 19966 30782 20018
rect 31378 19966 31390 20018
rect 31442 19966 31454 20018
rect 30270 19954 30322 19966
rect 33406 19954 33458 19966
rect 34078 20018 34130 20030
rect 34078 19954 34130 19966
rect 34750 20018 34802 20030
rect 35242 20022 35254 20074
rect 35306 20022 35318 20074
rect 40238 20066 40290 20078
rect 34750 19954 34802 19966
rect 38670 20018 38722 20030
rect 38670 19954 38722 19966
rect 39902 20018 39954 20030
rect 39902 19954 39954 19966
rect 40798 20018 40850 20030
rect 40798 19954 40850 19966
rect 41694 20018 41746 20030
rect 41694 19954 41746 19966
rect 42926 20018 42978 20030
rect 42926 19954 42978 19966
rect 43038 20018 43090 20030
rect 43038 19954 43090 19966
rect 43710 20018 43762 20030
rect 43710 19954 43762 19966
rect 8306 19854 8318 19906
rect 8370 19854 8382 19906
rect 15990 19898 16042 19910
rect 24726 19906 24778 19918
rect 44046 19906 44098 19918
rect 35970 19854 35982 19906
rect 36034 19854 36046 19906
rect 37874 19854 37886 19906
rect 37938 19854 37950 19906
rect 8038 19842 8090 19854
rect 24726 19842 24778 19854
rect 44046 19842 44098 19854
rect 22542 19794 22594 19806
rect 22542 19730 22594 19742
rect 26014 19794 26066 19806
rect 26014 19730 26066 19742
rect 27638 19794 27690 19806
rect 41134 19794 41186 19806
rect 31714 19742 31726 19794
rect 31778 19742 31790 19794
rect 27638 19730 27690 19742
rect 41134 19730 41186 19742
rect 42030 19794 42082 19806
rect 42030 19730 42082 19742
rect 42590 19794 42642 19806
rect 42590 19730 42642 19742
rect 43374 19794 43426 19806
rect 43374 19730 43426 19742
rect 1344 19626 44576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 44576 19626
rect 1344 19540 44576 19574
rect 9774 19458 9826 19470
rect 9774 19394 9826 19406
rect 22224 19458 22276 19470
rect 35870 19458 35922 19470
rect 26954 19406 26966 19458
rect 27018 19406 27030 19458
rect 22224 19394 22276 19406
rect 13806 19346 13858 19358
rect 13806 19282 13858 19294
rect 22822 19346 22874 19358
rect 22822 19282 22874 19294
rect 23494 19346 23546 19358
rect 29474 19350 29486 19402
rect 29538 19350 29550 19402
rect 35870 19394 35922 19406
rect 38558 19458 38610 19470
rect 38558 19394 38610 19406
rect 39772 19458 39824 19470
rect 39772 19394 39824 19406
rect 23494 19282 23546 19294
rect 35198 19346 35250 19358
rect 44214 19346 44266 19358
rect 35198 19282 35250 19294
rect 37158 19290 37210 19302
rect 11678 19234 11730 19246
rect 14142 19234 14194 19246
rect 8530 19182 8542 19234
rect 8594 19182 8606 19234
rect 9090 19154 9102 19206
rect 9154 19154 9166 19206
rect 12542 19182 12554 19234
rect 12606 19182 12618 19234
rect 13458 19182 13470 19234
rect 13522 19182 13534 19234
rect 11678 19170 11730 19182
rect 12798 19122 12850 19134
rect 13794 19126 13806 19178
rect 13858 19126 13870 19178
rect 14142 19170 14194 19182
rect 14478 19234 14530 19246
rect 15710 19234 15762 19246
rect 15026 19182 15038 19234
rect 15090 19182 15102 19234
rect 14478 19170 14530 19182
rect 15362 19126 15374 19178
rect 15426 19126 15438 19178
rect 15710 19170 15762 19182
rect 21478 19234 21530 19246
rect 21478 19170 21530 19182
rect 21982 19234 22034 19246
rect 21982 19170 22034 19182
rect 23774 19234 23826 19246
rect 27246 19234 27298 19246
rect 24546 19182 24558 19234
rect 24610 19182 24622 19234
rect 23774 19170 23826 19182
rect 27246 19170 27298 19182
rect 27470 19234 27522 19246
rect 34190 19234 34242 19246
rect 27794 19182 27806 19234
rect 27858 19182 27870 19234
rect 27470 19170 27522 19182
rect 28018 19138 28030 19190
rect 28082 19138 28094 19190
rect 29138 19182 29150 19234
rect 29202 19182 29214 19234
rect 29474 19182 29486 19234
rect 29538 19182 29550 19234
rect 34190 19170 34242 19182
rect 34862 19234 34914 19246
rect 34862 19170 34914 19182
rect 35534 19234 35586 19246
rect 40518 19290 40570 19302
rect 43586 19294 43598 19346
rect 43650 19294 43662 19346
rect 37158 19226 37210 19238
rect 37662 19234 37714 19246
rect 35534 19170 35586 19182
rect 37662 19170 37714 19182
rect 37904 19234 37956 19246
rect 37904 19170 37956 19182
rect 38222 19234 38274 19246
rect 38222 19170 38274 19182
rect 40014 19234 40066 19246
rect 44214 19282 44266 19294
rect 40518 19226 40570 19238
rect 40910 19234 40962 19246
rect 40014 19170 40066 19182
rect 41682 19182 41694 19234
rect 41746 19182 41758 19234
rect 40910 19170 40962 19182
rect 8374 19066 8426 19078
rect 12798 19058 12850 19070
rect 21310 19122 21362 19134
rect 15586 19014 15598 19066
rect 15650 19014 15662 19066
rect 21310 19058 21362 19070
rect 26462 19122 26514 19134
rect 26462 19058 26514 19070
rect 36990 19122 37042 19134
rect 8374 19002 8426 19014
rect 17110 19010 17162 19022
rect 27906 19014 27918 19066
rect 27970 19014 27982 19066
rect 36990 19058 37042 19070
rect 40686 19122 40738 19134
rect 40686 19058 40738 19070
rect 17110 18946 17162 18958
rect 28646 19010 28698 19022
rect 28646 18946 28698 18958
rect 34022 19010 34074 19022
rect 34022 18946 34074 18958
rect 34526 19010 34578 19022
rect 34526 18946 34578 18958
rect 1344 18842 44576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 44576 18842
rect 1344 18756 44576 18790
rect 18398 18562 18450 18574
rect 8866 18425 8878 18477
rect 8930 18425 8942 18477
rect 9874 18398 9886 18450
rect 9938 18398 9950 18450
rect 10210 18413 10222 18465
rect 10274 18413 10286 18465
rect 10434 18398 10446 18450
rect 10498 18398 10510 18450
rect 10994 18442 11006 18494
rect 11058 18442 11070 18494
rect 11218 18398 11230 18450
rect 11282 18398 11294 18450
rect 12002 18398 12014 18450
rect 12066 18398 12078 18450
rect 13906 18425 13918 18477
rect 13970 18425 13982 18477
rect 14914 18454 14926 18506
rect 14978 18454 14990 18506
rect 18398 18498 18450 18510
rect 21758 18562 21810 18574
rect 21758 18498 21810 18510
rect 28030 18489 28082 18501
rect 15262 18450 15314 18462
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 15262 18386 15314 18398
rect 16942 18450 16994 18462
rect 16942 18386 16994 18398
rect 17484 18450 17536 18462
rect 17484 18386 17536 18398
rect 17726 18450 17778 18462
rect 19070 18450 19122 18462
rect 22206 18450 22258 18462
rect 17726 18386 17778 18398
rect 18230 18394 18282 18406
rect 14926 18338 14978 18350
rect 9718 18282 9770 18294
rect 10098 18286 10110 18338
rect 10162 18286 10174 18338
rect 10882 18286 10894 18338
rect 10946 18286 10958 18338
rect 19842 18398 19854 18450
rect 19906 18398 19918 18450
rect 22878 18450 22930 18462
rect 19070 18386 19122 18398
rect 22206 18386 22258 18398
rect 22374 18394 22426 18406
rect 18230 18330 18282 18342
rect 18902 18338 18954 18350
rect 7982 18226 8034 18238
rect 14926 18274 14978 18286
rect 22878 18386 22930 18398
rect 23998 18450 24050 18462
rect 24670 18450 24722 18462
rect 23998 18386 24050 18398
rect 24502 18394 24554 18406
rect 22374 18330 22426 18342
rect 23756 18338 23808 18350
rect 18902 18274 18954 18286
rect 24670 18386 24722 18398
rect 25118 18450 25170 18462
rect 25118 18386 25170 18398
rect 25454 18450 25506 18462
rect 27022 18450 27074 18462
rect 26562 18398 26574 18450
rect 26626 18398 26638 18450
rect 25454 18386 25506 18398
rect 27022 18386 27074 18398
rect 27806 18450 27858 18462
rect 28030 18425 28082 18437
rect 28466 18398 28478 18450
rect 28530 18398 28542 18450
rect 28802 18398 28814 18450
rect 28866 18398 28878 18450
rect 29138 18413 29150 18465
rect 29202 18413 29214 18465
rect 30046 18450 30098 18462
rect 27806 18386 27858 18398
rect 30046 18386 30098 18398
rect 30270 18450 30322 18462
rect 33518 18450 33570 18462
rect 36206 18450 36258 18462
rect 31378 18398 31390 18450
rect 31442 18398 31454 18450
rect 32050 18398 32062 18450
rect 32114 18398 32126 18450
rect 34290 18398 34302 18450
rect 34354 18398 34366 18450
rect 30270 18386 30322 18398
rect 33518 18386 33570 18398
rect 36206 18386 36258 18398
rect 39454 18450 39506 18462
rect 39454 18386 39506 18398
rect 39790 18450 39842 18462
rect 39790 18386 39842 18398
rect 40126 18450 40178 18462
rect 40126 18386 40178 18398
rect 40798 18450 40850 18462
rect 43486 18450 43538 18462
rect 41570 18398 41582 18450
rect 41634 18398 41646 18450
rect 40798 18386 40850 18398
rect 43486 18386 43538 18398
rect 44214 18450 44266 18462
rect 44214 18386 44266 18398
rect 24502 18330 24554 18342
rect 26786 18286 26798 18338
rect 26850 18286 26862 18338
rect 28242 18286 28254 18338
rect 28306 18286 28318 18338
rect 29250 18286 29262 18338
rect 29314 18286 29326 18338
rect 36754 18286 36766 18338
rect 36818 18286 36830 18338
rect 38658 18286 38670 18338
rect 38722 18286 38734 18338
rect 23756 18274 23808 18286
rect 9718 18218 9770 18230
rect 16606 18226 16658 18238
rect 7982 18162 8034 18174
rect 16606 18162 16658 18174
rect 23120 18226 23172 18238
rect 30538 18174 30550 18226
rect 30602 18174 30614 18226
rect 32386 18174 32398 18226
rect 32450 18174 32462 18226
rect 23120 18162 23172 18174
rect 1344 18058 44576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 44576 18058
rect 1344 17972 44576 18006
rect 12686 17890 12738 17902
rect 12686 17826 12738 17838
rect 14590 17890 14642 17902
rect 14590 17826 14642 17838
rect 19070 17890 19122 17902
rect 28366 17890 28418 17902
rect 34060 17890 34112 17902
rect 19070 17826 19122 17838
rect 23662 17834 23714 17846
rect 21870 17778 21922 17790
rect 8306 17726 8318 17778
rect 8370 17726 8382 17778
rect 10210 17726 10222 17778
rect 10274 17726 10286 17778
rect 23662 17770 23714 17782
rect 24446 17834 24498 17846
rect 29866 17838 29878 17890
rect 29930 17838 29942 17890
rect 30650 17838 30662 17890
rect 30714 17838 30726 17890
rect 28366 17826 28418 17838
rect 31838 17834 31890 17846
rect 24446 17770 24498 17782
rect 25342 17778 25394 17790
rect 21870 17714 21922 17726
rect 25342 17714 25394 17726
rect 27582 17778 27634 17790
rect 32274 17782 32286 17834
rect 32338 17782 32350 17834
rect 34060 17826 34112 17838
rect 37214 17890 37266 17902
rect 37214 17826 37266 17838
rect 31838 17770 31890 17782
rect 43934 17778 43986 17790
rect 27582 17714 27634 17726
rect 34806 17722 34858 17734
rect 7534 17666 7586 17678
rect 7534 17602 7586 17614
rect 11566 17666 11618 17678
rect 11566 17602 11618 17614
rect 13470 17666 13522 17678
rect 15822 17666 15874 17678
rect 18510 17666 18562 17678
rect 14334 17614 14346 17666
rect 14398 17614 14410 17666
rect 16594 17614 16606 17666
rect 16658 17614 16670 17666
rect 12430 17558 12442 17610
rect 12494 17558 12506 17610
rect 13470 17602 13522 17614
rect 15822 17602 15874 17614
rect 18510 17602 18562 17614
rect 19406 17666 19458 17678
rect 19406 17602 19458 17614
rect 20862 17666 20914 17678
rect 20862 17602 20914 17614
rect 21534 17666 21586 17678
rect 27246 17666 27298 17678
rect 28702 17666 28754 17678
rect 22194 17614 22206 17666
rect 22258 17614 22270 17666
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 24098 17614 24110 17666
rect 24162 17614 24174 17666
rect 24546 17614 24558 17666
rect 24610 17614 24622 17666
rect 24882 17614 24894 17666
rect 24946 17614 24958 17666
rect 25442 17614 25454 17666
rect 25506 17614 25518 17666
rect 26114 17614 26126 17666
rect 26178 17614 26190 17666
rect 27906 17614 27918 17666
rect 27970 17614 27982 17666
rect 21534 17602 21586 17614
rect 21914 17558 21926 17610
rect 21978 17558 21990 17610
rect 27246 17602 27298 17614
rect 27458 17558 27470 17610
rect 27522 17558 27534 17610
rect 28702 17602 28754 17614
rect 29374 17666 29426 17678
rect 29374 17602 29426 17614
rect 29598 17666 29650 17678
rect 29598 17602 29650 17614
rect 30158 17666 30210 17678
rect 30158 17602 30210 17614
rect 30382 17666 30434 17678
rect 32846 17666 32898 17678
rect 31378 17614 31390 17666
rect 31442 17614 31454 17666
rect 31714 17614 31726 17666
rect 31778 17614 31790 17666
rect 32162 17614 32174 17666
rect 32226 17614 32238 17666
rect 32498 17614 32510 17666
rect 32562 17614 32574 17666
rect 30382 17602 30434 17614
rect 32846 17602 32898 17614
rect 34302 17666 34354 17678
rect 35590 17722 35642 17734
rect 40114 17726 40126 17778
rect 40178 17726 40190 17778
rect 42018 17726 42030 17778
rect 42082 17726 42094 17778
rect 34806 17658 34858 17670
rect 34974 17666 35026 17678
rect 34302 17602 34354 17614
rect 34974 17602 35026 17614
rect 35422 17666 35474 17678
rect 43318 17722 43370 17734
rect 35590 17658 35642 17670
rect 36094 17666 36146 17678
rect 35422 17602 35474 17614
rect 36094 17602 36146 17614
rect 36336 17666 36388 17678
rect 36336 17602 36388 17614
rect 36878 17666 36930 17678
rect 36878 17602 36930 17614
rect 39342 17666 39394 17678
rect 39342 17602 39394 17614
rect 42814 17666 42866 17678
rect 43934 17714 43986 17726
rect 43318 17658 43370 17670
rect 44270 17666 44322 17678
rect 42814 17602 42866 17614
rect 44270 17602 44322 17614
rect 42572 17554 42624 17566
rect 42572 17490 42624 17502
rect 20526 17442 20578 17454
rect 20526 17378 20578 17390
rect 33182 17442 33234 17454
rect 43138 17446 43150 17498
rect 43202 17446 43214 17498
rect 33182 17378 33234 17390
rect 1344 17274 44576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 44576 17274
rect 1344 17188 44576 17222
rect 8262 17106 8314 17118
rect 8262 17042 8314 17054
rect 8934 17106 8986 17118
rect 8934 17042 8986 17054
rect 16102 17106 16154 17118
rect 16102 17042 16154 17054
rect 16606 17106 16658 17118
rect 16606 17042 16658 17054
rect 34806 17106 34858 17118
rect 34806 17042 34858 17054
rect 35198 17106 35250 17118
rect 35198 17042 35250 17054
rect 35982 17106 36034 17118
rect 35982 17042 36034 17054
rect 40126 17106 40178 17118
rect 40126 17042 40178 17054
rect 41078 17106 41130 17118
rect 41078 17042 41130 17054
rect 42926 17106 42978 17118
rect 42926 17042 42978 17054
rect 43542 17106 43594 17118
rect 43542 17042 43594 17054
rect 43934 17106 43986 17118
rect 43934 17042 43986 17054
rect 18398 16994 18450 17006
rect 9438 16882 9490 16894
rect 8418 16830 8430 16882
rect 8482 16830 8494 16882
rect 9090 16830 9102 16882
rect 9154 16830 9166 16882
rect 9438 16818 9490 16830
rect 12126 16882 12178 16894
rect 12674 16857 12686 16909
rect 12738 16857 12750 16909
rect 16942 16882 16994 16894
rect 12126 16818 12178 16830
rect 16942 16818 16994 16830
rect 17484 16882 17536 16894
rect 17484 16818 17536 16830
rect 17726 16882 17778 16894
rect 18218 16886 18230 16938
rect 18282 16886 18294 16938
rect 18398 16930 18450 16942
rect 22430 16994 22482 17006
rect 22430 16930 22482 16942
rect 41452 16994 41504 17006
rect 17726 16818 17778 16830
rect 19742 16882 19794 16894
rect 23438 16882 23490 16894
rect 20514 16830 20526 16882
rect 20578 16830 20590 16882
rect 19742 16818 19794 16830
rect 23438 16818 23490 16830
rect 23756 16882 23808 16894
rect 23756 16818 23808 16830
rect 23998 16882 24050 16894
rect 24490 16886 24502 16938
rect 24554 16886 24566 16938
rect 23998 16818 24050 16830
rect 24670 16882 24722 16894
rect 26014 16882 26066 16894
rect 25778 16830 25790 16882
rect 25842 16830 25854 16882
rect 24670 16818 24722 16830
rect 26014 16818 26066 16830
rect 26910 16882 26962 16894
rect 26910 16818 26962 16830
rect 27246 16882 27298 16894
rect 27455 16869 27467 16921
rect 27519 16869 27531 16921
rect 29486 16882 29538 16894
rect 29810 16886 29822 16938
rect 29874 16886 29886 16938
rect 31838 16921 31890 16933
rect 41452 16930 41504 16942
rect 42366 16994 42418 17006
rect 31614 16882 31666 16894
rect 28466 16830 28478 16882
rect 28530 16830 28542 16882
rect 30146 16830 30158 16882
rect 30210 16830 30222 16882
rect 30482 16830 30494 16882
rect 30546 16830 30558 16882
rect 30818 16830 30830 16882
rect 30882 16830 30894 16882
rect 35534 16882 35586 16894
rect 31838 16857 31890 16869
rect 32274 16830 32286 16882
rect 32338 16830 32350 16882
rect 27246 16818 27298 16830
rect 29486 16818 29538 16830
rect 31614 16818 31666 16830
rect 35534 16818 35586 16830
rect 35646 16882 35698 16894
rect 35646 16818 35698 16830
rect 39678 16882 39730 16894
rect 39678 16818 39730 16830
rect 39790 16882 39842 16894
rect 39790 16818 39842 16830
rect 41694 16882 41746 16894
rect 42186 16886 42198 16938
rect 42250 16886 42262 16938
rect 42366 16930 42418 16942
rect 41694 16818 41746 16830
rect 42590 16882 42642 16894
rect 42590 16818 42642 16830
rect 44270 16882 44322 16894
rect 44270 16818 44322 16830
rect 27806 16770 27858 16782
rect 31950 16770 32002 16782
rect 10210 16718 10222 16770
rect 10274 16718 10286 16770
rect 25890 16718 25902 16770
rect 25954 16718 25966 16770
rect 29922 16718 29934 16770
rect 29986 16718 29998 16770
rect 27806 16706 27858 16718
rect 13582 16658 13634 16670
rect 13582 16594 13634 16606
rect 23102 16658 23154 16670
rect 30818 16662 30830 16714
rect 30882 16662 30894 16714
rect 31950 16706 32002 16718
rect 23102 16594 23154 16606
rect 39342 16658 39394 16670
rect 39342 16594 39394 16606
rect 1344 16490 44576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 44576 16490
rect 1344 16404 44576 16438
rect 12798 16322 12850 16334
rect 28534 16322 28586 16334
rect 26282 16270 26294 16322
rect 26346 16270 26358 16322
rect 12798 16258 12850 16270
rect 27022 16266 27074 16278
rect 31950 16322 32002 16334
rect 28534 16258 28586 16270
rect 31502 16266 31554 16278
rect 16146 16158 16158 16210
rect 16210 16158 16222 16210
rect 23650 16158 23662 16210
rect 23714 16158 23726 16210
rect 25554 16158 25566 16210
rect 25618 16158 25630 16210
rect 27022 16202 27074 16214
rect 31950 16258 32002 16270
rect 33742 16322 33794 16334
rect 33742 16258 33794 16270
rect 37662 16322 37714 16334
rect 37662 16258 37714 16270
rect 29586 16158 29598 16210
rect 29650 16158 29662 16210
rect 29922 16158 29934 16210
rect 29986 16158 29998 16210
rect 31502 16202 31554 16214
rect 40294 16210 40346 16222
rect 40294 16146 40346 16158
rect 43542 16210 43594 16222
rect 43542 16146 43594 16158
rect 44214 16210 44266 16222
rect 44214 16146 44266 16158
rect 7870 16098 7922 16110
rect 11454 16098 11506 16110
rect 8642 16046 8654 16098
rect 8706 16046 8718 16098
rect 7870 16034 7922 16046
rect 11454 16034 11506 16046
rect 11678 16098 11730 16110
rect 11678 16034 11730 16046
rect 13470 16098 13522 16110
rect 15374 16098 15426 16110
rect 14334 16046 14346 16098
rect 14398 16046 14410 16098
rect 10558 15986 10610 15998
rect 12542 15990 12554 16042
rect 12606 15990 12618 16042
rect 13470 16034 13522 16046
rect 15374 16034 15426 16046
rect 18062 16098 18114 16110
rect 18062 16034 18114 16046
rect 19854 16098 19906 16110
rect 19854 16034 19906 16046
rect 22878 16098 22930 16110
rect 22878 16034 22930 16046
rect 26574 16098 26626 16110
rect 26574 16034 26626 16046
rect 26798 16098 26850 16110
rect 27694 16098 27746 16110
rect 32286 16098 32338 16110
rect 27122 16046 27134 16098
rect 27186 16046 27198 16098
rect 27458 16046 27470 16098
rect 27522 16046 27534 16098
rect 28354 16046 28366 16098
rect 28418 16046 28430 16098
rect 29138 16046 29150 16098
rect 29202 16046 29214 16098
rect 26798 16034 26850 16046
rect 27694 16034 27746 16046
rect 29474 16002 29486 16054
rect 29538 16002 29550 16054
rect 30034 16031 30046 16083
rect 30098 16031 30110 16083
rect 30258 16046 30270 16098
rect 30322 16046 30334 16098
rect 31042 16046 31054 16098
rect 31106 16046 31118 16098
rect 31378 16046 31390 16098
rect 31442 16046 31454 16098
rect 32286 16034 32338 16046
rect 34078 16098 34130 16110
rect 34078 16034 34130 16046
rect 34190 16098 34242 16110
rect 34190 16034 34242 16046
rect 35646 16098 35698 16110
rect 35646 16034 35698 16046
rect 37326 16098 37378 16110
rect 37326 16034 37378 16046
rect 38446 16098 38498 16110
rect 38446 16034 38498 16046
rect 10558 15922 10610 15934
rect 14590 15986 14642 15998
rect 14590 15922 14642 15934
rect 34526 15986 34578 15998
rect 34526 15922 34578 15934
rect 38204 15986 38256 15998
rect 38938 15990 38950 16042
rect 39002 15990 39014 16042
rect 38204 15922 38256 15934
rect 39118 15986 39170 15998
rect 39118 15922 39170 15934
rect 39846 15986 39898 15998
rect 39846 15922 39898 15934
rect 11118 15874 11170 15886
rect 11118 15810 11170 15822
rect 19518 15874 19570 15886
rect 19518 15810 19570 15822
rect 28030 15874 28082 15886
rect 28030 15810 28082 15822
rect 32678 15874 32730 15886
rect 32678 15810 32730 15822
rect 35310 15874 35362 15886
rect 35310 15810 35362 15822
rect 1344 15706 44576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 44576 15706
rect 1344 15620 44576 15654
rect 7366 15538 7418 15550
rect 7366 15474 7418 15486
rect 11566 15538 11618 15550
rect 11566 15474 11618 15486
rect 24278 15538 24330 15550
rect 24278 15474 24330 15486
rect 25398 15538 25450 15550
rect 25398 15474 25450 15486
rect 43654 15538 43706 15550
rect 43654 15474 43706 15486
rect 23774 15426 23826 15438
rect 7522 15262 7534 15314
rect 7586 15262 7598 15314
rect 7858 15262 7870 15314
rect 7922 15262 7934 15314
rect 8082 15277 8094 15329
rect 8146 15277 8158 15329
rect 8642 15262 8654 15314
rect 8706 15262 8718 15314
rect 8866 15306 8878 15358
rect 8930 15306 8942 15358
rect 13694 15353 13746 15365
rect 10210 15289 10222 15341
rect 10274 15289 10286 15341
rect 12898 15262 12910 15314
rect 12962 15262 12974 15314
rect 13234 15262 13246 15314
rect 13298 15262 13310 15314
rect 13694 15289 13746 15301
rect 13918 15314 13970 15326
rect 13918 15250 13970 15262
rect 14254 15314 14306 15326
rect 14254 15250 14306 15262
rect 14814 15314 14866 15326
rect 15486 15314 15538 15326
rect 14814 15250 14866 15262
rect 14982 15258 15034 15270
rect 13582 15202 13634 15214
rect 8194 15150 8206 15202
rect 8258 15150 8270 15202
rect 8978 15150 8990 15202
rect 9042 15150 9054 15202
rect 15486 15250 15538 15262
rect 16942 15314 16994 15326
rect 16942 15250 16994 15262
rect 17484 15314 17536 15326
rect 17484 15250 17536 15262
rect 17726 15314 17778 15326
rect 18218 15318 18230 15370
rect 18282 15318 18294 15370
rect 23774 15362 23826 15374
rect 29486 15426 29538 15438
rect 29486 15362 29538 15374
rect 32006 15426 32058 15438
rect 17726 15250 17778 15262
rect 18398 15314 18450 15326
rect 18398 15250 18450 15262
rect 19182 15314 19234 15326
rect 19182 15250 19234 15262
rect 21758 15314 21810 15326
rect 21758 15250 21810 15262
rect 22542 15314 22594 15326
rect 22542 15250 22594 15262
rect 22860 15314 22912 15326
rect 22860 15250 22912 15262
rect 23102 15314 23154 15326
rect 26126 15314 26178 15326
rect 23102 15250 23154 15262
rect 23606 15258 23658 15270
rect 14982 15194 15034 15206
rect 18846 15202 18898 15214
rect 13582 15138 13634 15150
rect 18846 15138 18898 15150
rect 19574 15202 19626 15214
rect 19574 15138 19626 15150
rect 21422 15202 21474 15214
rect 26126 15250 26178 15262
rect 26798 15314 26850 15326
rect 26798 15250 26850 15262
rect 30158 15314 30210 15326
rect 30482 15318 30494 15370
rect 30546 15318 30558 15370
rect 32006 15362 32058 15374
rect 39902 15426 39954 15438
rect 39902 15362 39954 15374
rect 41470 15426 41522 15438
rect 41470 15362 41522 15374
rect 31054 15314 31106 15326
rect 30706 15262 30718 15314
rect 30770 15262 30782 15314
rect 30158 15250 30210 15262
rect 31054 15250 31106 15262
rect 32958 15314 33010 15326
rect 32958 15250 33010 15262
rect 34862 15314 34914 15326
rect 34862 15250 34914 15262
rect 35198 15314 35250 15326
rect 35198 15250 35250 15262
rect 36766 15314 36818 15326
rect 36766 15250 36818 15262
rect 37102 15314 37154 15326
rect 37102 15250 37154 15262
rect 37214 15314 37266 15326
rect 37214 15250 37266 15262
rect 41638 15314 41690 15326
rect 41638 15250 41690 15262
rect 42142 15314 42194 15326
rect 42142 15250 42194 15262
rect 42702 15314 42754 15326
rect 42702 15250 42754 15262
rect 23606 15194 23658 15206
rect 26462 15202 26514 15214
rect 31390 15202 31442 15214
rect 21422 15138 21474 15150
rect 27570 15150 27582 15202
rect 27634 15150 27646 15202
rect 30594 15150 30606 15202
rect 30658 15150 30670 15202
rect 26462 15138 26514 15150
rect 31390 15138 31442 15150
rect 33294 15202 33346 15214
rect 33294 15138 33346 15150
rect 36374 15202 36426 15214
rect 43038 15202 43090 15214
rect 37986 15150 37998 15202
rect 38050 15150 38062 15202
rect 36374 15138 36426 15150
rect 43038 15138 43090 15150
rect 12742 15090 12794 15102
rect 12742 15026 12794 15038
rect 15728 15090 15780 15102
rect 15728 15026 15780 15038
rect 16606 15090 16658 15102
rect 16606 15026 16658 15038
rect 22206 15090 22258 15102
rect 22206 15026 22258 15038
rect 34526 15090 34578 15102
rect 34526 15026 34578 15038
rect 35534 15090 35586 15102
rect 35534 15026 35586 15038
rect 42384 15090 42436 15102
rect 42384 15026 42436 15038
rect 1344 14922 44576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 44576 14922
rect 1344 14836 44576 14870
rect 11454 14754 11506 14766
rect 11454 14690 11506 14702
rect 14590 14754 14642 14766
rect 14590 14690 14642 14702
rect 19276 14754 19328 14766
rect 19276 14690 19328 14702
rect 28384 14754 28436 14766
rect 28384 14690 28436 14702
rect 34956 14754 35008 14766
rect 34956 14690 35008 14702
rect 38782 14754 38834 14766
rect 38782 14690 38834 14702
rect 31334 14642 31386 14654
rect 8754 14590 8766 14642
rect 8818 14590 8830 14642
rect 16818 14590 16830 14642
rect 16882 14590 16894 14642
rect 18722 14590 18734 14642
rect 18786 14590 18798 14642
rect 27638 14586 27690 14598
rect 8990 14530 9042 14542
rect 7746 14478 7758 14530
rect 7810 14478 7822 14530
rect 8418 14478 8430 14530
rect 8482 14478 8494 14530
rect 8642 14434 8654 14486
rect 8706 14434 8718 14486
rect 13470 14530 13522 14542
rect 8990 14466 9042 14478
rect 10098 14450 10110 14502
rect 10162 14450 10174 14502
rect 13470 14466 13522 14478
rect 15598 14530 15650 14542
rect 14334 14422 14346 14474
rect 14398 14422 14410 14474
rect 15598 14466 15650 14478
rect 15934 14530 15986 14542
rect 15934 14466 15986 14478
rect 16046 14530 16098 14542
rect 16046 14466 16098 14478
rect 19518 14530 19570 14542
rect 24446 14530 24498 14542
rect 19518 14466 19570 14478
rect 20010 14422 20022 14474
rect 20074 14422 20086 14474
rect 21410 14450 21422 14502
rect 21474 14450 21486 14502
rect 24446 14466 24498 14478
rect 25118 14530 25170 14542
rect 24204 14418 24256 14430
rect 24938 14422 24950 14474
rect 25002 14422 25014 14474
rect 25118 14466 25170 14478
rect 27246 14530 27298 14542
rect 27246 14466 27298 14478
rect 27470 14530 27522 14542
rect 41570 14590 41582 14642
rect 41634 14590 41646 14642
rect 31334 14578 31386 14590
rect 27638 14522 27690 14534
rect 28142 14530 28194 14542
rect 27470 14466 27522 14478
rect 28142 14466 28194 14478
rect 29486 14530 29538 14542
rect 29486 14466 29538 14478
rect 30942 14530 30994 14542
rect 7926 14306 7978 14318
rect 19842 14310 19854 14362
rect 19906 14310 19918 14362
rect 24204 14354 24256 14366
rect 29244 14418 29296 14430
rect 29978 14422 29990 14474
rect 30042 14422 30054 14474
rect 30942 14466 30994 14478
rect 34190 14530 34242 14542
rect 34190 14466 34242 14478
rect 35198 14530 35250 14542
rect 35198 14466 35250 14478
rect 36374 14530 36426 14542
rect 29244 14354 29296 14366
rect 30606 14418 30658 14430
rect 35690 14422 35702 14474
rect 35754 14422 35766 14474
rect 36374 14466 36426 14478
rect 37662 14530 37714 14542
rect 7926 14242 7978 14254
rect 22654 14306 22706 14318
rect 22654 14242 22706 14254
rect 26518 14306 26570 14318
rect 26518 14242 26570 14254
rect 26910 14306 26962 14318
rect 29810 14310 29822 14362
rect 29874 14310 29886 14362
rect 30606 14354 30658 14366
rect 35870 14418 35922 14430
rect 35870 14354 35922 14366
rect 36990 14418 37042 14430
rect 37146 14422 37158 14474
rect 37210 14422 37222 14474
rect 37662 14466 37714 14478
rect 38446 14530 38498 14542
rect 38446 14466 38498 14478
rect 40798 14530 40850 14542
rect 40798 14466 40850 14478
rect 36990 14354 37042 14366
rect 37904 14418 37956 14430
rect 37904 14354 37956 14366
rect 43486 14418 43538 14430
rect 43486 14354 43538 14366
rect 26910 14242 26962 14254
rect 33854 14306 33906 14318
rect 33854 14242 33906 14254
rect 44102 14306 44154 14318
rect 44102 14242 44154 14254
rect 1344 14138 44576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 44576 14138
rect 1344 14052 44576 14086
rect 41190 13970 41242 13982
rect 9662 13858 9714 13870
rect 9662 13794 9714 13806
rect 14254 13858 14306 13870
rect 16482 13862 16494 13914
rect 16546 13862 16558 13914
rect 41190 13906 41242 13918
rect 14254 13794 14306 13806
rect 19966 13858 20018 13870
rect 19966 13794 20018 13806
rect 21310 13858 21362 13870
rect 21310 13794 21362 13806
rect 30382 13858 30434 13870
rect 30382 13794 30434 13806
rect 41470 13858 41522 13870
rect 41470 13794 41522 13806
rect 42384 13858 42436 13870
rect 43474 13862 43486 13914
rect 43538 13862 43550 13914
rect 42384 13794 42436 13806
rect 7522 13694 7534 13746
rect 7586 13694 7598 13746
rect 7746 13694 7758 13746
rect 7810 13694 7822 13746
rect 8082 13709 8094 13761
rect 8146 13709 8158 13761
rect 8530 13694 8542 13746
rect 8594 13694 8606 13746
rect 8866 13738 8878 13790
rect 8930 13738 8942 13790
rect 12350 13746 12402 13758
rect 11554 13694 11566 13746
rect 11618 13694 11630 13746
rect 12350 13682 12402 13694
rect 13134 13746 13186 13758
rect 15598 13746 15650 13758
rect 13998 13694 14010 13746
rect 14062 13694 14074 13746
rect 13134 13682 13186 13694
rect 15598 13682 15650 13694
rect 15916 13746 15968 13758
rect 15916 13682 15968 13694
rect 16158 13746 16210 13758
rect 17278 13746 17330 13758
rect 23998 13746 24050 13758
rect 16158 13682 16210 13694
rect 16662 13690 16714 13702
rect 18050 13694 18062 13746
rect 18114 13694 18126 13746
rect 17278 13682 17330 13694
rect 23998 13682 24050 13694
rect 24110 13746 24162 13758
rect 24110 13682 24162 13694
rect 27694 13746 27746 13758
rect 27694 13682 27746 13694
rect 32062 13746 32114 13758
rect 32062 13682 32114 13694
rect 33070 13746 33122 13758
rect 33070 13682 33122 13694
rect 36094 13746 36146 13758
rect 39118 13746 39170 13758
rect 36866 13694 36878 13746
rect 36930 13694 36942 13746
rect 36094 13682 36146 13694
rect 39118 13682 39170 13694
rect 40462 13746 40514 13758
rect 42142 13746 42194 13758
rect 40462 13682 40514 13694
rect 41638 13690 41690 13702
rect 8194 13582 8206 13634
rect 8258 13582 8270 13634
rect 8978 13582 8990 13634
rect 9042 13582 9054 13634
rect 16662 13626 16714 13638
rect 24446 13634 24498 13646
rect 42142 13682 42194 13694
rect 42908 13746 42960 13758
rect 42908 13682 42960 13694
rect 43150 13746 43202 13758
rect 43150 13682 43202 13694
rect 43654 13690 43706 13702
rect 23202 13582 23214 13634
rect 23266 13582 23278 13634
rect 28466 13582 28478 13634
rect 28530 13582 28542 13634
rect 33842 13582 33854 13634
rect 33906 13582 33918 13634
rect 35746 13582 35758 13634
rect 35810 13582 35822 13634
rect 38770 13582 38782 13634
rect 38834 13582 38846 13634
rect 41638 13626 41690 13638
rect 43654 13626 43706 13638
rect 24446 13570 24498 13582
rect 7366 13522 7418 13534
rect 7366 13458 7418 13470
rect 15262 13522 15314 13534
rect 15262 13458 15314 13470
rect 31726 13522 31778 13534
rect 31726 13458 31778 13470
rect 39454 13522 39506 13534
rect 39454 13458 39506 13470
rect 40126 13522 40178 13534
rect 40126 13458 40178 13470
rect 1344 13354 44576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 44576 13354
rect 1344 13268 44576 13302
rect 29374 13186 29426 13198
rect 29374 13122 29426 13134
rect 30606 13186 30658 13198
rect 30606 13122 30658 13134
rect 32044 13186 32096 13198
rect 32044 13122 32096 13134
rect 18230 13074 18282 13086
rect 33462 13074 33514 13086
rect 9762 13022 9774 13074
rect 9826 13022 9838 13074
rect 11666 13022 11678 13074
rect 11730 13022 11742 13074
rect 14466 13022 14478 13074
rect 14530 13022 14542 13074
rect 16370 13022 16382 13074
rect 16434 13022 16446 13074
rect 21970 13022 21982 13074
rect 22034 13022 22046 13074
rect 38994 13022 39006 13074
rect 39058 13022 39070 13074
rect 41346 13022 41358 13074
rect 41410 13022 41422 13074
rect 18230 13010 18282 13022
rect 33462 13010 33514 13022
rect 8990 12962 9042 12974
rect 8990 12898 9042 12910
rect 17166 12962 17218 12974
rect 17166 12898 17218 12910
rect 17278 12962 17330 12974
rect 17278 12898 17330 12910
rect 20302 12962 20354 12974
rect 20302 12898 20354 12910
rect 21198 12962 21250 12974
rect 21198 12898 21250 12910
rect 25678 12962 25730 12974
rect 25678 12898 25730 12910
rect 27358 12962 27410 12974
rect 23886 12850 23938 12862
rect 23886 12786 23938 12798
rect 26686 12850 26738 12862
rect 26842 12854 26854 12906
rect 26906 12854 26918 12906
rect 27358 12898 27410 12910
rect 29038 12962 29090 12974
rect 29038 12898 29090 12910
rect 30270 12962 30322 12974
rect 30270 12898 30322 12910
rect 31502 12962 31554 12974
rect 31502 12898 31554 12910
rect 32286 12962 32338 12974
rect 32286 12898 32338 12910
rect 32958 12962 33010 12974
rect 26686 12786 26738 12798
rect 27600 12850 27652 12862
rect 32778 12854 32790 12906
rect 32842 12854 32854 12906
rect 32958 12898 33010 12910
rect 34190 12962 34242 12974
rect 34190 12898 34242 12910
rect 34358 12962 34410 12974
rect 34358 12898 34410 12910
rect 34862 12962 34914 12974
rect 39790 12962 39842 12974
rect 35746 12910 35758 12962
rect 35810 12910 35822 12962
rect 34862 12898 34914 12910
rect 39790 12898 39842 12910
rect 40574 12962 40626 12974
rect 40574 12898 40626 12910
rect 43598 12962 43650 12974
rect 43598 12898 43650 12910
rect 27600 12786 27652 12798
rect 35104 12850 35156 12862
rect 35104 12786 35156 12798
rect 37102 12850 37154 12862
rect 37102 12786 37154 12798
rect 43262 12850 43314 12862
rect 43262 12786 43314 12798
rect 17614 12738 17666 12750
rect 17614 12674 17666 12686
rect 19966 12738 20018 12750
rect 19966 12674 20018 12686
rect 25342 12738 25394 12750
rect 25342 12674 25394 12686
rect 26406 12738 26458 12750
rect 26406 12674 26458 12686
rect 31166 12738 31218 12750
rect 31166 12674 31218 12686
rect 35590 12738 35642 12750
rect 35590 12674 35642 12686
rect 36150 12738 36202 12750
rect 36150 12674 36202 12686
rect 43934 12738 43986 12750
rect 43934 12674 43986 12686
rect 1344 12570 44576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 44576 12570
rect 1344 12484 44576 12518
rect 28870 12402 28922 12414
rect 28870 12338 28922 12350
rect 36430 12402 36482 12414
rect 36430 12338 36482 12350
rect 12126 12290 12178 12302
rect 12126 12226 12178 12238
rect 13694 12290 13746 12302
rect 9438 12178 9490 12190
rect 12574 12178 12626 12190
rect 13438 12182 13450 12234
rect 13502 12182 13514 12234
rect 13694 12226 13746 12238
rect 14254 12290 14306 12302
rect 14254 12226 14306 12238
rect 25230 12290 25282 12302
rect 25230 12226 25282 12238
rect 26574 12290 26626 12302
rect 26574 12226 26626 12238
rect 43598 12290 43650 12302
rect 43598 12226 43650 12238
rect 16942 12178 16994 12190
rect 10210 12126 10222 12178
rect 10274 12126 10286 12178
rect 16146 12126 16158 12178
rect 16210 12126 16222 12178
rect 18386 12126 18398 12178
rect 18450 12126 18462 12178
rect 18722 12141 18734 12193
rect 18786 12141 18798 12193
rect 19394 12153 19406 12205
rect 19458 12153 19470 12205
rect 21870 12178 21922 12190
rect 21410 12126 21422 12178
rect 21474 12126 21486 12178
rect 25902 12178 25954 12190
rect 9438 12114 9490 12126
rect 12574 12114 12626 12126
rect 16942 12114 16994 12126
rect 21870 12114 21922 12126
rect 25398 12122 25450 12134
rect 27246 12178 27298 12190
rect 25902 12114 25954 12126
rect 26742 12122 26794 12134
rect 18834 12014 18846 12066
rect 18898 12014 18910 12066
rect 22642 12014 22654 12066
rect 22706 12014 22718 12066
rect 24546 12014 24558 12066
rect 24610 12014 24622 12066
rect 25398 12058 25450 12070
rect 27246 12114 27298 12126
rect 27806 12178 27858 12190
rect 27806 12114 27858 12126
rect 29710 12178 29762 12190
rect 30482 12126 30494 12178
rect 30546 12126 30558 12178
rect 33618 12153 33630 12205
rect 33682 12153 33694 12205
rect 35086 12178 35138 12190
rect 29710 12114 29762 12126
rect 35086 12114 35138 12126
rect 36094 12178 36146 12190
rect 37314 12153 37326 12205
rect 37378 12153 37390 12205
rect 40910 12178 40962 12190
rect 36094 12114 36146 12126
rect 41682 12126 41694 12178
rect 41746 12126 41758 12178
rect 40910 12114 40962 12126
rect 26742 12058 26794 12070
rect 44214 12066 44266 12078
rect 32386 12014 32398 12066
rect 32450 12014 32462 12066
rect 44214 12002 44266 12014
rect 26144 11954 26196 11966
rect 26144 11890 26196 11902
rect 27488 11954 27540 11966
rect 27488 11890 27540 11902
rect 28142 11954 28194 11966
rect 28142 11890 28194 11902
rect 39006 11954 39058 11966
rect 39006 11890 39058 11902
rect 1344 11786 44576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 44576 11786
rect 1344 11700 44576 11734
rect 11342 11618 11394 11630
rect 11342 11554 11394 11566
rect 22318 11618 22370 11630
rect 22318 11554 22370 11566
rect 43934 11618 43986 11630
rect 43934 11554 43986 11566
rect 24670 11506 24722 11518
rect 39902 11506 39954 11518
rect 18722 11454 18734 11506
rect 18786 11454 18798 11506
rect 20626 11454 20638 11506
rect 20690 11454 20702 11506
rect 26002 11454 26014 11506
rect 26066 11454 26078 11506
rect 27906 11454 27918 11506
rect 27970 11454 27982 11506
rect 34514 11454 34526 11506
rect 34578 11454 34590 11506
rect 35858 11454 35870 11506
rect 35922 11454 35934 11506
rect 24670 11442 24722 11454
rect 39902 11442 39954 11454
rect 17950 11394 18002 11406
rect 12002 11314 12014 11366
rect 12066 11314 12078 11366
rect 24334 11394 24386 11406
rect 28702 11394 28754 11406
rect 17950 11330 18002 11342
rect 21634 11314 21646 11366
rect 21698 11314 21710 11366
rect 24882 11342 24894 11394
rect 24946 11342 24958 11394
rect 24334 11330 24386 11342
rect 24546 11286 24558 11338
rect 24610 11286 24622 11338
rect 28702 11330 28754 11342
rect 29038 11394 29090 11406
rect 41022 11394 41074 11406
rect 42590 11394 42642 11406
rect 43542 11394 43594 11406
rect 29810 11342 29822 11394
rect 29874 11342 29886 11394
rect 29038 11330 29090 11342
rect 32274 11298 32286 11350
rect 32338 11298 32350 11350
rect 32498 11342 32510 11394
rect 32562 11342 32574 11394
rect 35522 11314 35534 11366
rect 35586 11314 35598 11366
rect 35970 11327 35982 11379
rect 36034 11327 36046 11379
rect 36194 11342 36206 11394
rect 36258 11342 36270 11394
rect 37202 11342 37214 11394
rect 37266 11342 37278 11394
rect 39218 11314 39230 11366
rect 39282 11314 39294 11366
rect 40133 11342 40145 11394
rect 40197 11342 40209 11394
rect 41701 11342 41713 11394
rect 41765 11342 41777 11394
rect 42802 11342 42814 11394
rect 42866 11342 42878 11394
rect 41022 11330 41074 11342
rect 42590 11330 42642 11342
rect 43542 11330 43594 11342
rect 44270 11394 44322 11406
rect 44270 11330 44322 11342
rect 31726 11282 31778 11294
rect 31726 11218 31778 11230
rect 41470 11282 41522 11294
rect 17110 11170 17162 11182
rect 32498 11174 32510 11226
rect 32562 11174 32574 11226
rect 41470 11218 41522 11230
rect 17110 11106 17162 11118
rect 42982 11170 43034 11182
rect 42982 11106 43034 11118
rect 1344 11002 44576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 44576 11002
rect 1344 10916 44576 10950
rect 24446 10834 24498 10846
rect 24446 10770 24498 10782
rect 23886 10722 23938 10734
rect 14030 10610 14082 10622
rect 14030 10546 14082 10558
rect 16718 10610 16770 10622
rect 17490 10573 17502 10625
rect 17554 10573 17566 10625
rect 18958 10610 19010 10622
rect 17826 10558 17838 10610
rect 17890 10558 17902 10610
rect 16718 10546 16770 10558
rect 18958 10546 19010 10558
rect 21982 10610 22034 10622
rect 22766 10610 22818 10622
rect 23630 10614 23642 10666
rect 23694 10614 23706 10666
rect 23886 10658 23938 10670
rect 25342 10722 25394 10734
rect 25342 10658 25394 10670
rect 22418 10558 22430 10610
rect 22482 10558 22494 10610
rect 21982 10546 22034 10558
rect 22766 10546 22818 10558
rect 24782 10610 24834 10622
rect 24782 10546 24834 10558
rect 28030 10610 28082 10622
rect 28030 10546 28082 10558
rect 28142 10610 28194 10622
rect 31826 10585 31838 10637
rect 31890 10585 31902 10637
rect 33070 10610 33122 10622
rect 33934 10614 33946 10666
rect 33998 10614 34010 10666
rect 32610 10558 32622 10610
rect 32674 10558 32686 10610
rect 28142 10546 28194 10558
rect 33070 10546 33122 10558
rect 34190 10610 34242 10622
rect 34906 10614 34918 10666
rect 34970 10614 34982 10666
rect 39342 10649 39394 10661
rect 35422 10610 35474 10622
rect 34626 10558 34638 10610
rect 34690 10558 34702 10610
rect 34190 10546 34242 10558
rect 35422 10546 35474 10558
rect 38782 10610 38834 10622
rect 38782 10546 38834 10558
rect 39118 10610 39170 10622
rect 41246 10610 41298 10622
rect 41477 10614 41489 10666
rect 41541 10614 41553 10666
rect 39342 10585 39394 10597
rect 39666 10558 39678 10610
rect 39730 10558 39742 10610
rect 40002 10558 40014 10610
rect 40066 10558 40078 10610
rect 39118 10546 39170 10558
rect 41246 10546 41298 10558
rect 42366 10610 42418 10622
rect 43045 10614 43057 10666
rect 43109 10614 43121 10666
rect 42366 10546 42418 10558
rect 43934 10610 43986 10622
rect 43934 10546 43986 10558
rect 28478 10498 28530 10510
rect 14802 10446 14814 10498
rect 14866 10446 14878 10498
rect 17378 10446 17390 10498
rect 17442 10446 17454 10498
rect 19282 10446 19294 10498
rect 19346 10446 19358 10498
rect 21186 10446 21198 10498
rect 21250 10446 21262 10498
rect 22262 10442 22314 10454
rect 27234 10446 27246 10498
rect 27298 10446 27310 10498
rect 35074 10446 35086 10498
rect 35138 10446 35150 10498
rect 36194 10446 36206 10498
rect 36258 10446 36270 10498
rect 38098 10446 38110 10498
rect 38162 10446 38174 10498
rect 39554 10446 39566 10498
rect 39618 10446 39630 10498
rect 18622 10386 18674 10398
rect 28478 10434 28530 10446
rect 22262 10378 22314 10390
rect 30942 10386 30994 10398
rect 18622 10322 18674 10334
rect 30942 10322 30994 10334
rect 32454 10386 32506 10398
rect 32454 10322 32506 10334
rect 40182 10386 40234 10398
rect 40182 10322 40234 10334
rect 42814 10386 42866 10398
rect 42814 10322 42866 10334
rect 1344 10218 44576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 44576 10218
rect 1344 10132 44576 10166
rect 22318 10050 22370 10062
rect 22318 9986 22370 9998
rect 30270 10050 30322 10062
rect 36318 10050 36370 10062
rect 30270 9986 30322 9998
rect 31446 9994 31498 10006
rect 36318 9986 36370 9998
rect 16930 9886 16942 9938
rect 16994 9886 17006 9938
rect 19730 9886 19742 9938
rect 19794 9886 19806 9938
rect 31446 9930 31498 9942
rect 32498 9886 32510 9938
rect 32562 9886 32574 9938
rect 34402 9886 34414 9938
rect 34466 9886 34478 9938
rect 24110 9826 24162 9838
rect 26238 9826 26290 9838
rect 30606 9826 30658 9838
rect 17938 9746 17950 9798
rect 18002 9746 18014 9798
rect 20402 9746 20414 9798
rect 20466 9746 20478 9798
rect 21298 9746 21310 9798
rect 21362 9746 21374 9798
rect 24974 9774 24986 9826
rect 25038 9774 25050 9826
rect 27102 9774 27114 9826
rect 27166 9774 27178 9826
rect 31726 9826 31778 9838
rect 24110 9762 24162 9774
rect 26238 9762 26290 9774
rect 30606 9762 30658 9774
rect 31614 9770 31666 9782
rect 25230 9714 25282 9726
rect 25230 9650 25282 9662
rect 27358 9714 27410 9726
rect 31726 9762 31778 9774
rect 35198 9826 35250 9838
rect 35198 9762 35250 9774
rect 36878 9826 36930 9838
rect 39566 9826 39618 9838
rect 37650 9774 37662 9826
rect 37714 9774 37726 9826
rect 36062 9718 36074 9770
rect 36126 9718 36138 9770
rect 36878 9762 36930 9774
rect 39566 9762 39618 9774
rect 39902 9826 39954 9838
rect 44270 9826 44322 9838
rect 40674 9774 40686 9826
rect 40738 9774 40750 9826
rect 42914 9774 42926 9826
rect 42978 9774 42990 9826
rect 39902 9762 39954 9774
rect 44270 9762 44322 9774
rect 31614 9706 31666 9718
rect 42590 9714 42642 9726
rect 27358 9650 27410 9662
rect 42590 9650 42642 9662
rect 43094 9602 43146 9614
rect 43094 9538 43146 9550
rect 43934 9602 43986 9614
rect 43934 9538 43986 9550
rect 1344 9434 44576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 44576 9434
rect 1344 9348 44576 9382
rect 16774 9266 16826 9278
rect 16774 9202 16826 9214
rect 23326 9266 23378 9278
rect 37998 9266 38050 9278
rect 23326 9202 23378 9214
rect 25566 9210 25618 9222
rect 37998 9202 38050 9214
rect 39554 9158 39566 9210
rect 39618 9158 39630 9210
rect 25566 9146 25618 9158
rect 18342 9071 18394 9083
rect 16482 8990 16494 9042
rect 16546 8990 16558 9042
rect 16930 8990 16942 9042
rect 16994 8990 17006 9042
rect 17938 8990 17950 9042
rect 18002 8990 18014 9042
rect 18846 9042 18898 9054
rect 18342 9007 18394 9019
rect 18610 8990 18622 9042
rect 18674 8990 18686 9042
rect 21970 9017 21982 9069
rect 22034 9017 22046 9069
rect 25330 8990 25342 9042
rect 25394 8990 25406 9042
rect 25554 9017 25566 9069
rect 25618 9017 25630 9069
rect 25902 9042 25954 9054
rect 18846 8978 18898 8990
rect 25902 8978 25954 8990
rect 29150 9042 29202 9054
rect 29150 8978 29202 8990
rect 29486 9042 29538 9054
rect 29486 8978 29538 8990
rect 31950 9042 32002 9054
rect 31950 8978 32002 8990
rect 33518 9042 33570 9054
rect 34290 8990 34302 9042
rect 34354 8990 34366 9042
rect 36642 9017 36654 9069
rect 36706 9017 36718 9069
rect 39722 9046 39734 9098
rect 39786 9046 39798 9098
rect 43822 9062 43874 9074
rect 40126 9042 40178 9054
rect 39442 8990 39454 9042
rect 39506 8990 39518 9042
rect 33518 8978 33570 8990
rect 40126 8978 40178 8990
rect 43710 9042 43762 9054
rect 43822 8998 43874 9010
rect 43710 8978 43762 8990
rect 16326 8874 16378 8886
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 19618 8878 19630 8930
rect 19682 8878 19694 8930
rect 21522 8878 21534 8930
rect 21586 8878 21598 8930
rect 36194 8878 36206 8930
rect 36258 8878 36270 8930
rect 41010 8878 41022 8930
rect 41074 8878 41086 8930
rect 42914 8878 42926 8930
rect 42978 8878 42990 8930
rect 16326 8810 16378 8822
rect 17782 8818 17834 8830
rect 17782 8754 17834 8766
rect 28814 8818 28866 8830
rect 28814 8754 28866 8766
rect 29822 8818 29874 8830
rect 29822 8754 29874 8766
rect 32286 8818 32338 8830
rect 32286 8754 32338 8766
rect 43990 8818 44042 8830
rect 43990 8754 44042 8766
rect 1344 8650 44576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 44576 8650
rect 1344 8564 44576 8598
rect 25230 8370 25282 8382
rect 34078 8370 34130 8382
rect 17266 8318 17278 8370
rect 17330 8318 17342 8370
rect 20066 8318 20078 8370
rect 20130 8318 20142 8370
rect 31154 8318 31166 8370
rect 31218 8318 31230 8370
rect 25230 8306 25282 8318
rect 34078 8306 34130 8318
rect 36374 8370 36426 8382
rect 36374 8306 36426 8318
rect 16494 8258 16546 8270
rect 20302 8258 20354 8270
rect 19730 8206 19742 8258
rect 19794 8206 19806 8258
rect 19910 8228 19962 8240
rect 16494 8194 16546 8206
rect 24110 8258 24162 8270
rect 26014 8258 26066 8270
rect 20302 8194 20354 8206
rect 23762 8178 23774 8230
rect 23826 8178 23838 8230
rect 24974 8206 24986 8258
rect 25038 8206 25050 8258
rect 24110 8194 24162 8206
rect 26014 8194 26066 8206
rect 26686 8258 26738 8270
rect 19910 8164 19962 8176
rect 19182 8146 19234 8158
rect 19182 8082 19234 8094
rect 25772 8146 25824 8158
rect 26506 8150 26518 8202
rect 26570 8150 26582 8202
rect 26686 8194 26738 8206
rect 29262 8258 29314 8270
rect 29262 8194 29314 8206
rect 31950 8258 32002 8270
rect 34638 8258 34690 8270
rect 43934 8258 43986 8270
rect 31950 8194 32002 8206
rect 34414 8202 34466 8214
rect 35502 8206 35514 8258
rect 35566 8206 35578 8258
rect 37202 8206 37214 8258
rect 37266 8206 37278 8258
rect 34638 8194 34690 8206
rect 37538 8178 37550 8230
rect 37602 8178 37614 8230
rect 39778 8206 39790 8258
rect 39842 8206 39854 8258
rect 40338 8178 40350 8230
rect 40402 8178 40414 8230
rect 43934 8194 43986 8206
rect 34414 8138 34466 8150
rect 35758 8146 35810 8158
rect 25772 8082 25824 8094
rect 35758 8082 35810 8094
rect 20638 8034 20690 8046
rect 20638 7970 20690 7982
rect 22094 8034 22146 8046
rect 22094 7970 22146 7982
rect 27190 8034 27242 8046
rect 27190 7970 27242 7982
rect 27638 8034 27690 8046
rect 27638 7970 27690 7982
rect 37046 8034 37098 8046
rect 37046 7970 37098 7982
rect 41694 8034 41746 8046
rect 41694 7970 41746 7982
rect 1344 7866 44576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 44576 7866
rect 1344 7780 44576 7814
rect 16774 7698 16826 7710
rect 16774 7634 16826 7646
rect 28646 7698 28698 7710
rect 18722 7590 18734 7642
rect 18786 7590 18798 7642
rect 28646 7634 28698 7646
rect 23438 7586 23490 7598
rect 16930 7422 16942 7474
rect 16994 7422 17006 7474
rect 17490 7466 17502 7518
rect 17554 7466 17566 7518
rect 17826 7422 17838 7474
rect 17890 7422 17902 7474
rect 18498 7437 18510 7489
rect 18562 7437 18574 7489
rect 19070 7474 19122 7486
rect 18834 7422 18846 7474
rect 18898 7422 18910 7474
rect 19070 7410 19122 7422
rect 22318 7474 22370 7486
rect 23182 7478 23194 7530
rect 23246 7478 23258 7530
rect 23438 7522 23490 7534
rect 25566 7586 25618 7598
rect 25566 7522 25618 7534
rect 29132 7586 29184 7598
rect 29132 7522 29184 7534
rect 30046 7586 30098 7598
rect 26238 7474 26290 7486
rect 22318 7410 22370 7422
rect 25734 7418 25786 7430
rect 26898 7422 26910 7474
rect 26962 7422 26974 7474
rect 27234 7449 27246 7501
rect 27298 7449 27310 7501
rect 27582 7474 27634 7486
rect 26238 7410 26290 7422
rect 27582 7410 27634 7422
rect 27918 7474 27970 7486
rect 27918 7410 27970 7422
rect 29374 7474 29426 7486
rect 29866 7478 29878 7530
rect 29930 7478 29942 7530
rect 30046 7522 30098 7534
rect 29374 7410 29426 7422
rect 30270 7474 30322 7486
rect 30270 7410 30322 7422
rect 35758 7474 35810 7486
rect 36082 7466 36094 7518
rect 36146 7466 36158 7518
rect 36990 7474 37042 7486
rect 36418 7422 36430 7474
rect 36482 7422 36494 7474
rect 35758 7410 35810 7422
rect 36990 7410 37042 7422
rect 37326 7474 37378 7486
rect 37706 7478 37718 7530
rect 37770 7478 37782 7530
rect 38677 7478 38689 7530
rect 38741 7478 38753 7530
rect 39566 7474 39618 7486
rect 37986 7422 37998 7474
rect 38050 7422 38062 7474
rect 40002 7466 40014 7518
rect 40066 7466 40078 7518
rect 40338 7422 40350 7474
rect 40402 7422 40414 7474
rect 40898 7449 40910 7501
rect 40962 7449 40974 7501
rect 42254 7474 42306 7486
rect 43810 7437 43822 7489
rect 43874 7437 43886 7489
rect 44034 7422 44046 7474
rect 44098 7422 44110 7474
rect 37326 7410 37378 7422
rect 39566 7410 39618 7422
rect 42254 7410 42306 7422
rect 17378 7310 17390 7362
rect 17442 7310 17454 7362
rect 19842 7310 19854 7362
rect 19906 7310 19918 7362
rect 21746 7310 21758 7362
rect 21810 7310 21822 7362
rect 25734 7354 25786 7366
rect 37662 7362 37714 7374
rect 27010 7310 27022 7362
rect 27074 7310 27086 7362
rect 35970 7310 35982 7362
rect 36034 7310 36046 7362
rect 37662 7298 37714 7310
rect 38446 7362 38498 7374
rect 39890 7310 39902 7362
rect 39954 7310 39966 7362
rect 43698 7310 43710 7362
rect 43762 7310 43774 7362
rect 38446 7298 38498 7310
rect 26480 7250 26532 7262
rect 26480 7186 26532 7198
rect 30606 7250 30658 7262
rect 30606 7186 30658 7198
rect 35422 7250 35474 7262
rect 35422 7186 35474 7198
rect 1344 7082 44576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 44576 7082
rect 1344 6996 44576 7030
rect 22318 6914 22370 6926
rect 22318 6850 22370 6862
rect 28366 6914 28418 6926
rect 28366 6850 28418 6862
rect 24210 6750 24222 6802
rect 24274 6750 24286 6802
rect 37090 6750 37102 6802
rect 37154 6750 37166 6802
rect 43250 6750 43262 6802
rect 43314 6750 43326 6802
rect 15822 6690 15874 6702
rect 19518 6690 19570 6702
rect 16594 6638 16606 6690
rect 16658 6638 16670 6690
rect 18946 6638 18958 6690
rect 19010 6638 19022 6690
rect 15822 6626 15874 6638
rect 19518 6626 19570 6638
rect 20638 6690 20690 6702
rect 24782 6690 24834 6702
rect 18510 6578 18562 6590
rect 20382 6582 20394 6634
rect 20446 6582 20458 6634
rect 20638 6626 20690 6638
rect 21634 6610 21646 6662
rect 21698 6610 21710 6662
rect 24098 6638 24110 6690
rect 24162 6638 24174 6690
rect 24434 6611 24446 6663
rect 24498 6611 24510 6663
rect 24782 6626 24834 6638
rect 25118 6690 25170 6702
rect 25118 6626 25170 6638
rect 26910 6690 26962 6702
rect 18510 6514 18562 6526
rect 25790 6578 25842 6590
rect 26021 6582 26033 6634
rect 26085 6582 26097 6634
rect 26910 6626 26962 6638
rect 27246 6690 27298 6702
rect 29486 6690 29538 6702
rect 28110 6638 28122 6690
rect 28174 6638 28186 6690
rect 27246 6626 27298 6638
rect 29486 6626 29538 6638
rect 29654 6690 29706 6702
rect 29654 6626 29706 6638
rect 30158 6690 30210 6702
rect 30158 6626 30210 6638
rect 30400 6690 30452 6702
rect 30400 6626 30452 6638
rect 30718 6690 30770 6702
rect 30718 6626 30770 6638
rect 34078 6690 34130 6702
rect 34078 6626 34130 6638
rect 35758 6690 35810 6702
rect 37662 6690 37714 6702
rect 36978 6638 36990 6690
rect 37042 6638 37054 6690
rect 44046 6690 44098 6702
rect 25790 6514 25842 6526
rect 33836 6578 33888 6590
rect 34570 6582 34582 6634
rect 34634 6582 34646 6634
rect 33836 6514 33888 6526
rect 34750 6578 34802 6590
rect 34750 6514 34802 6526
rect 35086 6578 35138 6590
rect 35242 6582 35254 6634
rect 35306 6582 35318 6634
rect 35758 6626 35810 6638
rect 35086 6514 35138 6526
rect 36000 6578 36052 6590
rect 37314 6582 37326 6634
rect 37378 6582 37390 6634
rect 37662 6626 37714 6638
rect 38770 6610 38782 6662
rect 38834 6610 38846 6662
rect 44046 6626 44098 6638
rect 36000 6514 36052 6526
rect 41358 6578 41410 6590
rect 41358 6514 41410 6526
rect 19126 6466 19178 6478
rect 19126 6402 19178 6414
rect 31054 6466 31106 6478
rect 31054 6402 31106 6414
rect 31670 6466 31722 6478
rect 31670 6402 31722 6414
rect 40126 6466 40178 6478
rect 40126 6402 40178 6414
rect 1344 6298 44576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 44576 6298
rect 1344 6212 44576 6246
rect 16326 6130 16378 6142
rect 16326 6066 16378 6078
rect 24558 6018 24610 6030
rect 24558 5954 24610 5966
rect 26462 6018 26514 6030
rect 26462 5954 26514 5966
rect 28814 6018 28866 6030
rect 28814 5954 28866 5966
rect 29374 6018 29426 6030
rect 29374 5954 29426 5966
rect 33742 6018 33794 6030
rect 33742 5954 33794 5966
rect 35422 6018 35474 6030
rect 37314 6022 37326 6074
rect 37378 6022 37390 6074
rect 35422 5954 35474 5966
rect 16482 5854 16494 5906
rect 16546 5854 16558 5906
rect 16930 5854 16942 5906
rect 16994 5854 17006 5906
rect 17490 5869 17502 5921
rect 17554 5869 17566 5921
rect 17714 5854 17726 5906
rect 17778 5854 17790 5906
rect 18274 5854 18286 5906
rect 18338 5854 18350 5906
rect 18498 5898 18510 5950
rect 18562 5898 18574 5950
rect 18946 5854 18958 5906
rect 19010 5854 19022 5906
rect 19282 5898 19294 5950
rect 19346 5898 19358 5950
rect 19630 5906 19682 5918
rect 19630 5842 19682 5854
rect 23214 5906 23266 5918
rect 23214 5842 23266 5854
rect 23438 5906 23490 5918
rect 25342 5906 25394 5918
rect 26798 5906 26850 5918
rect 24302 5854 24314 5906
rect 24366 5854 24378 5906
rect 26206 5854 26218 5906
rect 26270 5854 26282 5906
rect 23438 5842 23490 5854
rect 25342 5842 25394 5854
rect 26798 5842 26850 5854
rect 27694 5906 27746 5918
rect 32062 5906 32114 5918
rect 28558 5854 28570 5906
rect 28622 5854 28634 5906
rect 31266 5854 31278 5906
rect 31330 5854 31342 5906
rect 27694 5842 27746 5854
rect 32062 5842 32114 5854
rect 33910 5906 33962 5918
rect 33910 5842 33962 5854
rect 34414 5906 34466 5918
rect 36542 5906 36594 5918
rect 35653 5854 35665 5906
rect 35717 5854 35729 5906
rect 37090 5898 37102 5950
rect 37154 5898 37166 5950
rect 37426 5854 37438 5906
rect 37490 5854 37502 5906
rect 40226 5881 40238 5933
rect 40290 5881 40302 5933
rect 40898 5854 40910 5906
rect 40962 5854 40974 5906
rect 41234 5869 41246 5921
rect 41298 5869 41310 5921
rect 41682 5881 41694 5933
rect 41746 5881 41758 5933
rect 34414 5842 34466 5854
rect 36542 5842 36594 5854
rect 17378 5742 17390 5794
rect 17442 5742 17454 5794
rect 18610 5742 18622 5794
rect 18674 5742 18686 5794
rect 19394 5742 19406 5794
rect 19458 5742 19470 5794
rect 20402 5742 20414 5794
rect 20466 5742 20478 5794
rect 22306 5742 22318 5794
rect 22370 5742 22382 5794
rect 39330 5742 39342 5794
rect 39394 5742 39406 5794
rect 41346 5742 41358 5794
rect 41410 5742 41422 5794
rect 42690 5742 42702 5794
rect 42754 5742 42766 5794
rect 16774 5682 16826 5694
rect 16774 5618 16826 5630
rect 22878 5682 22930 5694
rect 22878 5618 22930 5630
rect 27134 5682 27186 5694
rect 27134 5618 27186 5630
rect 34656 5682 34708 5694
rect 34656 5618 34708 5630
rect 1344 5514 44576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 44576 5514
rect 1344 5428 44576 5462
rect 43934 5346 43986 5358
rect 43934 5282 43986 5294
rect 15138 5182 15150 5234
rect 15202 5182 15214 5234
rect 17042 5182 17054 5234
rect 17106 5182 17118 5234
rect 20626 5182 20638 5234
rect 20690 5182 20702 5234
rect 22530 5182 22542 5234
rect 22594 5182 22606 5234
rect 24434 5182 24446 5234
rect 24498 5182 24510 5234
rect 24994 5182 25006 5234
rect 25058 5182 25070 5234
rect 26898 5182 26910 5234
rect 26962 5182 26974 5234
rect 29586 5182 29598 5234
rect 29650 5182 29662 5234
rect 31490 5182 31502 5234
rect 31554 5182 31566 5234
rect 35634 5182 35646 5234
rect 35698 5182 35710 5234
rect 39554 5182 39566 5234
rect 39618 5182 39630 5234
rect 43474 5182 43486 5234
rect 43538 5182 43550 5234
rect 17838 5122 17890 5134
rect 17838 5058 17890 5070
rect 17950 5122 18002 5134
rect 21758 5122 21810 5134
rect 18722 5070 18734 5122
rect 18786 5070 18798 5122
rect 21522 5070 21534 5122
rect 21586 5070 21598 5122
rect 17950 5058 18002 5070
rect 21758 5058 21810 5070
rect 27694 5122 27746 5134
rect 27694 5058 27746 5070
rect 28030 5122 28082 5134
rect 28030 5058 28082 5070
rect 28366 5122 28418 5134
rect 28366 5058 28418 5070
rect 32286 5122 32338 5134
rect 32286 5058 32338 5070
rect 32958 5122 33010 5134
rect 35982 5122 36034 5134
rect 33730 5070 33742 5122
rect 33794 5070 33806 5122
rect 32958 5058 33010 5070
rect 35982 5058 36034 5070
rect 36318 5122 36370 5134
rect 36318 5058 36370 5070
rect 36878 5122 36930 5134
rect 39902 5122 39954 5134
rect 44270 5122 44322 5134
rect 37650 5070 37662 5122
rect 37714 5070 37726 5122
rect 40674 5070 40686 5122
rect 40738 5070 40750 5122
rect 43026 5070 43038 5122
rect 43090 5070 43102 5122
rect 43318 5092 43370 5104
rect 36878 5058 36930 5070
rect 39902 5058 39954 5070
rect 44270 5058 44322 5070
rect 43318 5028 43370 5040
rect 42590 5010 42642 5022
rect 42590 4946 42642 4958
rect 21366 4898 21418 4910
rect 21366 4834 21418 4846
rect 1344 4730 44576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 44576 4730
rect 1344 4644 44576 4678
rect 38502 4562 38554 4574
rect 38502 4498 38554 4510
rect 28702 4450 28754 4462
rect 28702 4386 28754 4398
rect 29598 4450 29650 4462
rect 29598 4386 29650 4398
rect 30512 4450 30564 4462
rect 17602 4286 17614 4338
rect 17666 4286 17678 4338
rect 17938 4301 17950 4353
rect 18002 4301 18014 4353
rect 18286 4338 18338 4350
rect 18286 4274 18338 4286
rect 22206 4338 22258 4350
rect 22530 4301 22542 4353
rect 22594 4301 22606 4353
rect 26014 4338 26066 4350
rect 29754 4342 29766 4394
rect 29818 4342 29830 4394
rect 30512 4386 30564 4398
rect 36094 4450 36146 4462
rect 36094 4386 36146 4398
rect 36990 4450 37042 4462
rect 36990 4386 37042 4398
rect 39230 4450 39282 4462
rect 30270 4338 30322 4350
rect 22866 4286 22878 4338
rect 22930 4286 22942 4338
rect 26786 4286 26798 4338
rect 26850 4286 26862 4338
rect 22206 4274 22258 4286
rect 26014 4274 26066 4286
rect 30270 4274 30322 4286
rect 33406 4338 33458 4350
rect 37221 4342 37233 4394
rect 37285 4342 37297 4394
rect 39230 4386 39282 4398
rect 33406 4274 33458 4286
rect 38110 4338 38162 4350
rect 39461 4342 39473 4394
rect 39525 4342 39537 4394
rect 40350 4338 40402 4350
rect 38322 4286 38334 4338
rect 38386 4286 38398 4338
rect 38110 4274 38162 4286
rect 40350 4274 40402 4286
rect 44046 4338 44098 4350
rect 44046 4274 44098 4286
rect 18050 4174 18062 4226
rect 18114 4174 18126 4226
rect 19506 4174 19518 4226
rect 19570 4174 19582 4226
rect 21410 4174 21422 4226
rect 21474 4174 21486 4226
rect 22418 4174 22430 4226
rect 22482 4174 22494 4226
rect 34178 4174 34190 4226
rect 34242 4174 34254 4226
rect 41346 4174 41358 4226
rect 41410 4174 41422 4226
rect 43250 4174 43262 4226
rect 43314 4174 43326 4226
rect 1344 3946 44576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 44576 3946
rect 1344 3860 44576 3894
rect 17334 3778 17386 3790
rect 17334 3714 17386 3726
rect 25566 3778 25618 3790
rect 25566 3714 25618 3726
rect 29280 3778 29332 3790
rect 34638 3778 34690 3790
rect 32274 3726 32286 3778
rect 32338 3775 32350 3778
rect 33394 3775 33406 3778
rect 32338 3729 33406 3775
rect 32338 3726 32350 3729
rect 33394 3726 33406 3729
rect 33458 3726 33470 3778
rect 29280 3714 29332 3726
rect 34638 3714 34690 3726
rect 36766 3778 36818 3790
rect 36766 3714 36818 3726
rect 42870 3722 42922 3734
rect 27862 3666 27914 3678
rect 38502 3666 38554 3678
rect 27862 3602 27914 3614
rect 28534 3610 28586 3622
rect 18174 3554 18226 3566
rect 28366 3554 28418 3566
rect 17490 3502 17502 3554
rect 17554 3502 17566 3554
rect 18174 3490 18226 3502
rect 19842 3474 19854 3526
rect 19906 3474 19918 3526
rect 21074 3474 21086 3526
rect 21138 3474 21150 3526
rect 22978 3502 22990 3554
rect 23042 3502 23054 3554
rect 24546 3474 24558 3526
rect 24610 3474 24622 3526
rect 38770 3614 38782 3666
rect 38834 3614 38846 3666
rect 39890 3614 39902 3666
rect 39954 3614 39966 3666
rect 41794 3614 41806 3666
rect 41858 3614 41870 3666
rect 42870 3658 42922 3670
rect 43586 3614 43598 3666
rect 43650 3614 43662 3666
rect 38502 3602 38554 3614
rect 28534 3546 28586 3558
rect 29038 3554 29090 3566
rect 28366 3490 28418 3502
rect 29038 3490 29090 3502
rect 34302 3554 34354 3566
rect 34302 3490 34354 3502
rect 36430 3554 36482 3566
rect 42590 3554 42642 3566
rect 36430 3490 36482 3502
rect 38882 3487 38894 3539
rect 38946 3487 38958 3539
rect 39106 3502 39118 3554
rect 39170 3502 39182 3554
rect 42590 3490 42642 3502
rect 42702 3498 42754 3510
rect 43698 3487 43710 3539
rect 43762 3487 43774 3539
rect 43922 3502 43934 3554
rect 43986 3502 43998 3554
rect 42702 3434 42754 3446
rect 1344 3162 44576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 44576 3162
rect 1344 3076 44576 3110
<< via1 >>
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 41694 42142 41746 42194
rect 31278 41933 31330 41985
rect 31614 41918 31666 41970
rect 32286 41956 32338 42008
rect 32622 41918 32674 41970
rect 32846 41918 32898 41970
rect 33014 41862 33066 41914
rect 36878 41918 36930 41970
rect 37102 41918 37154 41970
rect 43038 41945 43090 41997
rect 31166 41806 31218 41858
rect 33630 41694 33682 41746
rect 34638 41694 34690 41746
rect 36598 41694 36650 41746
rect 37438 41694 37490 41746
rect 38334 41694 38386 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 35422 41358 35474 41410
rect 22990 41246 23042 41298
rect 26462 41246 26514 41298
rect 30942 41246 30994 41298
rect 33294 41246 33346 41298
rect 35982 41246 36034 41298
rect 37438 41246 37490 41298
rect 22542 41134 22594 41186
rect 22654 41134 22706 41186
rect 23102 41090 23154 41142
rect 23326 41134 23378 41186
rect 26014 41134 26066 41186
rect 26238 41134 26290 41186
rect 26574 41090 26626 41142
rect 26910 41134 26962 41186
rect 30158 41134 30210 41186
rect 33406 41119 33458 41171
rect 33630 41134 33682 41186
rect 35758 41134 35810 41186
rect 36094 41119 36146 41171
rect 36430 41134 36482 41186
rect 36990 41134 37042 41186
rect 37326 41119 37378 41171
rect 37662 41134 37714 41186
rect 22262 41022 22314 41074
rect 25734 41022 25786 41074
rect 32846 41022 32898 41074
rect 40798 41078 40850 41130
rect 41022 41078 41074 41130
rect 41246 41078 41298 41130
rect 41358 41078 41410 41130
rect 42030 41106 42082 41158
rect 40518 41022 40570 41074
rect 37998 40910 38050 40962
rect 43374 40910 43426 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 23942 40518 23994 40570
rect 28646 40462 28698 40514
rect 32398 40462 32450 40514
rect 33182 40462 33234 40514
rect 37774 40462 37826 40514
rect 20750 40350 20802 40402
rect 23438 40350 23490 40402
rect 23774 40350 23826 40402
rect 24782 40350 24834 40402
rect 25118 40350 25170 40402
rect 27806 40350 27858 40402
rect 28142 40350 28194 40402
rect 28366 40350 28418 40402
rect 33425 40406 33477 40458
rect 29710 40350 29762 40402
rect 34302 40350 34354 40402
rect 35086 40350 35138 40402
rect 35870 40350 35922 40402
rect 38110 40350 38162 40402
rect 38334 40350 38386 40402
rect 38614 40350 38666 40402
rect 39790 40350 39842 40402
rect 40462 40350 40514 40402
rect 40798 40350 40850 40402
rect 43486 40350 43538 40402
rect 21534 40238 21586 40290
rect 24446 40238 24498 40290
rect 25902 40238 25954 40290
rect 29206 40238 29258 40290
rect 30494 40238 30546 40290
rect 40126 40238 40178 40290
rect 41582 40238 41634 40290
rect 39454 40126 39506 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 40294 39790 40346 39842
rect 21870 39734 21922 39786
rect 23102 39734 23154 39786
rect 34302 39734 34354 39786
rect 43934 39790 43986 39842
rect 27358 39678 27410 39730
rect 28646 39678 28698 39730
rect 41358 39678 41410 39730
rect 21982 39566 22034 39618
rect 22318 39566 22370 39618
rect 22650 39528 22702 39580
rect 23326 39566 23378 39618
rect 24110 39566 24162 39618
rect 24894 39566 24946 39618
rect 27246 39566 27298 39618
rect 27918 39566 27970 39618
rect 27694 39510 27746 39562
rect 30270 39566 30322 39618
rect 31054 39566 31106 39618
rect 33742 39566 33794 39618
rect 33854 39566 33906 39618
rect 34190 39566 34242 39618
rect 34526 39566 34578 39618
rect 35758 39566 35810 39618
rect 35982 39527 36034 39579
rect 36318 39566 36370 39618
rect 36990 39566 37042 39618
rect 26798 39454 26850 39506
rect 37438 39527 37490 39579
rect 37662 39566 37714 39618
rect 39454 39510 39506 39562
rect 39566 39538 39618 39590
rect 39790 39538 39842 39590
rect 40014 39538 40066 39590
rect 40574 39566 40626 39618
rect 43598 39566 43650 39618
rect 32958 39454 33010 39506
rect 33462 39454 33514 39506
rect 43262 39454 43314 39506
rect 35646 39398 35698 39450
rect 37550 39398 37602 39450
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 32398 39006 32450 39058
rect 34974 39006 35026 39058
rect 22430 38894 22482 38946
rect 19742 38782 19794 38834
rect 22822 38838 22874 38890
rect 22990 38894 23042 38946
rect 24614 38894 24666 38946
rect 38110 38894 38162 38946
rect 23214 38782 23266 38834
rect 23438 38810 23490 38862
rect 24110 38782 24162 38834
rect 24334 38782 24386 38834
rect 25118 38782 25170 38834
rect 25902 38782 25954 38834
rect 28702 38782 28754 38834
rect 30382 38809 30434 38861
rect 31726 38782 31778 38834
rect 31950 38782 32002 38834
rect 32062 38782 32114 38834
rect 33126 38782 33178 38834
rect 33406 38782 33458 38834
rect 33630 38782 33682 38834
rect 35310 38782 35362 38834
rect 35422 38782 35474 38834
rect 36206 38782 36258 38834
rect 39454 38817 39506 38869
rect 39566 38838 39618 38890
rect 39790 38810 39842 38862
rect 40014 38810 40066 38862
rect 43710 38782 43762 38834
rect 20526 38670 20578 38722
rect 27806 38670 27858 38722
rect 31446 38670 31498 38722
rect 41022 38670 41074 38722
rect 42926 38670 42978 38722
rect 40294 38558 40346 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 29542 38222 29594 38274
rect 31334 38222 31386 38274
rect 21870 38166 21922 38218
rect 24894 38166 24946 38218
rect 26238 38166 26290 38218
rect 20302 38110 20354 38162
rect 31838 38110 31890 38162
rect 34190 38166 34242 38218
rect 43710 38222 43762 38274
rect 40574 38110 40626 38162
rect 20414 37954 20466 38006
rect 20750 37998 20802 38050
rect 21982 37998 22034 38050
rect 22318 37998 22370 38050
rect 22990 37998 23042 38050
rect 23102 37998 23154 38050
rect 23326 37998 23378 38050
rect 23550 37998 23602 38050
rect 23830 37998 23882 38050
rect 24110 37998 24162 38050
rect 24446 37998 24498 38050
rect 25006 37998 25058 38050
rect 25678 37998 25730 38050
rect 26238 37998 26290 38050
rect 26462 37998 26514 38050
rect 26966 37998 27018 38050
rect 27246 37998 27298 38050
rect 27470 37998 27522 38050
rect 27582 37998 27634 38050
rect 29038 37998 29090 38050
rect 29262 37998 29314 38050
rect 30830 37998 30882 38050
rect 31054 37998 31106 38050
rect 32174 37998 32226 38050
rect 34302 37998 34354 38050
rect 34638 37998 34690 38050
rect 36542 37998 36594 38050
rect 37438 37998 37490 38050
rect 38670 37998 38722 38050
rect 41358 37998 41410 38050
rect 41582 37963 41634 38015
rect 41694 37942 41746 37994
rect 41918 37970 41970 38022
rect 42422 37998 42474 38050
rect 42142 37942 42194 37994
rect 42702 37998 42754 38050
rect 43374 37998 43426 38050
rect 22710 37886 22762 37938
rect 37102 37886 37154 37938
rect 36374 37774 36426 37826
rect 43038 37774 43090 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 34862 37438 34914 37490
rect 39566 37438 39618 37490
rect 40238 37438 40290 37490
rect 23942 37326 23994 37378
rect 30718 37326 30770 37378
rect 19630 37214 19682 37266
rect 22318 37214 22370 37266
rect 22654 37214 22706 37266
rect 22878 37214 22930 37266
rect 23438 37214 23490 37266
rect 23662 37214 23714 37266
rect 27134 37214 27186 37266
rect 27246 37214 27298 37266
rect 27414 37214 27466 37266
rect 27582 37214 27634 37266
rect 28030 37214 28082 37266
rect 31502 37214 31554 37266
rect 31614 37214 31666 37266
rect 31838 37214 31890 37266
rect 32062 37214 32114 37266
rect 33182 37214 33234 37266
rect 33518 37214 33570 37266
rect 33854 37214 33906 37266
rect 34190 37214 34242 37266
rect 34526 37214 34578 37266
rect 35870 37214 35922 37266
rect 36094 37229 36146 37281
rect 36654 37229 36706 37281
rect 36990 37214 37042 37266
rect 37214 37214 37266 37266
rect 37886 37214 37938 37266
rect 39230 37214 39282 37266
rect 39902 37214 39954 37266
rect 40910 37214 40962 37266
rect 41694 37214 41746 37266
rect 20414 37102 20466 37154
rect 28814 37102 28866 37154
rect 33070 37046 33122 37098
rect 23158 36990 23210 37042
rect 26854 36990 26906 37042
rect 31222 36990 31274 37042
rect 32342 36990 32394 37042
rect 36206 37102 36258 37154
rect 36542 37102 36594 37154
rect 43598 37102 43650 37154
rect 34302 37046 34354 37098
rect 37550 36990 37602 37042
rect 38222 36990 38274 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 21758 36598 21810 36650
rect 29934 36654 29986 36706
rect 33742 36598 33794 36650
rect 20302 36542 20354 36594
rect 22150 36542 22202 36594
rect 37998 36542 38050 36594
rect 43150 36542 43202 36594
rect 12126 36430 12178 36482
rect 20414 36415 20466 36467
rect 20638 36430 20690 36482
rect 21422 36430 21474 36482
rect 21646 36430 21698 36482
rect 22430 36430 22482 36482
rect 22654 36430 22706 36482
rect 22766 36430 22818 36482
rect 22990 36430 23042 36482
rect 26910 36430 26962 36482
rect 29038 36430 29090 36482
rect 27786 36374 27838 36426
rect 30270 36430 30322 36482
rect 30550 36430 30602 36482
rect 30830 36430 30882 36482
rect 31054 36430 31106 36482
rect 31670 36430 31722 36482
rect 31950 36430 32002 36482
rect 32174 36430 32226 36482
rect 32958 36430 33010 36482
rect 33518 36430 33570 36482
rect 34134 36430 34186 36482
rect 34414 36430 34466 36482
rect 34526 36430 34578 36482
rect 34862 36430 34914 36482
rect 34694 36374 34746 36426
rect 37214 36402 37266 36454
rect 23270 36318 23322 36370
rect 28030 36318 28082 36370
rect 40798 36374 40850 36426
rect 41022 36402 41074 36454
rect 41246 36402 41298 36454
rect 41358 36374 41410 36426
rect 43822 36402 43874 36454
rect 40518 36318 40570 36370
rect 11790 36206 11842 36258
rect 15374 36206 15426 36258
rect 16662 36206 16714 36258
rect 29374 36206 29426 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 30718 35870 30770 35922
rect 16662 35758 16714 35810
rect 20190 35758 20242 35810
rect 26630 35758 26682 35810
rect 29598 35758 29650 35810
rect 34302 35758 34354 35810
rect 34694 35758 34746 35810
rect 9550 35646 9602 35698
rect 10426 35646 10478 35698
rect 11697 35646 11749 35698
rect 12574 35646 12626 35698
rect 13134 35646 13186 35698
rect 15822 35646 15874 35698
rect 16158 35646 16210 35698
rect 16382 35646 16434 35698
rect 17278 35646 17330 35698
rect 22878 35646 22930 35698
rect 26126 35646 26178 35698
rect 26350 35646 26402 35698
rect 26910 35646 26962 35698
rect 27694 35646 27746 35698
rect 31054 35646 31106 35698
rect 31838 35646 31890 35698
rect 32062 35646 32114 35698
rect 32398 35646 32450 35698
rect 33070 35646 33122 35698
rect 33182 35646 33234 35698
rect 33966 35646 34018 35698
rect 13918 35534 13970 35586
rect 22094 35534 22146 35586
rect 23270 35534 23322 35586
rect 25958 35534 26010 35586
rect 34134 35590 34186 35642
rect 34414 35646 34466 35698
rect 34974 35646 35026 35698
rect 35198 35646 35250 35698
rect 35478 35646 35530 35698
rect 37326 35674 37378 35726
rect 37550 35702 37602 35754
rect 37774 35702 37826 35754
rect 37886 35702 37938 35754
rect 39790 35646 39842 35698
rect 39902 35646 39954 35698
rect 40798 35646 40850 35698
rect 31502 35534 31554 35586
rect 33462 35534 33514 35586
rect 39454 35534 39506 35586
rect 41582 35534 41634 35586
rect 43486 35534 43538 35586
rect 10670 35422 10722 35474
rect 11454 35422 11506 35474
rect 17614 35422 17666 35474
rect 32510 35478 32562 35530
rect 37046 35422 37098 35474
rect 40238 35422 40290 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 21422 35086 21474 35138
rect 31614 35086 31666 35138
rect 43150 35086 43202 35138
rect 10334 34974 10386 35026
rect 27974 34974 28026 35026
rect 32398 34974 32450 35026
rect 36318 34974 36370 35026
rect 37102 34974 37154 35026
rect 40686 34974 40738 35026
rect 12238 34862 12290 34914
rect 13022 34862 13074 34914
rect 13358 34862 13410 34914
rect 15150 34862 15202 34914
rect 17390 34862 17442 34914
rect 18174 34862 18226 34914
rect 18286 34862 18338 34914
rect 18622 34862 18674 34914
rect 21758 34862 21810 34914
rect 25678 34862 25730 34914
rect 31950 34862 32002 34914
rect 34302 34862 34354 34914
rect 35086 34862 35138 34914
rect 35646 34862 35698 34914
rect 35758 34862 35810 34914
rect 35926 34862 35978 34914
rect 39006 34862 39058 34914
rect 39790 34862 39842 34914
rect 39902 34862 39954 34914
rect 43486 34862 43538 34914
rect 15486 34750 15538 34802
rect 42590 34750 42642 34802
rect 13694 34638 13746 34690
rect 14814 34638 14866 34690
rect 31222 34638 31274 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 26910 34302 26962 34354
rect 13694 34190 13746 34242
rect 33070 34190 33122 34242
rect 9102 34078 9154 34130
rect 9905 34078 9957 34130
rect 10782 34078 10834 34130
rect 11006 34078 11058 34130
rect 11790 34078 11842 34130
rect 14030 34078 14082 34130
rect 14814 34078 14866 34130
rect 17278 34078 17330 34130
rect 18062 34078 18114 34130
rect 24558 34078 24610 34130
rect 24782 34078 24834 34130
rect 25454 34078 25506 34130
rect 28254 34105 28306 34157
rect 31950 34078 32002 34130
rect 32286 34078 32338 34130
rect 33208 34118 33260 34170
rect 33518 34111 33570 34163
rect 33854 34114 33906 34166
rect 34190 34134 34242 34186
rect 34750 34078 34802 34130
rect 35086 34078 35138 34130
rect 35310 34078 35362 34130
rect 36766 34106 36818 34158
rect 36990 34134 37042 34186
rect 37214 34106 37266 34158
rect 37326 34134 37378 34186
rect 37886 34105 37938 34157
rect 40798 34078 40850 34130
rect 41582 34078 41634 34130
rect 16718 33966 16770 34018
rect 19966 33966 20018 34018
rect 8766 33854 8818 33906
rect 9662 33854 9714 33906
rect 24278 33854 24330 33906
rect 25286 33854 25338 33906
rect 32398 33910 32450 33962
rect 43486 33966 43538 34018
rect 34638 33910 34690 33962
rect 35646 33854 35698 33906
rect 36486 33854 36538 33906
rect 38894 33854 38946 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 12294 33518 12346 33570
rect 15822 33518 15874 33570
rect 16774 33518 16826 33570
rect 17558 33518 17610 33570
rect 27694 33518 27746 33570
rect 28590 33462 28642 33514
rect 42814 33518 42866 33570
rect 8766 33406 8818 33458
rect 9886 33406 9938 33458
rect 11790 33406 11842 33458
rect 24222 33406 24274 33458
rect 26126 33406 26178 33458
rect 31614 33406 31666 33458
rect 6078 33294 6130 33346
rect 6862 33294 6914 33346
rect 9102 33294 9154 33346
rect 12462 33294 12514 33346
rect 16158 33294 16210 33346
rect 16382 33294 16434 33346
rect 16494 33294 16546 33346
rect 17054 33294 17106 33346
rect 17278 33294 17330 33346
rect 20078 33294 20130 33346
rect 20862 33294 20914 33346
rect 22990 33294 23042 33346
rect 23438 33294 23490 33346
rect 26574 33294 26626 33346
rect 27450 33294 27502 33346
rect 28142 33294 28194 33346
rect 28478 33294 28530 33346
rect 18174 33182 18226 33234
rect 29094 33238 29146 33290
rect 29262 33238 29314 33290
rect 29486 33255 29538 33307
rect 30046 33294 30098 33346
rect 31278 33294 31330 33346
rect 31502 33279 31554 33331
rect 32174 33294 32226 33346
rect 34414 33266 34466 33318
rect 34862 33294 34914 33346
rect 35534 33294 35586 33346
rect 37326 33266 37378 33318
rect 37550 33266 37602 33318
rect 37718 33259 37770 33311
rect 38110 33294 38162 33346
rect 39454 33294 39506 33346
rect 40238 33294 40290 33346
rect 42478 33294 42530 33346
rect 23158 33126 23210 33178
rect 37046 33182 37098 33234
rect 37886 33238 37938 33290
rect 43710 33294 43762 33346
rect 42142 33182 42194 33234
rect 35198 33070 35250 33122
rect 35870 33070 35922 33122
rect 36486 33070 36538 33122
rect 43374 33070 43426 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 20078 32734 20130 32786
rect 6414 32622 6466 32674
rect 25398 32678 25450 32730
rect 38334 32734 38386 32786
rect 38838 32734 38890 32786
rect 12238 32622 12290 32674
rect 19126 32622 19178 32674
rect 34022 32622 34074 32674
rect 9102 32510 9154 32562
rect 9550 32510 9602 32562
rect 10334 32510 10386 32562
rect 17726 32510 17778 32562
rect 17950 32510 18002 32562
rect 19406 32510 19458 32562
rect 19630 32510 19682 32562
rect 19742 32510 19794 32562
rect 20862 32510 20914 32562
rect 21646 32510 21698 32562
rect 24334 32510 24386 32562
rect 24558 32510 24610 32562
rect 25230 32510 25282 32562
rect 25678 32510 25730 32562
rect 28366 32510 28418 32562
rect 29038 32510 29090 32562
rect 30606 32510 30658 32562
rect 30718 32510 30770 32562
rect 30904 32547 30956 32599
rect 31726 32510 31778 32562
rect 31838 32510 31890 32562
rect 31984 32547 32036 32599
rect 34582 32566 34634 32618
rect 34750 32566 34802 32618
rect 37662 32622 37714 32674
rect 39510 32622 39562 32674
rect 33406 32510 33458 32562
rect 34302 32510 34354 32562
rect 34414 32510 34466 32562
rect 39790 32566 39842 32618
rect 34974 32510 35026 32562
rect 35758 32510 35810 32562
rect 37998 32510 38050 32562
rect 38670 32510 38722 32562
rect 40014 32538 40066 32590
rect 40182 32545 40234 32597
rect 40350 32566 40402 32618
rect 43822 32537 43874 32589
rect 8318 32398 8370 32450
rect 23550 32398 23602 32450
rect 26462 32398 26514 32450
rect 24670 32342 24722 32394
rect 17446 32286 17498 32338
rect 43150 32398 43202 32450
rect 28870 32342 28922 32394
rect 31278 32286 31330 32338
rect 32398 32286 32450 32338
rect 33574 32286 33626 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 18062 31838 18114 31890
rect 29654 31894 29706 31946
rect 34078 31950 34130 32002
rect 34582 31950 34634 32002
rect 18846 31838 18898 31890
rect 23886 31838 23938 31890
rect 24726 31838 24778 31890
rect 27918 31838 27970 31890
rect 33182 31838 33234 31890
rect 42254 31838 42306 31890
rect 15038 31726 15090 31778
rect 15598 31726 15650 31778
rect 15710 31726 15762 31778
rect 16830 31726 16882 31778
rect 17726 31726 17778 31778
rect 18398 31726 18450 31778
rect 18510 31726 18562 31778
rect 21198 31726 21250 31778
rect 21982 31726 22034 31778
rect 25006 31670 25058 31722
rect 25230 31670 25282 31722
rect 25454 31698 25506 31750
rect 25622 31710 25674 31762
rect 28702 31726 28754 31778
rect 29038 31726 29090 31778
rect 29486 31726 29538 31778
rect 30270 31726 30322 31778
rect 35142 31782 35194 31834
rect 31390 31726 31442 31778
rect 31838 31726 31890 31778
rect 32174 31726 32226 31778
rect 32734 31726 32786 31778
rect 32958 31726 33010 31778
rect 33406 31726 33458 31778
rect 33518 31726 33570 31778
rect 34862 31726 34914 31778
rect 34974 31726 35026 31778
rect 35310 31726 35362 31778
rect 31146 31670 31198 31722
rect 33686 31670 33738 31722
rect 35534 31726 35586 31778
rect 35758 31726 35810 31778
rect 39566 31726 39618 31778
rect 40350 31726 40402 31778
rect 15318 31614 15370 31666
rect 26014 31614 26066 31666
rect 36038 31614 36090 31666
rect 14702 31502 14754 31554
rect 16494 31502 16546 31554
rect 17390 31502 17442 31554
rect 29206 31502 29258 31554
rect 42870 31502 42922 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 18398 31166 18450 31218
rect 30326 31166 30378 31218
rect 15374 31054 15426 31106
rect 17446 31054 17498 31106
rect 28982 31054 29034 31106
rect 29598 31054 29650 31106
rect 37662 31054 37714 31106
rect 12686 30942 12738 30994
rect 13470 30942 13522 30994
rect 16270 30942 16322 30994
rect 16494 30942 16546 30994
rect 17726 30942 17778 30994
rect 17838 30942 17890 30994
rect 18062 30942 18114 30994
rect 20078 30962 20130 31014
rect 20190 30942 20242 30994
rect 20974 30942 21026 30994
rect 22878 30942 22930 30994
rect 25454 30942 25506 30994
rect 25790 30942 25842 30994
rect 26126 30969 26178 31021
rect 26462 30942 26514 30994
rect 26798 30942 26850 30994
rect 27246 30981 27298 31033
rect 27470 30942 27522 30994
rect 27806 30942 27858 30994
rect 28478 30942 28530 30994
rect 28702 30942 28754 30994
rect 29262 30942 29314 30994
rect 30158 30942 30210 30994
rect 30606 30942 30658 30994
rect 31614 30998 31666 31050
rect 31726 30998 31778 31050
rect 31950 30998 32002 31050
rect 30830 30942 30882 30994
rect 31110 30942 31162 30994
rect 32174 30970 32226 31022
rect 33070 30942 33122 30994
rect 33182 30942 33234 30994
rect 33350 30942 33402 30994
rect 34190 30942 34242 30994
rect 34526 30942 34578 30994
rect 34974 30942 35026 30994
rect 35758 30942 35810 30994
rect 41470 30942 41522 30994
rect 42366 30942 42418 30994
rect 26238 30830 26290 30882
rect 27134 30830 27186 30882
rect 16774 30718 16826 30770
rect 19910 30718 19962 30770
rect 32454 30718 32506 30770
rect 34414 30774 34466 30826
rect 33742 30718 33794 30770
rect 41302 30718 41354 30770
rect 42702 30718 42754 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 20638 30382 20690 30434
rect 28086 30382 28138 30434
rect 32734 30382 32786 30434
rect 33854 30382 33906 30434
rect 17838 30270 17890 30322
rect 19742 30270 19794 30322
rect 21982 30270 22034 30322
rect 40462 30270 40514 30322
rect 13918 30158 13970 30210
rect 14030 30158 14082 30210
rect 14814 30158 14866 30210
rect 16718 30158 16770 30210
rect 17054 30158 17106 30210
rect 20302 30158 20354 30210
rect 21198 30158 21250 30210
rect 23886 30158 23938 30210
rect 24222 30158 24274 30210
rect 25006 30158 25058 30210
rect 25230 30158 25282 30210
rect 25510 30158 25562 30210
rect 26350 30158 26402 30210
rect 27246 30123 27298 30175
rect 27414 30123 27466 30175
rect 27638 30123 27690 30175
rect 27862 30123 27914 30175
rect 31614 30158 31666 30210
rect 33182 30158 33234 30210
rect 33294 30158 33346 30210
rect 33462 30158 33514 30210
rect 32490 30102 32542 30154
rect 37774 30158 37826 30210
rect 38110 30158 38162 30210
rect 38558 30158 38610 30210
rect 39678 30158 39730 30210
rect 42366 30158 42418 30210
rect 13582 29934 13634 29986
rect 24558 29934 24610 29986
rect 26686 29934 26738 29986
rect 37606 29934 37658 29986
rect 38894 29934 38946 29986
rect 39510 29934 39562 29986
rect 42982 29934 43034 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 18622 29598 18674 29650
rect 25902 29598 25954 29650
rect 26686 29598 26738 29650
rect 27246 29598 27298 29650
rect 43374 29598 43426 29650
rect 16158 29486 16210 29538
rect 18118 29486 18170 29538
rect 19742 29486 19794 29538
rect 32398 29486 32450 29538
rect 13470 29374 13522 29426
rect 14254 29374 14306 29426
rect 17726 29374 17778 29426
rect 17838 29374 17890 29426
rect 18958 29374 19010 29426
rect 21646 29374 21698 29426
rect 22430 29374 22482 29426
rect 22822 29374 22874 29426
rect 23550 29374 23602 29426
rect 24222 29374 24274 29426
rect 25566 29374 25618 29426
rect 31278 29374 31330 29426
rect 32154 29374 32206 29426
rect 36318 29374 36370 29426
rect 36878 29374 36930 29426
rect 37214 29374 37266 29426
rect 37438 29389 37490 29441
rect 40014 29401 40066 29453
rect 40910 29374 40962 29426
rect 41246 29389 41298 29441
rect 41918 29401 41970 29453
rect 37550 29262 37602 29314
rect 39342 29262 39394 29314
rect 41358 29262 41410 29314
rect 23214 29150 23266 29202
rect 23886 29150 23938 29202
rect 36150 29150 36202 29202
rect 36710 29150 36762 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 25902 28814 25954 28866
rect 31894 28814 31946 28866
rect 31054 28758 31106 28810
rect 15934 28702 15986 28754
rect 17838 28702 17890 28754
rect 35870 28702 35922 28754
rect 36990 28702 37042 28754
rect 38670 28702 38722 28754
rect 43598 28702 43650 28754
rect 15150 28590 15202 28642
rect 20862 28590 20914 28642
rect 21310 28590 21362 28642
rect 22186 28590 22238 28642
rect 24110 28590 24162 28642
rect 24222 28590 24274 28642
rect 24558 28590 24610 28642
rect 25566 28590 25618 28642
rect 26238 28590 26290 28642
rect 26462 28590 26514 28642
rect 26798 28575 26850 28627
rect 27246 28590 27298 28642
rect 27582 28575 27634 28627
rect 30830 28590 30882 28642
rect 31054 28590 31106 28642
rect 31390 28590 31442 28642
rect 31614 28590 31666 28642
rect 34750 28562 34802 28614
rect 35422 28590 35474 28642
rect 35758 28546 35810 28598
rect 36430 28590 36482 28642
rect 37102 28546 37154 28598
rect 37326 28590 37378 28642
rect 37886 28590 37938 28642
rect 40910 28590 40962 28642
rect 41694 28590 41746 28642
rect 22430 28478 22482 28530
rect 40574 28478 40626 28530
rect 20526 28366 20578 28418
rect 23774 28366 23826 28418
rect 26574 28422 26626 28474
rect 27358 28422 27410 28474
rect 25230 28366 25282 28418
rect 33742 28366 33794 28418
rect 36262 28366 36314 28418
rect 44214 28366 44266 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 16494 28030 16546 28082
rect 31166 28030 31218 28082
rect 24110 27918 24162 27970
rect 33966 27974 34018 28026
rect 28254 27918 28306 27970
rect 34526 27918 34578 27970
rect 11790 27806 11842 27858
rect 16830 27806 16882 27858
rect 21422 27806 21474 27858
rect 22206 27806 22258 27858
rect 24726 27806 24778 27858
rect 25566 27806 25618 27858
rect 26350 27806 26402 27858
rect 28814 27850 28866 27902
rect 29150 27806 29202 27858
rect 29822 27806 29874 27858
rect 32510 27833 32562 27885
rect 33742 27850 33794 27902
rect 34078 27806 34130 27858
rect 36430 27806 36482 27858
rect 37214 27806 37266 27858
rect 39678 27806 39730 27858
rect 40462 27806 40514 27858
rect 41134 27806 41186 27858
rect 28702 27694 28754 27746
rect 37774 27694 37826 27746
rect 41918 27694 41970 27746
rect 43822 27694 43874 27746
rect 11622 27582 11674 27634
rect 29654 27582 29706 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 14142 27246 14194 27298
rect 20526 27246 20578 27298
rect 21422 27246 21474 27298
rect 22598 27246 22650 27298
rect 37998 27246 38050 27298
rect 27806 27190 27858 27242
rect 40854 27246 40906 27298
rect 12798 27134 12850 27186
rect 15598 27134 15650 27186
rect 23662 27134 23714 27186
rect 25566 27134 25618 27186
rect 30270 27134 30322 27186
rect 32174 27134 32226 27186
rect 33406 27134 33458 27186
rect 34414 27134 34466 27186
rect 36318 27134 36370 27186
rect 10110 27022 10162 27074
rect 10894 27022 10946 27074
rect 14478 27022 14530 27074
rect 16046 27022 16098 27074
rect 16606 27022 16658 27074
rect 19462 27022 19514 27074
rect 15766 26966 15818 27018
rect 19854 27022 19906 27074
rect 20190 27022 20242 27074
rect 20862 27022 20914 27074
rect 21758 27022 21810 27074
rect 22878 27022 22930 27074
rect 23102 27022 23154 27074
rect 26350 27022 26402 27074
rect 26574 27022 26626 27074
rect 27246 27022 27298 27074
rect 28030 27022 28082 27074
rect 28590 27022 28642 27074
rect 26910 26966 26962 27018
rect 29486 27022 29538 27074
rect 32958 27022 33010 27074
rect 33294 27007 33346 27059
rect 33630 27022 33682 27074
rect 36990 26994 37042 27046
rect 39678 27022 39730 27074
rect 40686 27022 40738 27074
rect 41134 27022 41186 27074
rect 41918 27022 41970 27074
rect 16774 26854 16826 26906
rect 22150 26910 22202 26962
rect 43822 26910 43874 26962
rect 26686 26854 26738 26906
rect 18566 26798 18618 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 9718 26462 9770 26514
rect 22318 26462 22370 26514
rect 16494 26350 16546 26402
rect 26238 26406 26290 26458
rect 33238 26462 33290 26514
rect 40182 26462 40234 26514
rect 42254 26462 42306 26514
rect 29710 26350 29762 26402
rect 9886 26238 9938 26290
rect 10222 26238 10274 26290
rect 10446 26282 10498 26334
rect 10782 26238 10834 26290
rect 13806 26238 13858 26290
rect 14590 26238 14642 26290
rect 17278 26238 17330 26290
rect 17838 26238 17890 26290
rect 18118 26267 18170 26319
rect 18734 26238 18786 26290
rect 19070 26238 19122 26290
rect 19742 26238 19794 26290
rect 20078 26238 20130 26290
rect 20414 26282 20466 26334
rect 37774 26350 37826 26402
rect 20794 26276 20846 26328
rect 21534 26238 21586 26290
rect 22654 26238 22706 26290
rect 23102 26238 23154 26290
rect 25118 26238 25170 26290
rect 25454 26238 25506 26290
rect 26014 26238 26066 26290
rect 26350 26277 26402 26329
rect 26574 26238 26626 26290
rect 27022 26238 27074 26290
rect 30942 26238 30994 26290
rect 32174 26282 32226 26334
rect 32510 26238 32562 26290
rect 33070 26238 33122 26290
rect 33630 26238 33682 26290
rect 34506 26238 34558 26290
rect 35086 26238 35138 26290
rect 35870 26238 35922 26290
rect 38558 26238 38610 26290
rect 39434 26238 39486 26290
rect 40350 26238 40402 26290
rect 41246 26265 41298 26317
rect 43878 26294 43930 26346
rect 44046 26294 44098 26346
rect 10558 26126 10610 26178
rect 11566 26126 11618 26178
rect 13470 26126 13522 26178
rect 18286 26126 18338 26178
rect 20526 26126 20578 26178
rect 27806 26126 27858 26178
rect 32062 26126 32114 26178
rect 43710 26126 43762 26178
rect 17446 26014 17498 26066
rect 19406 26014 19458 26066
rect 21646 26070 21698 26122
rect 22934 26014 22986 26066
rect 30606 26014 30658 26066
rect 34750 26014 34802 26066
rect 39678 26014 39730 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 14086 25622 14138 25674
rect 28142 25678 28194 25730
rect 36206 25678 36258 25730
rect 17054 25566 17106 25618
rect 18174 25566 18226 25618
rect 21982 25566 22034 25618
rect 23886 25566 23938 25618
rect 30718 25566 30770 25618
rect 32622 25566 32674 25618
rect 37998 25566 38050 25618
rect 40798 25566 40850 25618
rect 12238 25454 12290 25506
rect 13022 25454 13074 25506
rect 13806 25454 13858 25506
rect 10334 25342 10386 25394
rect 14254 25398 14306 25450
rect 14366 25454 14418 25506
rect 15150 25454 15202 25506
rect 17446 25454 17498 25506
rect 20862 25454 20914 25506
rect 21198 25454 21250 25506
rect 25566 25454 25618 25506
rect 26126 25454 26178 25506
rect 26686 25454 26738 25506
rect 27358 25454 27410 25506
rect 25902 25398 25954 25450
rect 27022 25398 27074 25450
rect 27806 25454 27858 25506
rect 29934 25454 29986 25506
rect 33294 25426 33346 25478
rect 36542 25454 36594 25506
rect 36990 25426 37042 25478
rect 39790 25426 39842 25478
rect 43822 25454 43874 25506
rect 20078 25342 20130 25394
rect 42945 25398 42997 25450
rect 29766 25342 29818 25394
rect 34974 25342 35026 25394
rect 42702 25342 42754 25394
rect 13638 25230 13690 25282
rect 25566 25286 25618 25338
rect 27470 25286 27522 25338
rect 20694 25230 20746 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 13526 24894 13578 24946
rect 37438 24894 37490 24946
rect 42366 24894 42418 24946
rect 19966 24782 20018 24834
rect 28646 24782 28698 24834
rect 13022 24697 13074 24749
rect 13358 24670 13410 24722
rect 14030 24670 14082 24722
rect 17278 24670 17330 24722
rect 23774 24697 23826 24749
rect 24782 24670 24834 24722
rect 25454 24697 25506 24749
rect 28142 24670 28194 24722
rect 28366 24670 28418 24722
rect 29262 24670 29314 24722
rect 29374 24670 29426 24722
rect 32510 24697 32562 24749
rect 32958 24670 33010 24722
rect 33742 24670 33794 24722
rect 36094 24697 36146 24749
rect 39118 24670 39170 24722
rect 39994 24670 40046 24722
rect 41022 24697 41074 24749
rect 44270 24670 44322 24722
rect 14814 24558 14866 24610
rect 16718 24558 16770 24610
rect 18062 24558 18114 24610
rect 35646 24558 35698 24610
rect 11678 24446 11730 24498
rect 22206 24446 22258 24498
rect 24446 24446 24498 24498
rect 26462 24446 26514 24498
rect 29654 24446 29706 24498
rect 31502 24446 31554 24498
rect 40238 24446 40290 24498
rect 43934 24446 43986 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 11062 24110 11114 24162
rect 19518 24110 19570 24162
rect 10278 23998 10330 24050
rect 11454 23998 11506 24050
rect 12238 23998 12290 24050
rect 15598 23998 15650 24050
rect 16830 23998 16882 24050
rect 18622 23998 18674 24050
rect 21982 23998 22034 24050
rect 23886 23998 23938 24050
rect 25342 23998 25394 24050
rect 30158 23998 30210 24050
rect 33630 23998 33682 24050
rect 35982 23998 36034 24050
rect 41022 23998 41074 24050
rect 10894 23886 10946 23938
rect 10782 23830 10834 23882
rect 11566 23842 11618 23894
rect 11902 23886 11954 23938
rect 12350 23871 12402 23923
rect 12686 23886 12738 23938
rect 15710 23871 15762 23923
rect 16046 23886 16098 23938
rect 16942 23871 16994 23923
rect 17166 23886 17218 23938
rect 18790 23856 18842 23908
rect 18958 23886 19010 23938
rect 19854 23886 19906 23938
rect 21198 23886 21250 23938
rect 24558 23886 24610 23938
rect 28702 23886 28754 23938
rect 29150 23858 29202 23910
rect 31838 23886 31890 23938
rect 32846 23886 32898 23938
rect 35534 23886 35586 23938
rect 36150 23856 36202 23908
rect 36318 23886 36370 23938
rect 37550 23886 37602 23938
rect 38222 23886 38274 23938
rect 39790 23886 39842 23938
rect 37942 23830 37994 23882
rect 27246 23774 27298 23826
rect 38913 23830 38965 23882
rect 40350 23886 40402 23938
rect 40686 23886 40738 23938
rect 40910 23847 40962 23899
rect 41246 23886 41298 23938
rect 41694 23858 41746 23910
rect 38670 23774 38722 23826
rect 10614 23662 10666 23714
rect 37662 23718 37714 23770
rect 32174 23662 32226 23714
rect 43374 23662 43426 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 32398 23326 32450 23378
rect 33126 23326 33178 23378
rect 33574 23326 33626 23378
rect 9662 23102 9714 23154
rect 9886 23146 9938 23198
rect 10558 23146 10610 23198
rect 10894 23102 10946 23154
rect 13694 23129 13746 23181
rect 14478 23102 14530 23154
rect 15710 23102 15762 23154
rect 16830 23102 16882 23154
rect 20582 23158 20634 23210
rect 20862 23130 20914 23182
rect 21086 23158 21138 23210
rect 21198 23158 21250 23210
rect 27806 23214 27858 23266
rect 31054 23214 31106 23266
rect 21758 23102 21810 23154
rect 23998 23129 24050 23181
rect 28702 23158 28754 23210
rect 25118 23102 25170 23154
rect 28142 23102 28194 23154
rect 28814 23130 28866 23182
rect 29038 23130 29090 23182
rect 29262 23158 29314 23210
rect 29934 23102 29986 23154
rect 30810 23102 30862 23154
rect 31390 23102 31442 23154
rect 32062 23102 32114 23154
rect 33294 23102 33346 23154
rect 33742 23102 33794 23154
rect 34862 23102 34914 23154
rect 35738 23102 35790 23154
rect 36430 23102 36482 23154
rect 37306 23102 37358 23154
rect 37550 23102 37602 23154
rect 37998 23102 38050 23154
rect 38334 23129 38386 23181
rect 38670 23102 38722 23154
rect 39006 23102 39058 23154
rect 39454 23102 39506 23154
rect 40462 23102 40514 23154
rect 41022 23102 41074 23154
rect 41358 23117 41410 23169
rect 42161 23102 42213 23154
rect 43038 23102 43090 23154
rect 43486 23146 43538 23198
rect 43822 23102 43874 23154
rect 9998 22990 10050 23042
rect 10446 22990 10498 23042
rect 25902 22990 25954 23042
rect 38110 22990 38162 23042
rect 41470 22990 41522 23042
rect 43374 22990 43426 23042
rect 12686 22878 12738 22930
rect 14142 22878 14194 22930
rect 15374 22878 15426 22930
rect 16494 22878 16546 22930
rect 17502 22878 17554 22930
rect 18286 22878 18338 22930
rect 20358 22878 20410 22930
rect 28310 22934 28362 22986
rect 29542 22878 29594 22930
rect 31726 22878 31778 22930
rect 35982 22878 36034 22930
rect 39790 22878 39842 22930
rect 40294 22878 40346 22930
rect 41918 22878 41970 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 16158 22542 16210 22594
rect 19630 22542 19682 22594
rect 22654 22542 22706 22594
rect 24446 22542 24498 22594
rect 36206 22542 36258 22594
rect 38110 22542 38162 22594
rect 42926 22542 42978 22594
rect 10894 22430 10946 22482
rect 12798 22430 12850 22482
rect 26238 22430 26290 22482
rect 27694 22430 27746 22482
rect 29150 22430 29202 22482
rect 38670 22430 38722 22482
rect 9774 22290 9826 22342
rect 10110 22318 10162 22370
rect 13582 22318 13634 22370
rect 14458 22262 14510 22314
rect 15150 22290 15202 22342
rect 19873 22318 19925 22370
rect 20750 22318 20802 22370
rect 22318 22318 22370 22370
rect 23550 22290 23602 22342
rect 26350 22274 26402 22326
rect 26686 22318 26738 22370
rect 27470 22318 27522 22370
rect 27750 22288 27802 22340
rect 28030 22318 28082 22370
rect 29262 22274 29314 22326
rect 29598 22318 29650 22370
rect 29934 22318 29986 22370
rect 30810 22318 30862 22370
rect 31950 22318 32002 22370
rect 34190 22318 34242 22370
rect 35086 22318 35138 22370
rect 36990 22318 37042 22370
rect 38558 22318 38610 22370
rect 39230 22318 39282 22370
rect 14702 22206 14754 22258
rect 35962 22262 36014 22314
rect 37866 22262 37918 22314
rect 38838 22262 38890 22314
rect 39678 22318 39730 22370
rect 40462 22318 40514 22370
rect 44046 22318 44098 22370
rect 31054 22206 31106 22258
rect 43169 22262 43221 22314
rect 42366 22206 42418 22258
rect 8430 22094 8482 22146
rect 27134 22094 27186 22146
rect 28646 22094 28698 22146
rect 31614 22094 31666 22146
rect 32342 22094 32394 22146
rect 33854 22094 33906 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 17950 21758 18002 21810
rect 19294 21758 19346 21810
rect 32006 21758 32058 21810
rect 28478 21702 28530 21754
rect 29206 21646 29258 21698
rect 37774 21646 37826 21698
rect 8094 21534 8146 21586
rect 8542 21534 8594 21586
rect 9438 21534 9490 21586
rect 10222 21534 10274 21586
rect 12574 21534 12626 21586
rect 13450 21534 13502 21586
rect 16158 21534 16210 21586
rect 16942 21534 16994 21586
rect 17614 21534 17666 21586
rect 18398 21534 18450 21586
rect 19630 21534 19682 21586
rect 20209 21534 20261 21586
rect 21086 21534 21138 21586
rect 24110 21534 24162 21586
rect 24334 21534 24386 21586
rect 25454 21561 25506 21613
rect 28366 21578 28418 21630
rect 29766 21590 29818 21642
rect 43822 21646 43874 21698
rect 28702 21534 28754 21586
rect 29486 21534 29538 21586
rect 29598 21534 29650 21586
rect 29934 21534 29986 21586
rect 30382 21534 30434 21586
rect 31122 21572 31174 21624
rect 32958 21534 33010 21586
rect 39678 21534 39730 21586
rect 40462 21534 40514 21586
rect 41134 21534 41186 21586
rect 12126 21422 12178 21474
rect 14254 21422 14306 21474
rect 26462 21422 26514 21474
rect 31558 21422 31610 21474
rect 33742 21422 33794 21474
rect 35646 21422 35698 21474
rect 41918 21422 41970 21474
rect 8262 21366 8314 21418
rect 8878 21310 8930 21362
rect 13694 21310 13746 21362
rect 18734 21310 18786 21362
rect 30606 21366 30658 21418
rect 19966 21310 20018 21362
rect 23830 21310 23882 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 18268 20974 18320 21026
rect 25398 20974 25450 21026
rect 29374 20974 29426 21026
rect 32062 20974 32114 21026
rect 12238 20862 12290 20914
rect 8206 20750 8258 20802
rect 8990 20750 9042 20802
rect 9102 20750 9154 20802
rect 9886 20750 9938 20802
rect 12350 20706 12402 20758
rect 12574 20750 12626 20802
rect 13582 20750 13634 20802
rect 14458 20750 14510 20802
rect 17166 20750 17218 20802
rect 17950 20750 18002 20802
rect 18510 20750 18562 20802
rect 19014 20806 19066 20858
rect 21404 20862 21456 20914
rect 30718 20918 30770 20970
rect 42254 20974 42306 21026
rect 20862 20750 20914 20802
rect 21646 20750 21698 20802
rect 22150 20806 22202 20858
rect 22822 20862 22874 20914
rect 26910 20862 26962 20914
rect 28142 20862 28194 20914
rect 33294 20862 33346 20914
rect 35198 20862 35250 20914
rect 24670 20750 24722 20802
rect 24838 20806 24890 20858
rect 25118 20750 25170 20802
rect 26574 20750 26626 20802
rect 27022 20706 27074 20758
rect 27246 20750 27298 20802
rect 27694 20750 27746 20802
rect 28030 20706 28082 20758
rect 29710 20750 29762 20802
rect 29934 20750 29986 20802
rect 30494 20750 30546 20802
rect 32398 20750 32450 20802
rect 32510 20750 32562 20802
rect 38614 20806 38666 20858
rect 39360 20862 39412 20914
rect 39118 20750 39170 20802
rect 40126 20750 40178 20802
rect 40630 20806 40682 20858
rect 41302 20750 41354 20802
rect 42590 20750 42642 20802
rect 42908 20750 42960 20802
rect 43150 20750 43202 20802
rect 43654 20806 43706 20858
rect 6302 20638 6354 20690
rect 11790 20638 11842 20690
rect 14702 20638 14754 20690
rect 15262 20638 15314 20690
rect 19182 20638 19234 20690
rect 22318 20638 22370 20690
rect 25006 20638 25058 20690
rect 39884 20638 39936 20690
rect 19686 20526 19738 20578
rect 20526 20526 20578 20578
rect 28646 20526 28698 20578
rect 31334 20526 31386 20578
rect 38782 20582 38834 20634
rect 40798 20638 40850 20690
rect 35814 20526 35866 20578
rect 43598 20582 43650 20634
rect 41862 20526 41914 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 13358 20190 13410 20242
rect 17614 20190 17666 20242
rect 25342 20190 25394 20242
rect 12126 20078 12178 20130
rect 15822 20078 15874 20130
rect 28366 20134 28418 20186
rect 21870 20078 21922 20130
rect 26854 20078 26906 20130
rect 29934 20078 29986 20130
rect 33164 20078 33216 20130
rect 35086 20134 35138 20186
rect 34508 20078 34560 20130
rect 8430 19981 8482 20033
rect 8766 19966 8818 20018
rect 9438 19966 9490 20018
rect 10222 19966 10274 20018
rect 14702 19993 14754 20045
rect 15990 19910 16042 19962
rect 16494 19966 16546 20018
rect 16736 19966 16788 20018
rect 17278 19966 17330 20018
rect 19182 19966 19234 20018
rect 19966 19966 20018 20018
rect 22206 19966 22258 20018
rect 24278 19966 24330 20018
rect 25678 19966 25730 20018
rect 26350 19966 26402 20018
rect 27134 19966 27186 20018
rect 27358 19966 27410 20018
rect 27470 19966 27522 20018
rect 28254 19966 28306 20018
rect 28702 20005 28754 20057
rect 28926 19966 28978 20018
rect 33910 20022 33962 20074
rect 40238 20078 40290 20130
rect 30270 19966 30322 20018
rect 30718 19966 30770 20018
rect 31390 19966 31442 20018
rect 33406 19966 33458 20018
rect 34078 19966 34130 20018
rect 35254 20022 35306 20074
rect 34750 19966 34802 20018
rect 38670 19966 38722 20018
rect 39902 19966 39954 20018
rect 40798 19966 40850 20018
rect 41694 19966 41746 20018
rect 42926 19966 42978 20018
rect 43038 19966 43090 20018
rect 43710 19966 43762 20018
rect 8038 19854 8090 19906
rect 8318 19854 8370 19906
rect 24726 19854 24778 19906
rect 35982 19854 36034 19906
rect 37886 19854 37938 19906
rect 44046 19854 44098 19906
rect 22542 19742 22594 19794
rect 26014 19742 26066 19794
rect 27638 19742 27690 19794
rect 31726 19742 31778 19794
rect 41134 19742 41186 19794
rect 42030 19742 42082 19794
rect 42590 19742 42642 19794
rect 43374 19742 43426 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 9774 19406 9826 19458
rect 22224 19406 22276 19458
rect 26966 19406 27018 19458
rect 35870 19406 35922 19458
rect 13806 19294 13858 19346
rect 22822 19294 22874 19346
rect 29486 19350 29538 19402
rect 38558 19406 38610 19458
rect 39772 19406 39824 19458
rect 23494 19294 23546 19346
rect 35198 19294 35250 19346
rect 8542 19182 8594 19234
rect 9102 19154 9154 19206
rect 11678 19182 11730 19234
rect 12554 19182 12606 19234
rect 13470 19182 13522 19234
rect 14142 19182 14194 19234
rect 13806 19126 13858 19178
rect 14478 19182 14530 19234
rect 15038 19182 15090 19234
rect 15710 19182 15762 19234
rect 15374 19126 15426 19178
rect 21478 19182 21530 19234
rect 21982 19182 22034 19234
rect 23774 19182 23826 19234
rect 24558 19182 24610 19234
rect 27246 19182 27298 19234
rect 27470 19182 27522 19234
rect 27806 19182 27858 19234
rect 28030 19138 28082 19190
rect 29150 19182 29202 19234
rect 29486 19182 29538 19234
rect 34190 19182 34242 19234
rect 34862 19182 34914 19234
rect 35534 19182 35586 19234
rect 37158 19238 37210 19290
rect 43598 19294 43650 19346
rect 44214 19294 44266 19346
rect 37662 19182 37714 19234
rect 37904 19182 37956 19234
rect 38222 19182 38274 19234
rect 40014 19182 40066 19234
rect 40518 19238 40570 19290
rect 40910 19182 40962 19234
rect 41694 19182 41746 19234
rect 8374 19014 8426 19066
rect 12798 19070 12850 19122
rect 21310 19070 21362 19122
rect 15598 19014 15650 19066
rect 26462 19070 26514 19122
rect 36990 19070 37042 19122
rect 27918 19014 27970 19066
rect 40686 19070 40738 19122
rect 17110 18958 17162 19010
rect 28646 18958 28698 19010
rect 34022 18958 34074 19010
rect 34526 18958 34578 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 18398 18510 18450 18562
rect 8878 18425 8930 18477
rect 9886 18398 9938 18450
rect 10222 18413 10274 18465
rect 10446 18398 10498 18450
rect 11006 18442 11058 18494
rect 11230 18398 11282 18450
rect 12014 18398 12066 18450
rect 13918 18425 13970 18477
rect 14926 18454 14978 18506
rect 21758 18510 21810 18562
rect 14590 18398 14642 18450
rect 15262 18398 15314 18450
rect 16942 18398 16994 18450
rect 17484 18398 17536 18450
rect 17726 18398 17778 18450
rect 10110 18286 10162 18338
rect 10894 18286 10946 18338
rect 14926 18286 14978 18338
rect 18230 18342 18282 18394
rect 19070 18398 19122 18450
rect 19854 18398 19906 18450
rect 22206 18398 22258 18450
rect 7982 18174 8034 18226
rect 9718 18230 9770 18282
rect 18902 18286 18954 18338
rect 22374 18342 22426 18394
rect 22878 18398 22930 18450
rect 23998 18398 24050 18450
rect 23756 18286 23808 18338
rect 24502 18342 24554 18394
rect 24670 18398 24722 18450
rect 25118 18398 25170 18450
rect 25454 18398 25506 18450
rect 26574 18398 26626 18450
rect 27022 18398 27074 18450
rect 27806 18398 27858 18450
rect 28030 18437 28082 18489
rect 28478 18398 28530 18450
rect 28814 18398 28866 18450
rect 29150 18413 29202 18465
rect 30046 18398 30098 18450
rect 30270 18398 30322 18450
rect 31390 18398 31442 18450
rect 32062 18398 32114 18450
rect 33518 18398 33570 18450
rect 34302 18398 34354 18450
rect 36206 18398 36258 18450
rect 39454 18398 39506 18450
rect 39790 18398 39842 18450
rect 40126 18398 40178 18450
rect 40798 18398 40850 18450
rect 41582 18398 41634 18450
rect 43486 18398 43538 18450
rect 44214 18398 44266 18450
rect 26798 18286 26850 18338
rect 28254 18286 28306 18338
rect 29262 18286 29314 18338
rect 36766 18286 36818 18338
rect 38670 18286 38722 18338
rect 16606 18174 16658 18226
rect 23120 18174 23172 18226
rect 30550 18174 30602 18226
rect 32398 18174 32450 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 12686 17838 12738 17890
rect 14590 17838 14642 17890
rect 19070 17838 19122 17890
rect 8318 17726 8370 17778
rect 10222 17726 10274 17778
rect 21870 17726 21922 17778
rect 23662 17782 23714 17834
rect 24446 17782 24498 17834
rect 28366 17838 28418 17890
rect 29878 17838 29930 17890
rect 30662 17838 30714 17890
rect 34060 17838 34112 17890
rect 25342 17726 25394 17778
rect 27582 17726 27634 17778
rect 31838 17782 31890 17834
rect 32286 17782 32338 17834
rect 37214 17838 37266 17890
rect 7534 17614 7586 17666
rect 11566 17614 11618 17666
rect 13470 17614 13522 17666
rect 14346 17614 14398 17666
rect 15822 17614 15874 17666
rect 16606 17614 16658 17666
rect 18510 17614 18562 17666
rect 12442 17558 12494 17610
rect 19406 17614 19458 17666
rect 20862 17614 20914 17666
rect 21534 17614 21586 17666
rect 22206 17614 22258 17666
rect 23774 17614 23826 17666
rect 24110 17614 24162 17666
rect 24558 17614 24610 17666
rect 24894 17614 24946 17666
rect 25454 17614 25506 17666
rect 26126 17614 26178 17666
rect 27246 17614 27298 17666
rect 27918 17614 27970 17666
rect 28702 17614 28754 17666
rect 21926 17558 21978 17610
rect 27470 17558 27522 17610
rect 29374 17614 29426 17666
rect 29598 17614 29650 17666
rect 30158 17614 30210 17666
rect 30382 17614 30434 17666
rect 31390 17614 31442 17666
rect 31726 17614 31778 17666
rect 32174 17614 32226 17666
rect 32510 17614 32562 17666
rect 32846 17614 32898 17666
rect 34302 17614 34354 17666
rect 34806 17670 34858 17722
rect 40126 17726 40178 17778
rect 42030 17726 42082 17778
rect 34974 17614 35026 17666
rect 35422 17614 35474 17666
rect 35590 17670 35642 17722
rect 36094 17614 36146 17666
rect 36336 17614 36388 17666
rect 36878 17614 36930 17666
rect 39342 17614 39394 17666
rect 42814 17614 42866 17666
rect 43318 17670 43370 17722
rect 43934 17726 43986 17778
rect 44270 17614 44322 17666
rect 42572 17502 42624 17554
rect 20526 17390 20578 17442
rect 43150 17446 43202 17498
rect 33182 17390 33234 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 8262 17054 8314 17106
rect 8934 17054 8986 17106
rect 16102 17054 16154 17106
rect 16606 17054 16658 17106
rect 34806 17054 34858 17106
rect 35198 17054 35250 17106
rect 35982 17054 36034 17106
rect 40126 17054 40178 17106
rect 41078 17054 41130 17106
rect 42926 17054 42978 17106
rect 43542 17054 43594 17106
rect 43934 17054 43986 17106
rect 18398 16942 18450 16994
rect 8430 16830 8482 16882
rect 9102 16830 9154 16882
rect 9438 16830 9490 16882
rect 12126 16830 12178 16882
rect 12686 16857 12738 16909
rect 16942 16830 16994 16882
rect 17484 16830 17536 16882
rect 18230 16886 18282 16938
rect 22430 16942 22482 16994
rect 41452 16942 41504 16994
rect 17726 16830 17778 16882
rect 19742 16830 19794 16882
rect 20526 16830 20578 16882
rect 23438 16830 23490 16882
rect 23756 16830 23808 16882
rect 24502 16886 24554 16938
rect 23998 16830 24050 16882
rect 24670 16830 24722 16882
rect 25790 16830 25842 16882
rect 26014 16830 26066 16882
rect 26910 16830 26962 16882
rect 27246 16830 27298 16882
rect 27467 16869 27519 16921
rect 29822 16886 29874 16938
rect 42366 16942 42418 16994
rect 28478 16830 28530 16882
rect 29486 16830 29538 16882
rect 30158 16830 30210 16882
rect 30494 16830 30546 16882
rect 30830 16830 30882 16882
rect 31614 16830 31666 16882
rect 31838 16869 31890 16921
rect 32286 16830 32338 16882
rect 35534 16830 35586 16882
rect 35646 16830 35698 16882
rect 39678 16830 39730 16882
rect 39790 16830 39842 16882
rect 42198 16886 42250 16938
rect 41694 16830 41746 16882
rect 42590 16830 42642 16882
rect 44270 16830 44322 16882
rect 10222 16718 10274 16770
rect 25902 16718 25954 16770
rect 27806 16718 27858 16770
rect 29934 16718 29986 16770
rect 31950 16718 32002 16770
rect 13582 16606 13634 16658
rect 30830 16662 30882 16714
rect 23102 16606 23154 16658
rect 39342 16606 39394 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 12798 16270 12850 16322
rect 26294 16270 26346 16322
rect 27022 16214 27074 16266
rect 28534 16270 28586 16322
rect 16158 16158 16210 16210
rect 23662 16158 23714 16210
rect 25566 16158 25618 16210
rect 31502 16214 31554 16266
rect 31950 16270 32002 16322
rect 33742 16270 33794 16322
rect 37662 16270 37714 16322
rect 29598 16158 29650 16210
rect 29934 16158 29986 16210
rect 40294 16158 40346 16210
rect 43542 16158 43594 16210
rect 44214 16158 44266 16210
rect 7870 16046 7922 16098
rect 8654 16046 8706 16098
rect 11454 16046 11506 16098
rect 11678 16046 11730 16098
rect 13470 16046 13522 16098
rect 14346 16046 14398 16098
rect 15374 16046 15426 16098
rect 12554 15990 12606 16042
rect 18062 16046 18114 16098
rect 19854 16046 19906 16098
rect 22878 16046 22930 16098
rect 26574 16046 26626 16098
rect 26798 16046 26850 16098
rect 27134 16046 27186 16098
rect 27470 16046 27522 16098
rect 27694 16046 27746 16098
rect 28366 16046 28418 16098
rect 29150 16046 29202 16098
rect 29486 16002 29538 16054
rect 30046 16031 30098 16083
rect 30270 16046 30322 16098
rect 31054 16046 31106 16098
rect 31390 16046 31442 16098
rect 32286 16046 32338 16098
rect 34078 16046 34130 16098
rect 34190 16046 34242 16098
rect 35646 16046 35698 16098
rect 37326 16046 37378 16098
rect 38446 16046 38498 16098
rect 10558 15934 10610 15986
rect 14590 15934 14642 15986
rect 34526 15934 34578 15986
rect 38950 15990 39002 16042
rect 38204 15934 38256 15986
rect 39118 15934 39170 15986
rect 39846 15934 39898 15986
rect 11118 15822 11170 15874
rect 19518 15822 19570 15874
rect 28030 15822 28082 15874
rect 32678 15822 32730 15874
rect 35310 15822 35362 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 7366 15486 7418 15538
rect 11566 15486 11618 15538
rect 24278 15486 24330 15538
rect 25398 15486 25450 15538
rect 43654 15486 43706 15538
rect 23774 15374 23826 15426
rect 7534 15262 7586 15314
rect 7870 15262 7922 15314
rect 8094 15277 8146 15329
rect 8654 15262 8706 15314
rect 8878 15306 8930 15358
rect 10222 15289 10274 15341
rect 12910 15262 12962 15314
rect 13246 15262 13298 15314
rect 13694 15301 13746 15353
rect 13918 15262 13970 15314
rect 14254 15262 14306 15314
rect 14814 15262 14866 15314
rect 8206 15150 8258 15202
rect 8990 15150 9042 15202
rect 13582 15150 13634 15202
rect 14982 15206 15034 15258
rect 15486 15262 15538 15314
rect 16942 15262 16994 15314
rect 17484 15262 17536 15314
rect 18230 15318 18282 15370
rect 29486 15374 29538 15426
rect 32006 15374 32058 15426
rect 17726 15262 17778 15314
rect 18398 15262 18450 15314
rect 19182 15262 19234 15314
rect 21758 15262 21810 15314
rect 22542 15262 22594 15314
rect 22860 15262 22912 15314
rect 23102 15262 23154 15314
rect 18846 15150 18898 15202
rect 19574 15150 19626 15202
rect 21422 15150 21474 15202
rect 23606 15206 23658 15258
rect 26126 15262 26178 15314
rect 26798 15262 26850 15314
rect 30494 15318 30546 15370
rect 39902 15374 39954 15426
rect 41470 15374 41522 15426
rect 30158 15262 30210 15314
rect 30718 15262 30770 15314
rect 31054 15262 31106 15314
rect 32958 15262 33010 15314
rect 34862 15262 34914 15314
rect 35198 15262 35250 15314
rect 36766 15262 36818 15314
rect 37102 15262 37154 15314
rect 37214 15262 37266 15314
rect 41638 15262 41690 15314
rect 42142 15262 42194 15314
rect 42702 15262 42754 15314
rect 26462 15150 26514 15202
rect 27582 15150 27634 15202
rect 30606 15150 30658 15202
rect 31390 15150 31442 15202
rect 33294 15150 33346 15202
rect 36374 15150 36426 15202
rect 37998 15150 38050 15202
rect 43038 15150 43090 15202
rect 12742 15038 12794 15090
rect 15728 15038 15780 15090
rect 16606 15038 16658 15090
rect 22206 15038 22258 15090
rect 34526 15038 34578 15090
rect 35534 15038 35586 15090
rect 42384 15038 42436 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 11454 14702 11506 14754
rect 14590 14702 14642 14754
rect 19276 14702 19328 14754
rect 28384 14702 28436 14754
rect 34956 14702 35008 14754
rect 38782 14702 38834 14754
rect 8766 14590 8818 14642
rect 16830 14590 16882 14642
rect 18734 14590 18786 14642
rect 7758 14478 7810 14530
rect 8430 14478 8482 14530
rect 8654 14434 8706 14486
rect 8990 14478 9042 14530
rect 10110 14450 10162 14502
rect 13470 14478 13522 14530
rect 15598 14478 15650 14530
rect 14346 14422 14398 14474
rect 15934 14478 15986 14530
rect 16046 14478 16098 14530
rect 19518 14478 19570 14530
rect 20022 14422 20074 14474
rect 21422 14450 21474 14502
rect 24446 14478 24498 14530
rect 25118 14478 25170 14530
rect 24950 14422 25002 14474
rect 27246 14478 27298 14530
rect 27470 14478 27522 14530
rect 27638 14534 27690 14586
rect 31334 14590 31386 14642
rect 41582 14590 41634 14642
rect 28142 14478 28194 14530
rect 29486 14478 29538 14530
rect 30942 14478 30994 14530
rect 24204 14366 24256 14418
rect 19854 14310 19906 14362
rect 29990 14422 30042 14474
rect 34190 14478 34242 14530
rect 35198 14478 35250 14530
rect 36374 14478 36426 14530
rect 29244 14366 29296 14418
rect 35702 14422 35754 14474
rect 37662 14478 37714 14530
rect 30606 14366 30658 14418
rect 7926 14254 7978 14306
rect 22654 14254 22706 14306
rect 26518 14254 26570 14306
rect 29822 14310 29874 14362
rect 35870 14366 35922 14418
rect 37158 14422 37210 14474
rect 38446 14478 38498 14530
rect 40798 14478 40850 14530
rect 36990 14366 37042 14418
rect 37904 14366 37956 14418
rect 43486 14366 43538 14418
rect 26910 14254 26962 14306
rect 33854 14254 33906 14306
rect 44102 14254 44154 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 41190 13918 41242 13970
rect 9662 13806 9714 13858
rect 16494 13862 16546 13914
rect 14254 13806 14306 13858
rect 19966 13806 20018 13858
rect 21310 13806 21362 13858
rect 30382 13806 30434 13858
rect 41470 13806 41522 13858
rect 43486 13862 43538 13914
rect 42384 13806 42436 13858
rect 7534 13694 7586 13746
rect 7758 13694 7810 13746
rect 8094 13709 8146 13761
rect 8542 13694 8594 13746
rect 8878 13738 8930 13790
rect 11566 13694 11618 13746
rect 12350 13694 12402 13746
rect 13134 13694 13186 13746
rect 14010 13694 14062 13746
rect 15598 13694 15650 13746
rect 15916 13694 15968 13746
rect 16158 13694 16210 13746
rect 16662 13638 16714 13690
rect 17278 13694 17330 13746
rect 18062 13694 18114 13746
rect 23998 13694 24050 13746
rect 24110 13694 24162 13746
rect 27694 13694 27746 13746
rect 32062 13694 32114 13746
rect 33070 13694 33122 13746
rect 36094 13694 36146 13746
rect 36878 13694 36930 13746
rect 39118 13694 39170 13746
rect 40462 13694 40514 13746
rect 8206 13582 8258 13634
rect 8990 13582 9042 13634
rect 41638 13638 41690 13690
rect 42142 13694 42194 13746
rect 42908 13694 42960 13746
rect 43150 13694 43202 13746
rect 23214 13582 23266 13634
rect 24446 13582 24498 13634
rect 28478 13582 28530 13634
rect 33854 13582 33906 13634
rect 35758 13582 35810 13634
rect 38782 13582 38834 13634
rect 43654 13638 43706 13690
rect 7366 13470 7418 13522
rect 15262 13470 15314 13522
rect 31726 13470 31778 13522
rect 39454 13470 39506 13522
rect 40126 13470 40178 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 29374 13134 29426 13186
rect 30606 13134 30658 13186
rect 32044 13134 32096 13186
rect 9774 13022 9826 13074
rect 11678 13022 11730 13074
rect 14478 13022 14530 13074
rect 16382 13022 16434 13074
rect 18230 13022 18282 13074
rect 21982 13022 22034 13074
rect 33462 13022 33514 13074
rect 39006 13022 39058 13074
rect 41358 13022 41410 13074
rect 8990 12910 9042 12962
rect 17166 12910 17218 12962
rect 17278 12910 17330 12962
rect 20302 12910 20354 12962
rect 21198 12910 21250 12962
rect 25678 12910 25730 12962
rect 27358 12910 27410 12962
rect 23886 12798 23938 12850
rect 26854 12854 26906 12906
rect 29038 12910 29090 12962
rect 30270 12910 30322 12962
rect 31502 12910 31554 12962
rect 32286 12910 32338 12962
rect 32958 12910 33010 12962
rect 26686 12798 26738 12850
rect 32790 12854 32842 12906
rect 34190 12910 34242 12962
rect 34358 12910 34410 12962
rect 34862 12910 34914 12962
rect 35758 12910 35810 12962
rect 39790 12910 39842 12962
rect 40574 12910 40626 12962
rect 43598 12910 43650 12962
rect 27600 12798 27652 12850
rect 35104 12798 35156 12850
rect 37102 12798 37154 12850
rect 43262 12798 43314 12850
rect 17614 12686 17666 12738
rect 19966 12686 20018 12738
rect 25342 12686 25394 12738
rect 26406 12686 26458 12738
rect 31166 12686 31218 12738
rect 35590 12686 35642 12738
rect 36150 12686 36202 12738
rect 43934 12686 43986 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 28870 12350 28922 12402
rect 36430 12350 36482 12402
rect 12126 12238 12178 12290
rect 13694 12238 13746 12290
rect 13450 12182 13502 12234
rect 14254 12238 14306 12290
rect 25230 12238 25282 12290
rect 26574 12238 26626 12290
rect 43598 12238 43650 12290
rect 9438 12126 9490 12178
rect 10222 12126 10274 12178
rect 12574 12126 12626 12178
rect 16158 12126 16210 12178
rect 16942 12126 16994 12178
rect 18398 12126 18450 12178
rect 18734 12141 18786 12193
rect 19406 12153 19458 12205
rect 21422 12126 21474 12178
rect 21870 12126 21922 12178
rect 25398 12070 25450 12122
rect 25902 12126 25954 12178
rect 18846 12014 18898 12066
rect 22654 12014 22706 12066
rect 24558 12014 24610 12066
rect 26742 12070 26794 12122
rect 27246 12126 27298 12178
rect 27806 12126 27858 12178
rect 29710 12126 29762 12178
rect 30494 12126 30546 12178
rect 33630 12153 33682 12205
rect 35086 12126 35138 12178
rect 36094 12126 36146 12178
rect 37326 12153 37378 12205
rect 40910 12126 40962 12178
rect 41694 12126 41746 12178
rect 32398 12014 32450 12066
rect 44214 12014 44266 12066
rect 26144 11902 26196 11954
rect 27488 11902 27540 11954
rect 28142 11902 28194 11954
rect 39006 11902 39058 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 11342 11566 11394 11618
rect 22318 11566 22370 11618
rect 43934 11566 43986 11618
rect 18734 11454 18786 11506
rect 20638 11454 20690 11506
rect 24670 11454 24722 11506
rect 26014 11454 26066 11506
rect 27918 11454 27970 11506
rect 34526 11454 34578 11506
rect 35870 11454 35922 11506
rect 39902 11454 39954 11506
rect 12014 11314 12066 11366
rect 17950 11342 18002 11394
rect 21646 11314 21698 11366
rect 24334 11342 24386 11394
rect 24894 11342 24946 11394
rect 28702 11342 28754 11394
rect 24558 11286 24610 11338
rect 29038 11342 29090 11394
rect 29822 11342 29874 11394
rect 32286 11298 32338 11350
rect 32510 11342 32562 11394
rect 35534 11314 35586 11366
rect 35982 11327 36034 11379
rect 36206 11342 36258 11394
rect 37214 11342 37266 11394
rect 39230 11314 39282 11366
rect 40145 11342 40197 11394
rect 41022 11342 41074 11394
rect 41713 11342 41765 11394
rect 42590 11342 42642 11394
rect 42814 11342 42866 11394
rect 43542 11342 43594 11394
rect 44270 11342 44322 11394
rect 31726 11230 31778 11282
rect 41470 11230 41522 11282
rect 32510 11174 32562 11226
rect 17110 11118 17162 11170
rect 42982 11118 43034 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 24446 10782 24498 10834
rect 23886 10670 23938 10722
rect 14030 10558 14082 10610
rect 16718 10558 16770 10610
rect 17502 10573 17554 10625
rect 17838 10558 17890 10610
rect 18958 10558 19010 10610
rect 23642 10614 23694 10666
rect 25342 10670 25394 10722
rect 21982 10558 22034 10610
rect 22430 10558 22482 10610
rect 22766 10558 22818 10610
rect 24782 10558 24834 10610
rect 28030 10558 28082 10610
rect 28142 10558 28194 10610
rect 31838 10585 31890 10637
rect 33946 10614 33998 10666
rect 32622 10558 32674 10610
rect 33070 10558 33122 10610
rect 34918 10614 34970 10666
rect 34190 10558 34242 10610
rect 34638 10558 34690 10610
rect 35422 10558 35474 10610
rect 38782 10558 38834 10610
rect 39118 10558 39170 10610
rect 39342 10597 39394 10649
rect 41489 10614 41541 10666
rect 39678 10558 39730 10610
rect 40014 10558 40066 10610
rect 41246 10558 41298 10610
rect 43057 10614 43109 10666
rect 42366 10558 42418 10610
rect 43934 10558 43986 10610
rect 14814 10446 14866 10498
rect 17390 10446 17442 10498
rect 19294 10446 19346 10498
rect 21198 10446 21250 10498
rect 27246 10446 27298 10498
rect 28478 10446 28530 10498
rect 35086 10446 35138 10498
rect 36206 10446 36258 10498
rect 38110 10446 38162 10498
rect 39566 10446 39618 10498
rect 18622 10334 18674 10386
rect 22262 10390 22314 10442
rect 30942 10334 30994 10386
rect 32454 10334 32506 10386
rect 40182 10334 40234 10386
rect 42814 10334 42866 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 22318 9998 22370 10050
rect 30270 9998 30322 10050
rect 31446 9942 31498 9994
rect 36318 9998 36370 10050
rect 16942 9886 16994 9938
rect 19742 9886 19794 9938
rect 32510 9886 32562 9938
rect 34414 9886 34466 9938
rect 17950 9746 18002 9798
rect 20414 9746 20466 9798
rect 21310 9746 21362 9798
rect 24110 9774 24162 9826
rect 24986 9774 25038 9826
rect 26238 9774 26290 9826
rect 27114 9774 27166 9826
rect 30606 9774 30658 9826
rect 25230 9662 25282 9714
rect 27358 9662 27410 9714
rect 31614 9718 31666 9770
rect 31726 9774 31778 9826
rect 35198 9774 35250 9826
rect 36878 9774 36930 9826
rect 37662 9774 37714 9826
rect 39566 9774 39618 9826
rect 36074 9718 36126 9770
rect 39902 9774 39954 9826
rect 40686 9774 40738 9826
rect 42926 9774 42978 9826
rect 44270 9774 44322 9826
rect 42590 9662 42642 9714
rect 43094 9550 43146 9602
rect 43934 9550 43986 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 16774 9214 16826 9266
rect 23326 9214 23378 9266
rect 25566 9158 25618 9210
rect 37998 9214 38050 9266
rect 39566 9158 39618 9210
rect 16494 8990 16546 9042
rect 16942 8990 16994 9042
rect 17950 8990 18002 9042
rect 18342 9019 18394 9071
rect 18622 8990 18674 9042
rect 18846 8990 18898 9042
rect 21982 9017 22034 9069
rect 25342 8990 25394 9042
rect 25566 9017 25618 9069
rect 25902 8990 25954 9042
rect 29150 8990 29202 9042
rect 29486 8990 29538 9042
rect 31950 8990 32002 9042
rect 33518 8990 33570 9042
rect 34302 8990 34354 9042
rect 36654 9017 36706 9069
rect 39734 9046 39786 9098
rect 39454 8990 39506 9042
rect 40126 8990 40178 9042
rect 43710 8990 43762 9042
rect 43822 9010 43874 9062
rect 18174 8878 18226 8930
rect 19630 8878 19682 8930
rect 21534 8878 21586 8930
rect 36206 8878 36258 8930
rect 41022 8878 41074 8930
rect 42926 8878 42978 8930
rect 16326 8822 16378 8874
rect 17782 8766 17834 8818
rect 28814 8766 28866 8818
rect 29822 8766 29874 8818
rect 32286 8766 32338 8818
rect 43990 8766 44042 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 17278 8318 17330 8370
rect 20078 8318 20130 8370
rect 25230 8318 25282 8370
rect 31166 8318 31218 8370
rect 34078 8318 34130 8370
rect 36374 8318 36426 8370
rect 16494 8206 16546 8258
rect 19742 8206 19794 8258
rect 19910 8176 19962 8228
rect 20302 8206 20354 8258
rect 23774 8178 23826 8230
rect 24110 8206 24162 8258
rect 24986 8206 25038 8258
rect 26014 8206 26066 8258
rect 26686 8206 26738 8258
rect 19182 8094 19234 8146
rect 26518 8150 26570 8202
rect 29262 8206 29314 8258
rect 31950 8206 32002 8258
rect 34414 8150 34466 8202
rect 34638 8206 34690 8258
rect 35514 8206 35566 8258
rect 37214 8206 37266 8258
rect 37550 8178 37602 8230
rect 39790 8206 39842 8258
rect 40350 8178 40402 8230
rect 43934 8206 43986 8258
rect 25772 8094 25824 8146
rect 35758 8094 35810 8146
rect 20638 7982 20690 8034
rect 22094 7982 22146 8034
rect 27190 7982 27242 8034
rect 27638 7982 27690 8034
rect 37046 7982 37098 8034
rect 41694 7982 41746 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 16774 7646 16826 7698
rect 28646 7646 28698 7698
rect 18734 7590 18786 7642
rect 23438 7534 23490 7586
rect 16942 7422 16994 7474
rect 17502 7466 17554 7518
rect 17838 7422 17890 7474
rect 18510 7437 18562 7489
rect 18846 7422 18898 7474
rect 19070 7422 19122 7474
rect 23194 7478 23246 7530
rect 25566 7534 25618 7586
rect 29132 7534 29184 7586
rect 30046 7534 30098 7586
rect 22318 7422 22370 7474
rect 25734 7366 25786 7418
rect 26238 7422 26290 7474
rect 26910 7422 26962 7474
rect 27246 7449 27298 7501
rect 27582 7422 27634 7474
rect 27918 7422 27970 7474
rect 29878 7478 29930 7530
rect 29374 7422 29426 7474
rect 30270 7422 30322 7474
rect 35758 7422 35810 7474
rect 36094 7466 36146 7518
rect 36430 7422 36482 7474
rect 36990 7422 37042 7474
rect 37718 7478 37770 7530
rect 38689 7478 38741 7530
rect 37326 7422 37378 7474
rect 37998 7422 38050 7474
rect 39566 7422 39618 7474
rect 40014 7466 40066 7518
rect 40350 7422 40402 7474
rect 40910 7449 40962 7501
rect 42254 7422 42306 7474
rect 43822 7437 43874 7489
rect 44046 7422 44098 7474
rect 17390 7310 17442 7362
rect 19854 7310 19906 7362
rect 21758 7310 21810 7362
rect 27022 7310 27074 7362
rect 35982 7310 36034 7362
rect 37662 7310 37714 7362
rect 38446 7310 38498 7362
rect 39902 7310 39954 7362
rect 43710 7310 43762 7362
rect 26480 7198 26532 7250
rect 30606 7198 30658 7250
rect 35422 7198 35474 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 22318 6862 22370 6914
rect 28366 6862 28418 6914
rect 24222 6750 24274 6802
rect 37102 6750 37154 6802
rect 43262 6750 43314 6802
rect 15822 6638 15874 6690
rect 16606 6638 16658 6690
rect 18958 6638 19010 6690
rect 19518 6638 19570 6690
rect 20638 6638 20690 6690
rect 20394 6582 20446 6634
rect 21646 6610 21698 6662
rect 24110 6638 24162 6690
rect 24446 6611 24498 6663
rect 24782 6638 24834 6690
rect 25118 6638 25170 6690
rect 26910 6638 26962 6690
rect 18510 6526 18562 6578
rect 26033 6582 26085 6634
rect 27246 6638 27298 6690
rect 28122 6638 28174 6690
rect 29486 6638 29538 6690
rect 29654 6638 29706 6690
rect 30158 6638 30210 6690
rect 30400 6638 30452 6690
rect 30718 6638 30770 6690
rect 34078 6638 34130 6690
rect 35758 6638 35810 6690
rect 36990 6638 37042 6690
rect 37662 6638 37714 6690
rect 25790 6526 25842 6578
rect 34582 6582 34634 6634
rect 33836 6526 33888 6578
rect 34750 6526 34802 6578
rect 35254 6582 35306 6634
rect 35086 6526 35138 6578
rect 37326 6582 37378 6634
rect 38782 6610 38834 6662
rect 44046 6638 44098 6690
rect 36000 6526 36052 6578
rect 41358 6526 41410 6578
rect 19126 6414 19178 6466
rect 31054 6414 31106 6466
rect 31670 6414 31722 6466
rect 40126 6414 40178 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 16326 6078 16378 6130
rect 24558 5966 24610 6018
rect 26462 5966 26514 6018
rect 28814 5966 28866 6018
rect 29374 5966 29426 6018
rect 33742 5966 33794 6018
rect 37326 6022 37378 6074
rect 35422 5966 35474 6018
rect 16494 5854 16546 5906
rect 16942 5854 16994 5906
rect 17502 5869 17554 5921
rect 17726 5854 17778 5906
rect 18286 5854 18338 5906
rect 18510 5898 18562 5950
rect 18958 5854 19010 5906
rect 19294 5898 19346 5950
rect 19630 5854 19682 5906
rect 23214 5854 23266 5906
rect 23438 5854 23490 5906
rect 24314 5854 24366 5906
rect 25342 5854 25394 5906
rect 26218 5854 26270 5906
rect 26798 5854 26850 5906
rect 27694 5854 27746 5906
rect 28570 5854 28622 5906
rect 31278 5854 31330 5906
rect 32062 5854 32114 5906
rect 33910 5854 33962 5906
rect 34414 5854 34466 5906
rect 35665 5854 35717 5906
rect 36542 5854 36594 5906
rect 37102 5898 37154 5950
rect 37438 5854 37490 5906
rect 40238 5881 40290 5933
rect 40910 5854 40962 5906
rect 41246 5869 41298 5921
rect 41694 5881 41746 5933
rect 17390 5742 17442 5794
rect 18622 5742 18674 5794
rect 19406 5742 19458 5794
rect 20414 5742 20466 5794
rect 22318 5742 22370 5794
rect 39342 5742 39394 5794
rect 41358 5742 41410 5794
rect 42702 5742 42754 5794
rect 16774 5630 16826 5682
rect 22878 5630 22930 5682
rect 27134 5630 27186 5682
rect 34656 5630 34708 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 43934 5294 43986 5346
rect 15150 5182 15202 5234
rect 17054 5182 17106 5234
rect 20638 5182 20690 5234
rect 22542 5182 22594 5234
rect 24446 5182 24498 5234
rect 25006 5182 25058 5234
rect 26910 5182 26962 5234
rect 29598 5182 29650 5234
rect 31502 5182 31554 5234
rect 35646 5182 35698 5234
rect 39566 5182 39618 5234
rect 43486 5182 43538 5234
rect 17838 5070 17890 5122
rect 17950 5070 18002 5122
rect 18734 5070 18786 5122
rect 21534 5070 21586 5122
rect 21758 5070 21810 5122
rect 27694 5070 27746 5122
rect 28030 5070 28082 5122
rect 28366 5070 28418 5122
rect 32286 5070 32338 5122
rect 32958 5070 33010 5122
rect 33742 5070 33794 5122
rect 35982 5070 36034 5122
rect 36318 5070 36370 5122
rect 36878 5070 36930 5122
rect 37662 5070 37714 5122
rect 39902 5070 39954 5122
rect 40686 5070 40738 5122
rect 43038 5070 43090 5122
rect 43318 5040 43370 5092
rect 44270 5070 44322 5122
rect 42590 4958 42642 5010
rect 21366 4846 21418 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 38502 4510 38554 4562
rect 28702 4398 28754 4450
rect 29598 4398 29650 4450
rect 30512 4398 30564 4450
rect 17614 4286 17666 4338
rect 17950 4301 18002 4353
rect 18286 4286 18338 4338
rect 22206 4286 22258 4338
rect 22542 4301 22594 4353
rect 29766 4342 29818 4394
rect 36094 4398 36146 4450
rect 36990 4398 37042 4450
rect 39230 4398 39282 4450
rect 22878 4286 22930 4338
rect 26014 4286 26066 4338
rect 26798 4286 26850 4338
rect 30270 4286 30322 4338
rect 37233 4342 37285 4394
rect 33406 4286 33458 4338
rect 39473 4342 39525 4394
rect 38110 4286 38162 4338
rect 38334 4286 38386 4338
rect 40350 4286 40402 4338
rect 44046 4286 44098 4338
rect 18062 4174 18114 4226
rect 19518 4174 19570 4226
rect 21422 4174 21474 4226
rect 22430 4174 22482 4226
rect 34190 4174 34242 4226
rect 41358 4174 41410 4226
rect 43262 4174 43314 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 17334 3726 17386 3778
rect 25566 3726 25618 3778
rect 29280 3726 29332 3778
rect 32286 3726 32338 3778
rect 33406 3726 33458 3778
rect 34638 3726 34690 3778
rect 36766 3726 36818 3778
rect 27862 3614 27914 3666
rect 42870 3670 42922 3722
rect 17502 3502 17554 3554
rect 18174 3502 18226 3554
rect 19854 3474 19906 3526
rect 21086 3474 21138 3526
rect 22990 3502 23042 3554
rect 24558 3474 24610 3526
rect 28366 3502 28418 3554
rect 28534 3558 28586 3610
rect 38502 3614 38554 3666
rect 38782 3614 38834 3666
rect 39902 3614 39954 3666
rect 41806 3614 41858 3666
rect 43598 3614 43650 3666
rect 29038 3502 29090 3554
rect 34302 3502 34354 3554
rect 36430 3502 36482 3554
rect 38894 3487 38946 3539
rect 39118 3502 39170 3554
rect 42590 3502 42642 3554
rect 42702 3446 42754 3498
rect 43710 3487 43762 3539
rect 43934 3502 43986 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 41692 43092 41748 43102
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 41692 42194 41748 43036
rect 41692 42142 41694 42194
rect 41746 42142 41748 42194
rect 41692 42130 41748 42142
rect 32844 42028 33236 42084
rect 32284 42008 32340 42020
rect 31276 41985 31332 41997
rect 31276 41933 31278 41985
rect 31330 41933 31332 41985
rect 31164 41860 31220 41870
rect 30492 41858 31220 41860
rect 30492 41806 31166 41858
rect 31218 41806 31220 41858
rect 30492 41804 31220 41806
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 22540 41356 23044 41412
rect 22540 41186 22596 41356
rect 22988 41298 23044 41356
rect 22988 41246 22990 41298
rect 23042 41246 23044 41298
rect 22540 41134 22542 41186
rect 22594 41134 22596 41186
rect 22540 41122 22596 41134
rect 22652 41186 22708 41198
rect 22652 41134 22654 41186
rect 22706 41134 22708 41186
rect 22260 41076 22316 41086
rect 21868 41074 22316 41076
rect 21868 41022 22262 41074
rect 22314 41022 22316 41074
rect 21868 41020 22316 41022
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 21868 40628 21924 41020
rect 22260 41010 22316 41020
rect 21756 40572 21924 40628
rect 20748 40402 20804 40414
rect 20748 40350 20750 40402
rect 20802 40350 20804 40402
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 20748 39620 20804 40350
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19740 38836 19796 38846
rect 19628 38780 19740 38836
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 19628 37266 19684 38780
rect 19740 38742 19796 38780
rect 20748 38836 20804 39564
rect 21532 40290 21588 40302
rect 21532 40238 21534 40290
rect 21586 40238 21588 40290
rect 21532 39172 21588 40238
rect 21756 40068 21812 40572
rect 21756 40012 22036 40068
rect 21532 39106 21588 39116
rect 21868 39786 21924 39798
rect 21868 39734 21870 39786
rect 21922 39734 21924 39786
rect 20748 38770 20804 38780
rect 20188 38724 20244 38734
rect 20524 38722 20580 38734
rect 20524 38670 20526 38722
rect 20578 38670 20580 38722
rect 20524 38668 20580 38670
rect 20188 37940 20244 38668
rect 20300 38612 20580 38668
rect 21868 38724 21924 39734
rect 21980 39618 22036 40012
rect 22652 39732 22708 41134
rect 22428 39676 22708 39732
rect 21980 39566 21982 39618
rect 22034 39566 22036 39618
rect 21980 39554 22036 39566
rect 22316 39618 22372 39630
rect 22316 39566 22318 39618
rect 22370 39566 22372 39618
rect 21868 38658 21924 38668
rect 20300 38162 20356 38612
rect 20300 38110 20302 38162
rect 20354 38110 20356 38162
rect 20300 38098 20356 38110
rect 21868 38218 21924 38230
rect 21868 38166 21870 38218
rect 21922 38166 21924 38218
rect 20748 38052 20804 38062
rect 20412 38006 20468 38018
rect 20412 37954 20414 38006
rect 20466 37954 20468 38006
rect 20748 37958 20804 37996
rect 20412 37940 20468 37954
rect 20188 37884 20468 37940
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37214 19630 37266
rect 19682 37214 19684 37266
rect 19628 37202 19684 37214
rect 20188 37380 20244 37390
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 12124 36484 12180 36494
rect 12124 36482 12964 36484
rect 12124 36430 12126 36482
rect 12178 36430 12964 36482
rect 12124 36428 12964 36430
rect 12124 36418 12180 36428
rect 11788 36260 11844 36270
rect 11788 36258 11956 36260
rect 11788 36206 11790 36258
rect 11842 36206 11956 36258
rect 11788 36204 11956 36206
rect 11788 36194 11844 36204
rect 9548 35700 9604 35710
rect 8876 35698 9604 35700
rect 8876 35646 9550 35698
rect 9602 35646 9604 35698
rect 8876 35644 9604 35646
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 8764 33908 8820 33918
rect 8652 33906 8820 33908
rect 8652 33854 8766 33906
rect 8818 33854 8820 33906
rect 8652 33852 8820 33854
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 6076 33348 6132 33358
rect 6860 33348 6916 33358
rect 6076 33254 6132 33292
rect 6412 33346 6916 33348
rect 6412 33294 6862 33346
rect 6914 33294 6916 33346
rect 6412 33292 6916 33294
rect 6412 32674 6468 33292
rect 6860 33282 6916 33292
rect 8652 33348 8708 33852
rect 8764 33842 8820 33852
rect 8764 33460 8820 33470
rect 8876 33460 8932 35644
rect 9548 35634 9604 35644
rect 10424 35700 10480 35710
rect 10424 35606 10480 35644
rect 11116 35700 11172 35710
rect 10668 35474 10724 35486
rect 10668 35422 10670 35474
rect 10722 35422 10724 35474
rect 10332 35364 10388 35374
rect 9100 35140 9156 35150
rect 9100 34130 9156 35084
rect 10332 35026 10388 35308
rect 10332 34974 10334 35026
rect 10386 34974 10388 35026
rect 10332 34962 10388 34974
rect 9903 34132 9959 34142
rect 9100 34078 9102 34130
rect 9154 34078 9156 34130
rect 9100 34066 9156 34078
rect 9772 34130 9959 34132
rect 9772 34078 9905 34130
rect 9957 34078 9959 34130
rect 9772 34076 9959 34078
rect 8764 33458 8932 33460
rect 8764 33406 8766 33458
rect 8818 33406 8932 33458
rect 8764 33404 8932 33406
rect 9660 33906 9716 33918
rect 9660 33854 9662 33906
rect 9714 33854 9716 33906
rect 8764 33394 8820 33404
rect 8652 33282 8708 33292
rect 9100 33348 9156 33358
rect 6412 32622 6414 32674
rect 6466 32622 6468 32674
rect 6412 32610 6468 32622
rect 9100 32564 9156 33292
rect 9548 32564 9604 32574
rect 9100 32562 9604 32564
rect 9100 32510 9102 32562
rect 9154 32510 9550 32562
rect 9602 32510 9604 32562
rect 9100 32508 9604 32510
rect 9100 32498 9156 32508
rect 9548 32498 9604 32508
rect 9660 32564 9716 33854
rect 9772 33460 9828 34076
rect 9903 34066 9959 34076
rect 10668 34132 10724 35422
rect 11004 35252 11060 35262
rect 11004 34580 11060 35196
rect 11004 34514 11060 34524
rect 11116 34356 11172 35644
rect 11695 35698 11751 35710
rect 11695 35646 11697 35698
rect 11749 35646 11751 35698
rect 11452 35474 11508 35486
rect 11452 35422 11454 35474
rect 11506 35422 11508 35474
rect 11452 35252 11508 35422
rect 11695 35364 11751 35646
rect 11695 35298 11751 35308
rect 11900 35252 11956 36204
rect 12572 35700 12628 35738
rect 12572 35634 12628 35644
rect 11900 35196 12068 35252
rect 11452 35186 11508 35196
rect 12012 35140 12068 35196
rect 12012 35074 12068 35084
rect 12236 34916 12292 34926
rect 12012 34914 12292 34916
rect 12012 34862 12238 34914
rect 12290 34862 12292 34914
rect 12012 34860 12292 34862
rect 10668 34066 10724 34076
rect 10780 34300 11172 34356
rect 10780 34130 10836 34300
rect 10780 34078 10782 34130
rect 10834 34078 10836 34130
rect 10780 34066 10836 34078
rect 11004 34132 11060 34142
rect 11004 34038 11060 34076
rect 9772 33394 9828 33404
rect 9884 33908 9940 33918
rect 9884 33458 9940 33852
rect 11116 33796 11172 34300
rect 11788 34580 11844 34590
rect 11788 34130 11844 34524
rect 11788 34078 11790 34130
rect 11842 34078 11844 34130
rect 11788 34066 11844 34078
rect 11116 33730 11172 33740
rect 9884 33406 9886 33458
rect 9938 33406 9940 33458
rect 9884 33394 9940 33406
rect 11788 33460 11844 33470
rect 11788 33366 11844 33404
rect 12012 32900 12068 34860
rect 12236 34850 12292 34860
rect 12292 33796 12348 33806
rect 12292 33570 12348 33740
rect 12292 33518 12294 33570
rect 12346 33518 12348 33570
rect 12292 33506 12348 33518
rect 12908 33460 12964 36428
rect 15372 36260 15428 36270
rect 15148 36258 15428 36260
rect 15148 36206 15374 36258
rect 15426 36206 15428 36258
rect 15148 36204 15428 36206
rect 13132 35698 13188 35710
rect 13132 35646 13134 35698
rect 13186 35646 13188 35698
rect 13020 34914 13076 34926
rect 13020 34862 13022 34914
rect 13074 34862 13076 34914
rect 13020 34692 13076 34862
rect 13020 34132 13076 34636
rect 13020 34066 13076 34076
rect 13132 33684 13188 35646
rect 13916 35588 13972 35598
rect 13804 35586 13972 35588
rect 13804 35534 13918 35586
rect 13970 35534 13972 35586
rect 13804 35532 13972 35534
rect 13356 35140 13412 35150
rect 13356 34914 13412 35084
rect 13356 34862 13358 34914
rect 13410 34862 13412 34914
rect 13356 34850 13412 34862
rect 13692 34692 13748 34702
rect 13692 34598 13748 34636
rect 13692 34244 13748 34254
rect 13804 34244 13860 35532
rect 13916 35522 13972 35532
rect 15148 34914 15204 36204
rect 15372 36194 15428 36204
rect 16660 36258 16716 36270
rect 16660 36206 16662 36258
rect 16714 36206 16716 36258
rect 16660 35810 16716 36206
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 16660 35758 16662 35810
rect 16714 35758 16716 35810
rect 16660 35746 16716 35758
rect 20188 35810 20244 37324
rect 21532 37380 21588 37390
rect 20412 37154 20468 37166
rect 20412 37102 20414 37154
rect 20466 37102 20468 37154
rect 20300 36596 20356 36606
rect 20412 36596 20468 37102
rect 20636 37156 20692 37166
rect 20300 36594 20468 36596
rect 20300 36542 20302 36594
rect 20354 36542 20468 36594
rect 20300 36540 20468 36542
rect 20524 37044 20580 37054
rect 20300 36530 20356 36540
rect 20524 36484 20580 36988
rect 20412 36467 20580 36484
rect 20412 36415 20414 36467
rect 20466 36428 20580 36467
rect 20636 36482 20692 37100
rect 20636 36430 20638 36482
rect 20690 36430 20692 36482
rect 20466 36415 20468 36428
rect 20636 36418 20692 36430
rect 21420 36484 21476 36494
rect 21532 36484 21588 37324
rect 21420 36482 21588 36484
rect 21420 36430 21422 36482
rect 21474 36430 21588 36482
rect 21420 36428 21588 36430
rect 21644 37156 21700 37166
rect 21644 36482 21700 37100
rect 21868 37044 21924 38166
rect 21980 38050 22036 38062
rect 21980 37998 21982 38050
rect 22034 37998 22036 38050
rect 21980 37604 22036 37998
rect 22316 38050 22372 39566
rect 22428 38948 22484 39676
rect 22988 39620 23044 41246
rect 26460 41298 26516 41310
rect 26460 41246 26462 41298
rect 26514 41246 26516 41298
rect 23324 41188 23380 41198
rect 23212 41186 23380 41188
rect 23100 41142 23156 41154
rect 23100 41090 23102 41142
rect 23154 41090 23156 41142
rect 23100 40180 23156 41090
rect 23100 40114 23156 40124
rect 23212 41134 23326 41186
rect 23378 41134 23380 41186
rect 23212 41132 23380 41134
rect 23212 40404 23268 41132
rect 23324 41122 23380 41132
rect 24668 41188 24724 41198
rect 23940 40570 23996 40582
rect 23940 40518 23942 40570
rect 23994 40518 23996 40570
rect 22648 39580 23044 39620
rect 22648 39528 22650 39580
rect 22702 39564 23044 39580
rect 23100 39786 23156 39798
rect 23100 39734 23102 39786
rect 23154 39734 23156 39786
rect 22702 39528 22704 39564
rect 22648 39508 22704 39528
rect 22648 39442 22704 39452
rect 23100 39396 23156 39734
rect 22820 39340 23156 39396
rect 22428 38946 22708 38948
rect 22428 38894 22430 38946
rect 22482 38894 22708 38946
rect 22428 38892 22708 38894
rect 22428 38882 22484 38892
rect 22652 38668 22708 38892
rect 22820 38890 22876 39340
rect 22820 38838 22822 38890
rect 22874 38838 22876 38890
rect 22988 39172 23044 39182
rect 22988 38946 23044 39116
rect 22988 38894 22990 38946
rect 23042 38894 23044 38946
rect 22988 38882 23044 38894
rect 22820 38826 22876 38838
rect 23212 38834 23268 40348
rect 23436 40404 23492 40414
rect 23772 40404 23828 40414
rect 23436 40402 23828 40404
rect 23436 40350 23438 40402
rect 23490 40350 23774 40402
rect 23826 40350 23828 40402
rect 23436 40348 23828 40350
rect 23436 40338 23492 40348
rect 23772 40338 23828 40348
rect 23940 40404 23996 40518
rect 23940 40338 23996 40348
rect 24444 40292 24500 40302
rect 24444 40198 24500 40236
rect 23436 40180 23492 40190
rect 23212 38782 23214 38834
rect 23266 38782 23268 38834
rect 23212 38770 23268 38782
rect 23324 39618 23380 39630
rect 23324 39566 23326 39618
rect 23378 39566 23380 39618
rect 23324 38724 23380 39566
rect 23436 38948 23492 40124
rect 24332 39732 24388 39742
rect 24108 39620 24164 39630
rect 24108 39526 24164 39564
rect 23436 38862 23492 38892
rect 23436 38810 23438 38862
rect 23490 38810 23492 38862
rect 23436 38798 23492 38810
rect 23548 39508 23604 39518
rect 23324 38668 23492 38724
rect 22652 38612 23268 38668
rect 22316 37998 22318 38050
rect 22370 37998 22372 38050
rect 22316 37828 22372 37998
rect 22988 38052 23044 38062
rect 22988 37958 23044 37996
rect 23100 38050 23156 38062
rect 23100 37998 23102 38050
rect 23154 37998 23156 38050
rect 22708 37940 22764 37950
rect 22708 37938 22932 37940
rect 22708 37886 22710 37938
rect 22762 37886 22932 37938
rect 22708 37884 22932 37886
rect 22708 37874 22764 37884
rect 22316 37762 22372 37772
rect 21980 37538 22036 37548
rect 22652 37380 22708 37390
rect 22316 37268 22372 37278
rect 22316 37174 22372 37212
rect 22652 37266 22708 37324
rect 22652 37214 22654 37266
rect 22706 37214 22708 37266
rect 22652 37202 22708 37214
rect 22876 37266 22932 37884
rect 22876 37214 22878 37266
rect 22930 37214 22932 37266
rect 22876 37156 22932 37214
rect 23100 37268 23156 37998
rect 23212 38052 23268 38612
rect 23324 38052 23380 38062
rect 23212 38050 23380 38052
rect 23212 37998 23326 38050
rect 23378 37998 23380 38050
rect 23212 37996 23380 37998
rect 23324 37986 23380 37996
rect 23436 37940 23492 38668
rect 23548 38050 23604 39452
rect 24332 38948 24388 39676
rect 24668 38958 24724 41132
rect 26012 41188 26068 41198
rect 26012 41094 26068 41132
rect 26236 41186 26292 41198
rect 26236 41134 26238 41186
rect 26290 41134 26292 41186
rect 24780 41076 24836 41086
rect 24780 40402 24836 41020
rect 25732 41076 25788 41086
rect 25732 40982 25788 41020
rect 26236 40964 26292 41134
rect 26236 40898 26292 40908
rect 26460 40740 26516 41246
rect 26908 41188 26964 41198
rect 26908 41186 27076 41188
rect 26012 40684 26516 40740
rect 26572 41142 26628 41154
rect 26572 41090 26574 41142
rect 26626 41090 26628 41142
rect 26908 41134 26910 41186
rect 26962 41134 27076 41186
rect 26908 41132 27076 41134
rect 26908 41122 26964 41132
rect 24780 40350 24782 40402
rect 24834 40350 24836 40402
rect 24780 40338 24836 40350
rect 25116 40404 25172 40414
rect 24108 38834 24164 38846
rect 24108 38782 24110 38834
rect 24162 38782 24164 38834
rect 24108 38164 24164 38782
rect 24332 38834 24388 38892
rect 24612 38946 24724 38958
rect 24612 38894 24614 38946
rect 24666 38894 24724 38946
rect 24612 38892 24724 38894
rect 24892 39618 24948 39630
rect 24892 39566 24894 39618
rect 24946 39566 24948 39618
rect 24612 38882 24668 38892
rect 24332 38782 24334 38834
rect 24386 38782 24388 38834
rect 24332 38770 24388 38782
rect 24892 38218 24948 39566
rect 24892 38166 24894 38218
rect 24946 38166 24948 38218
rect 24892 38154 24948 38166
rect 25116 38834 25172 40348
rect 25900 40292 25956 40302
rect 25900 40198 25956 40236
rect 25116 38782 25118 38834
rect 25170 38782 25172 38834
rect 23548 37998 23550 38050
rect 23602 37998 23604 38050
rect 23548 37986 23604 37998
rect 23660 38052 23716 38062
rect 23436 37874 23492 37884
rect 23100 37202 23156 37212
rect 23436 37268 23492 37278
rect 23436 37174 23492 37212
rect 23660 37266 23716 37996
rect 23828 38052 23884 38062
rect 23828 37958 23884 37996
rect 24108 38050 24164 38108
rect 24108 37998 24110 38050
rect 24162 37998 24164 38050
rect 23940 37604 23996 37614
rect 23940 37378 23996 37548
rect 23940 37326 23942 37378
rect 23994 37326 23996 37378
rect 23940 37314 23996 37326
rect 23660 37214 23662 37266
rect 23714 37214 23716 37266
rect 23660 37202 23716 37214
rect 22876 37090 22932 37100
rect 21868 36978 21924 36988
rect 22652 37044 22708 37054
rect 23156 37044 23212 37054
rect 21644 36430 21646 36482
rect 21698 36430 21700 36482
rect 21420 36418 21476 36428
rect 21644 36418 21700 36430
rect 21756 36650 21812 36662
rect 21756 36598 21758 36650
rect 21810 36598 21812 36650
rect 21756 36484 21812 36598
rect 22148 36596 22204 36606
rect 22148 36502 22204 36540
rect 21756 36418 21812 36428
rect 21980 36484 22036 36494
rect 20412 36403 20468 36415
rect 20188 35758 20190 35810
rect 20242 35758 20244 35810
rect 20188 35746 20244 35758
rect 21868 36372 21924 36382
rect 15820 35700 15876 35710
rect 16156 35700 16212 35710
rect 16380 35700 16436 35710
rect 15820 35698 16212 35700
rect 15820 35646 15822 35698
rect 15874 35646 16158 35698
rect 16210 35646 16212 35698
rect 15820 35644 16212 35646
rect 15820 35634 15876 35644
rect 16156 35634 16212 35644
rect 16268 35698 16436 35700
rect 16268 35646 16382 35698
rect 16434 35646 16436 35698
rect 16268 35644 16436 35646
rect 15148 34862 15150 34914
rect 15202 34862 15204 34914
rect 15148 34850 15204 34862
rect 15484 34804 15540 34814
rect 15484 34802 15988 34804
rect 15484 34750 15486 34802
rect 15538 34750 15988 34802
rect 15484 34748 15988 34750
rect 15484 34738 15540 34748
rect 13692 34242 13860 34244
rect 13692 34190 13694 34242
rect 13746 34190 13860 34242
rect 13692 34188 13860 34190
rect 14812 34690 14868 34702
rect 14812 34638 14814 34690
rect 14866 34638 14868 34690
rect 13692 34178 13748 34188
rect 14028 34130 14084 34142
rect 14028 34078 14030 34130
rect 14082 34078 14084 34130
rect 14028 33796 14084 34078
rect 14812 34130 14868 34638
rect 14812 34078 14814 34130
rect 14866 34078 14868 34130
rect 14812 34066 14868 34078
rect 14028 33730 14084 33740
rect 14812 33796 14868 33806
rect 13132 33618 13188 33628
rect 12908 33394 12964 33404
rect 12460 33346 12516 33358
rect 12460 33294 12462 33346
rect 12514 33294 12516 33346
rect 12460 33236 12516 33294
rect 12012 32844 12292 32900
rect 12236 32674 12292 32844
rect 12236 32622 12238 32674
rect 12290 32622 12292 32674
rect 12236 32610 12292 32622
rect 9660 32498 9716 32508
rect 10332 32564 10388 32574
rect 10332 32470 10388 32508
rect 8316 32450 8372 32462
rect 8316 32398 8318 32450
rect 8370 32398 8372 32450
rect 8316 32340 8372 32398
rect 8316 32274 8372 32284
rect 12460 32340 12516 33180
rect 12460 32274 12516 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 14700 31556 14756 31566
rect 13468 31554 14756 31556
rect 13468 31502 14702 31554
rect 14754 31502 14756 31554
rect 13468 31500 14756 31502
rect 12684 30994 12740 31006
rect 12684 30942 12686 30994
rect 12738 30942 12740 30994
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 12684 29204 12740 30942
rect 13468 30994 13524 31500
rect 14700 31490 14756 31500
rect 14812 31108 14868 33740
rect 15820 33684 15876 33694
rect 15820 33570 15876 33628
rect 15820 33518 15822 33570
rect 15874 33518 15876 33570
rect 15820 33506 15876 33518
rect 15932 33348 15988 34748
rect 15932 33282 15988 33292
rect 16156 33460 16212 33470
rect 16156 33346 16212 33404
rect 16156 33294 16158 33346
rect 16210 33294 16212 33346
rect 16156 33282 16212 33294
rect 15036 32340 15092 32350
rect 15036 31778 15092 32284
rect 15036 31726 15038 31778
rect 15090 31726 15092 31778
rect 15036 31714 15092 31726
rect 15596 31780 15652 31790
rect 15596 31686 15652 31724
rect 15708 31778 15764 31790
rect 15708 31726 15710 31778
rect 15762 31726 15764 31778
rect 15316 31668 15372 31678
rect 13468 30942 13470 30994
rect 13522 30942 13524 30994
rect 13468 30930 13524 30942
rect 14700 31052 14868 31108
rect 15148 31666 15372 31668
rect 15148 31614 15318 31666
rect 15370 31614 15372 31666
rect 15148 31612 15372 31614
rect 13916 30548 13972 30558
rect 13916 30210 13972 30492
rect 13916 30158 13918 30210
rect 13970 30158 13972 30210
rect 13916 30146 13972 30158
rect 14028 30212 14084 30222
rect 14700 30212 14756 31052
rect 15148 30548 15204 31612
rect 15316 31602 15372 31612
rect 15708 31332 15764 31726
rect 16268 31780 16324 35644
rect 16380 35634 16436 35644
rect 17276 35700 17332 35710
rect 17276 35698 17556 35700
rect 17276 35646 17278 35698
rect 17330 35646 17556 35698
rect 17276 35644 17556 35646
rect 17276 35634 17332 35644
rect 17388 34916 17444 34926
rect 17388 34822 17444 34860
rect 17276 34130 17332 34142
rect 17276 34078 17278 34130
rect 17330 34078 17332 34130
rect 16716 34020 16772 34030
rect 16380 34018 16772 34020
rect 16380 33966 16718 34018
rect 16770 33966 16772 34018
rect 16380 33964 16772 33966
rect 16380 33346 16436 33964
rect 16716 33954 16772 33964
rect 17276 33684 17332 34078
rect 17276 33618 17332 33628
rect 17500 33582 17556 35644
rect 17612 35476 17668 35486
rect 17612 35474 18116 35476
rect 17612 35422 17614 35474
rect 17666 35422 18116 35474
rect 17612 35420 18116 35422
rect 17612 35410 17668 35420
rect 18060 34130 18116 35420
rect 21420 35364 21476 35374
rect 21868 35364 21924 36316
rect 21420 35138 21476 35308
rect 21420 35086 21422 35138
rect 21474 35086 21476 35138
rect 21420 35074 21476 35086
rect 21756 35308 21924 35364
rect 18060 34078 18062 34130
rect 18114 34078 18116 34130
rect 18060 34066 18116 34078
rect 18172 34914 18228 34926
rect 18172 34862 18174 34914
rect 18226 34862 18228 34914
rect 18172 33796 18228 34862
rect 18060 33740 18172 33796
rect 16772 33572 16828 33582
rect 17500 33570 17612 33582
rect 17500 33518 17558 33570
rect 17610 33518 17612 33570
rect 17500 33516 17612 33518
rect 16772 33478 16828 33516
rect 17556 33506 17612 33516
rect 16380 33294 16382 33346
rect 16434 33294 16436 33346
rect 16380 33282 16436 33294
rect 16492 33348 16548 33358
rect 17052 33348 17108 33358
rect 16492 33346 16660 33348
rect 16492 33294 16494 33346
rect 16546 33294 16660 33346
rect 16492 33292 16660 33294
rect 16492 33282 16548 33292
rect 16268 31714 16324 31724
rect 16604 32676 16660 33292
rect 17052 33254 17108 33292
rect 17276 33348 17332 33358
rect 17276 33346 17668 33348
rect 17276 33294 17278 33346
rect 17330 33294 17668 33346
rect 17276 33292 17668 33294
rect 17276 33282 17332 33292
rect 16492 31556 16548 31566
rect 15372 31276 15764 31332
rect 15932 31554 16548 31556
rect 15932 31502 16494 31554
rect 16546 31502 16548 31554
rect 15932 31500 16548 31502
rect 15372 31106 15428 31276
rect 15372 31054 15374 31106
rect 15426 31054 15428 31106
rect 15372 31042 15428 31054
rect 15148 30482 15204 30492
rect 14028 30210 14756 30212
rect 14028 30158 14030 30210
rect 14082 30158 14756 30210
rect 14028 30156 14756 30158
rect 14812 30212 14868 30222
rect 14028 30146 14084 30156
rect 14812 30118 14868 30156
rect 13580 29988 13636 29998
rect 13580 29986 14308 29988
rect 13580 29934 13582 29986
rect 13634 29934 14308 29986
rect 13580 29932 14308 29934
rect 13580 29922 13636 29932
rect 12684 29138 12740 29148
rect 13468 29426 13524 29438
rect 13468 29374 13470 29426
rect 13522 29374 13524 29426
rect 13468 29204 13524 29374
rect 14252 29426 14308 29932
rect 14252 29374 14254 29426
rect 14306 29374 14308 29426
rect 14252 29362 14308 29374
rect 13468 29138 13524 29148
rect 15148 29092 15204 29102
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 15148 28642 15204 29036
rect 15932 28754 15988 31500
rect 16492 31490 16548 31500
rect 16268 30994 16324 31006
rect 16268 30942 16270 30994
rect 16322 30942 16324 30994
rect 15932 28702 15934 28754
rect 15986 28702 15988 28754
rect 15932 28690 15988 28702
rect 16044 30212 16100 30222
rect 15148 28590 15150 28642
rect 15202 28590 15204 28642
rect 15148 28578 15204 28590
rect 16044 28420 16100 30156
rect 16156 29540 16212 29550
rect 16268 29540 16324 30942
rect 16492 30996 16548 31006
rect 16604 30996 16660 32620
rect 17444 32340 17500 32350
rect 17444 32246 17500 32284
rect 16828 31780 16884 31790
rect 17612 31780 17668 33292
rect 17948 33124 18004 33134
rect 17724 32676 17780 32686
rect 17724 32562 17780 32620
rect 17724 32510 17726 32562
rect 17778 32510 17780 32562
rect 17724 32498 17780 32510
rect 17948 32562 18004 33068
rect 17948 32510 17950 32562
rect 18002 32510 18004 32562
rect 17948 32498 18004 32510
rect 18060 31892 18116 33740
rect 18172 33730 18228 33740
rect 18284 34914 18340 34926
rect 18284 34862 18286 34914
rect 18338 34862 18340 34914
rect 18284 33572 18340 34862
rect 18620 34916 18676 34926
rect 18620 34822 18676 34860
rect 21756 34914 21812 35308
rect 21980 35252 22036 36428
rect 22428 36482 22484 36494
rect 22428 36430 22430 36482
rect 22482 36430 22484 36482
rect 22428 36260 22484 36430
rect 22652 36482 22708 36988
rect 23100 37042 23212 37044
rect 23100 36990 23158 37042
rect 23210 36990 23212 37042
rect 23100 36978 23212 36990
rect 24108 37044 24164 37998
rect 24444 38052 24500 38062
rect 24444 37958 24500 37996
rect 25004 38050 25060 38062
rect 25004 37998 25006 38050
rect 25058 37998 25060 38050
rect 25004 37940 25060 37998
rect 25004 37874 25060 37884
rect 24108 36978 24164 36988
rect 22988 36596 23044 36606
rect 22652 36430 22654 36482
rect 22706 36430 22708 36482
rect 22652 36418 22708 36430
rect 22764 36484 22820 36494
rect 22764 36390 22820 36428
rect 22988 36482 23044 36540
rect 22988 36430 22990 36482
rect 23042 36430 23044 36482
rect 22988 36418 23044 36430
rect 23100 36260 23156 36978
rect 23268 36372 23324 36382
rect 23268 36278 23324 36316
rect 22428 36204 23156 36260
rect 22876 35698 22932 35710
rect 22876 35646 22878 35698
rect 22930 35646 22932 35698
rect 22092 35586 22148 35598
rect 22092 35534 22094 35586
rect 22146 35534 22148 35586
rect 22092 35364 22148 35534
rect 22092 35298 22148 35308
rect 22876 35588 22932 35646
rect 23436 35700 23492 35710
rect 23268 35588 23324 35598
rect 22876 35586 23324 35588
rect 22876 35534 23270 35586
rect 23322 35534 23324 35586
rect 22876 35532 23324 35534
rect 21756 34862 21758 34914
rect 21810 34862 21812 34914
rect 21756 34850 21812 34862
rect 21868 35196 22036 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 18284 33506 18340 33516
rect 19964 34018 20020 34030
rect 19964 33966 19966 34018
rect 20018 33966 20020 34018
rect 18396 33348 18452 33358
rect 18172 33236 18228 33246
rect 18172 32564 18228 33180
rect 18172 32498 18228 32508
rect 16828 31778 17556 31780
rect 16828 31726 16830 31778
rect 16882 31726 17556 31778
rect 16828 31724 17556 31726
rect 16828 31714 16884 31724
rect 17388 31556 17444 31566
rect 16492 30994 16660 30996
rect 16492 30942 16494 30994
rect 16546 30942 16660 30994
rect 16492 30940 16660 30942
rect 17052 31554 17444 31556
rect 17052 31502 17390 31554
rect 17442 31502 17444 31554
rect 17052 31500 17444 31502
rect 16492 30930 16548 30940
rect 16772 30772 16828 30782
rect 16772 30770 16996 30772
rect 16772 30718 16774 30770
rect 16826 30718 16996 30770
rect 16772 30716 16996 30718
rect 16772 30706 16828 30716
rect 16716 30548 16772 30558
rect 16716 30210 16772 30492
rect 16716 30158 16718 30210
rect 16770 30158 16772 30210
rect 16716 30146 16772 30158
rect 16156 29538 16324 29540
rect 16156 29486 16158 29538
rect 16210 29486 16324 29538
rect 16156 29484 16324 29486
rect 16156 29474 16212 29484
rect 16940 28980 16996 30716
rect 17052 30210 17108 31500
rect 17388 31490 17444 31500
rect 17500 31118 17556 31724
rect 17444 31106 17556 31118
rect 17444 31054 17446 31106
rect 17498 31054 17556 31106
rect 17444 31052 17556 31054
rect 17444 31042 17500 31052
rect 17612 30996 17668 31724
rect 17724 31890 18116 31892
rect 17724 31838 18062 31890
rect 18114 31838 18116 31890
rect 17724 31836 18116 31838
rect 17724 31778 17780 31836
rect 18060 31826 18116 31836
rect 18396 32004 18452 33292
rect 19964 33124 20020 33966
rect 20076 33346 20132 33358
rect 20860 33348 20916 33358
rect 20076 33294 20078 33346
rect 20130 33294 20132 33346
rect 20076 33124 20132 33294
rect 20412 33346 20916 33348
rect 20412 33294 20862 33346
rect 20914 33294 20916 33346
rect 20412 33292 20916 33294
rect 20076 33068 20244 33124
rect 19964 33058 20020 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19124 32844 19684 32900
rect 19836 32890 20100 32900
rect 19124 32674 19180 32844
rect 19628 32788 19684 32844
rect 20076 32788 20132 32798
rect 20188 32788 20244 33068
rect 19628 32732 19796 32788
rect 19124 32622 19126 32674
rect 19178 32622 19180 32674
rect 19124 32610 19180 32622
rect 19292 32676 19348 32686
rect 19292 32564 19348 32620
rect 19404 32564 19460 32574
rect 19292 32562 19460 32564
rect 19292 32510 19406 32562
rect 19458 32510 19460 32562
rect 19292 32508 19460 32510
rect 18396 31948 18900 32004
rect 17724 31726 17726 31778
rect 17778 31726 17780 31778
rect 17724 31714 17780 31726
rect 18396 31778 18452 31948
rect 18844 31890 18900 31948
rect 18844 31838 18846 31890
rect 18898 31838 18900 31890
rect 18844 31826 18900 31838
rect 18396 31726 18398 31778
rect 18450 31726 18452 31778
rect 18396 31714 18452 31726
rect 18508 31780 18564 31790
rect 18508 31778 18788 31780
rect 18508 31726 18510 31778
rect 18562 31726 18788 31778
rect 18508 31724 18788 31726
rect 18508 31714 18564 31724
rect 18396 31220 18452 31230
rect 17948 31218 18452 31220
rect 17948 31166 18398 31218
rect 18450 31166 18452 31218
rect 17948 31164 18452 31166
rect 17724 30996 17780 31006
rect 17612 30994 17780 30996
rect 17612 30942 17726 30994
rect 17778 30942 17780 30994
rect 17612 30940 17780 30942
rect 17724 30324 17780 30940
rect 17836 30994 17892 31006
rect 17836 30942 17838 30994
rect 17890 30942 17892 30994
rect 17836 30660 17892 30942
rect 17836 30594 17892 30604
rect 17724 30258 17780 30268
rect 17836 30324 17892 30334
rect 17948 30324 18004 31164
rect 18396 31154 18452 31164
rect 17836 30322 18004 30324
rect 17836 30270 17838 30322
rect 17890 30270 18004 30322
rect 17836 30268 18004 30270
rect 18060 30994 18116 31006
rect 18060 30942 18062 30994
rect 18114 30942 18116 30994
rect 17836 30258 17892 30268
rect 17052 30158 17054 30210
rect 17106 30158 17108 30210
rect 17052 29204 17108 30158
rect 18060 29550 18116 30942
rect 18732 30548 18788 31724
rect 18732 30492 19012 30548
rect 18620 29988 18676 29998
rect 18620 29650 18676 29932
rect 18956 29652 19012 30492
rect 18620 29598 18622 29650
rect 18674 29598 18676 29650
rect 18620 29586 18676 29598
rect 18844 29596 19012 29652
rect 18060 29538 18172 29550
rect 18060 29486 18118 29538
rect 18170 29486 18172 29538
rect 18060 29484 18172 29486
rect 18116 29474 18172 29484
rect 17052 29138 17108 29148
rect 17724 29426 17780 29438
rect 17724 29374 17726 29426
rect 17778 29374 17780 29426
rect 16940 28924 17108 28980
rect 16044 28364 16548 28420
rect 16492 28082 16548 28364
rect 16492 28030 16494 28082
rect 16546 28030 16548 28082
rect 16492 28018 16548 28030
rect 10444 27860 10500 27870
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 10108 27076 10164 27086
rect 9716 27074 10164 27076
rect 9716 27022 10110 27074
rect 10162 27022 10164 27074
rect 9716 27020 10164 27022
rect 9716 26514 9772 27020
rect 10108 27010 10164 27020
rect 9716 26462 9718 26514
rect 9770 26462 9772 26514
rect 9716 26450 9772 26462
rect 10444 26334 10500 27804
rect 11788 27860 11844 27870
rect 11788 27766 11844 27804
rect 12796 27860 12852 27870
rect 11620 27636 11676 27646
rect 11004 27634 11676 27636
rect 11004 27582 11622 27634
rect 11674 27582 11676 27634
rect 11004 27580 11676 27582
rect 10892 27076 10948 27086
rect 9884 26290 9940 26302
rect 9884 26238 9886 26290
rect 9938 26238 9940 26290
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 9884 25284 9940 26238
rect 10220 26292 10276 26302
rect 10444 26282 10446 26334
rect 10498 26282 10500 26334
rect 10444 26270 10500 26282
rect 10556 27074 10948 27076
rect 10556 27022 10894 27074
rect 10946 27022 10948 27074
rect 10556 27020 10948 27022
rect 10220 26198 10276 26236
rect 10556 26178 10612 27020
rect 10892 27010 10948 27020
rect 10780 26292 10836 26302
rect 11004 26292 11060 27580
rect 11620 27570 11676 27580
rect 12796 27186 12852 27804
rect 16828 27860 16884 27870
rect 17052 27860 17108 28924
rect 17724 28756 17780 29374
rect 17836 29426 17892 29438
rect 17836 29374 17838 29426
rect 17890 29374 17892 29426
rect 17836 29316 17892 29374
rect 17836 29250 17892 29260
rect 17836 28756 17892 28766
rect 17724 28754 17892 28756
rect 17724 28702 17838 28754
rect 17890 28702 17892 28754
rect 17724 28700 17892 28702
rect 17836 28690 17892 28700
rect 16828 27858 17108 27860
rect 16828 27806 16830 27858
rect 16882 27806 17108 27858
rect 16828 27804 17108 27806
rect 16828 27794 16884 27804
rect 14140 27300 14196 27310
rect 18844 27300 18900 29596
rect 18956 29426 19012 29438
rect 18956 29374 18958 29426
rect 19010 29374 19012 29426
rect 18956 29316 19012 29374
rect 18956 29250 19012 29260
rect 12796 27134 12798 27186
rect 12850 27134 12852 27186
rect 12796 27122 12852 27134
rect 13916 27244 14140 27300
rect 10780 26290 11060 26292
rect 10780 26238 10782 26290
rect 10834 26238 11060 26290
rect 10780 26236 11060 26238
rect 12684 26292 12740 26302
rect 13804 26292 13860 26302
rect 10780 26226 10836 26236
rect 10556 26126 10558 26178
rect 10610 26126 10612 26178
rect 10556 26114 10612 26126
rect 11564 26178 11620 26190
rect 11564 26126 11566 26178
rect 11618 26126 11620 26178
rect 11564 25844 11620 26126
rect 11564 25788 12068 25844
rect 11116 25508 11172 25518
rect 9884 25218 9940 25228
rect 10332 25394 10388 25406
rect 10332 25342 10334 25394
rect 10386 25342 10388 25394
rect 10332 25284 10388 25342
rect 10332 25218 10388 25228
rect 10892 25172 10948 25182
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 10276 24052 10332 24062
rect 10276 23958 10332 23996
rect 10892 24052 10948 25116
rect 11116 24174 11172 25452
rect 11060 24162 11172 24174
rect 11060 24110 11062 24162
rect 11114 24110 11172 24162
rect 11060 24108 11172 24110
rect 11228 25284 11284 25294
rect 11060 24098 11116 24108
rect 10892 23938 10948 23996
rect 10780 23882 10836 23894
rect 10780 23830 10782 23882
rect 10834 23830 10836 23882
rect 10892 23886 10894 23938
rect 10946 23886 10948 23938
rect 10892 23874 10948 23886
rect 10612 23716 10668 23726
rect 10444 23714 10668 23716
rect 10444 23662 10614 23714
rect 10666 23662 10668 23714
rect 10444 23660 10668 23662
rect 9884 23268 9940 23278
rect 10444 23268 10500 23660
rect 10612 23650 10668 23660
rect 9884 23198 9940 23212
rect 9660 23154 9716 23166
rect 9660 23102 9662 23154
rect 9714 23102 9716 23154
rect 9884 23146 9886 23198
rect 9938 23146 9940 23198
rect 9884 23134 9940 23146
rect 10108 23212 10500 23268
rect 10556 23268 10612 23278
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 8428 22146 8484 22158
rect 8428 22094 8430 22146
rect 8482 22094 8484 22146
rect 8092 21586 8148 21598
rect 8092 21534 8094 21586
rect 8146 21534 8148 21586
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 6300 20692 6356 20702
rect 6300 20598 6356 20636
rect 8092 20692 8148 21534
rect 8260 21588 8316 21598
rect 8428 21588 8484 22094
rect 8540 21588 8596 21598
rect 8428 21586 8596 21588
rect 8428 21534 8542 21586
rect 8594 21534 8596 21586
rect 8428 21532 8596 21534
rect 8260 21418 8316 21532
rect 8540 21522 8596 21532
rect 9436 21588 9492 21598
rect 9436 21494 9492 21532
rect 8260 21366 8262 21418
rect 8314 21366 8316 21418
rect 9660 21476 9716 23102
rect 9996 23042 10052 23054
rect 9996 22990 9998 23042
rect 10050 22990 10052 23042
rect 9772 22932 9828 22942
rect 9772 22342 9828 22876
rect 9772 22290 9774 22342
rect 9826 22290 9828 22342
rect 9772 22278 9828 22290
rect 9996 21812 10052 22990
rect 10108 22370 10164 23212
rect 10556 23198 10612 23212
rect 10556 23146 10558 23198
rect 10610 23146 10612 23198
rect 10556 23134 10612 23146
rect 10444 23044 10500 23054
rect 10780 23044 10836 23830
rect 11228 23828 11284 25228
rect 11452 25284 11508 25294
rect 11452 24050 11508 25228
rect 11452 23998 11454 24050
rect 11506 23998 11508 24050
rect 11452 23986 11508 23998
rect 11676 24498 11732 24510
rect 11676 24446 11678 24498
rect 11730 24446 11732 24498
rect 11564 23894 11620 23906
rect 11564 23842 11566 23894
rect 11618 23842 11620 23894
rect 11564 23828 11620 23842
rect 11228 23772 11620 23828
rect 11676 23268 11732 24446
rect 12012 24052 12068 25788
rect 12236 25506 12292 25518
rect 12236 25454 12238 25506
rect 12290 25454 12292 25506
rect 12236 25284 12292 25454
rect 12236 25218 12292 25228
rect 12348 25396 12404 25406
rect 12236 24052 12292 24062
rect 12012 24050 12292 24052
rect 12012 23998 12238 24050
rect 12290 23998 12292 24050
rect 12012 23996 12292 23998
rect 12236 23986 12292 23996
rect 11900 23938 11956 23950
rect 11900 23886 11902 23938
rect 11954 23886 11956 23938
rect 11900 23716 11956 23886
rect 12348 23923 12404 25340
rect 12684 23940 12740 26236
rect 13580 26290 13860 26292
rect 13580 26238 13806 26290
rect 13858 26238 13860 26290
rect 13580 26236 13860 26238
rect 13468 26180 13524 26190
rect 13356 26178 13524 26180
rect 13356 26126 13470 26178
rect 13522 26126 13524 26178
rect 13356 26124 13524 26126
rect 13020 25508 13076 25518
rect 13020 25414 13076 25452
rect 13356 25396 13412 26124
rect 13468 26114 13524 26124
rect 13580 25508 13636 26236
rect 13804 26226 13860 26236
rect 12348 23871 12350 23923
rect 12402 23871 12404 23923
rect 12348 23859 12404 23871
rect 12460 23938 12740 23940
rect 12460 23886 12686 23938
rect 12738 23886 12740 23938
rect 12460 23884 12740 23886
rect 12460 23716 12516 23884
rect 12684 23874 12740 23884
rect 13020 24749 13076 24761
rect 13020 24697 13022 24749
rect 13074 24697 13076 24749
rect 11900 23660 12516 23716
rect 11676 23202 11732 23212
rect 10892 23156 10948 23166
rect 10892 23062 10948 23100
rect 12796 23156 12852 23166
rect 10444 23042 10724 23044
rect 10444 22990 10446 23042
rect 10498 22990 10724 23042
rect 10444 22988 10724 22990
rect 10444 22978 10500 22988
rect 10668 22708 10724 22988
rect 10780 22978 10836 22988
rect 12572 23044 12628 23054
rect 10668 22652 10948 22708
rect 10892 22482 10948 22652
rect 10892 22430 10894 22482
rect 10946 22430 10948 22482
rect 10892 22418 10948 22430
rect 10108 22318 10110 22370
rect 10162 22318 10164 22370
rect 10108 22306 10164 22318
rect 9996 21756 10276 21812
rect 10220 21586 10276 21756
rect 12572 21588 12628 22988
rect 12684 22932 12740 22942
rect 12684 22838 12740 22876
rect 12796 22482 12852 23100
rect 12796 22430 12798 22482
rect 12850 22430 12852 22482
rect 12796 22372 12852 22430
rect 12796 22306 12852 22316
rect 13020 21924 13076 24697
rect 13356 24722 13412 25340
rect 13524 25452 13636 25508
rect 13804 25508 13860 25518
rect 13916 25508 13972 27244
rect 14140 27206 14196 27244
rect 15932 27244 16660 27300
rect 14588 27188 14644 27198
rect 14476 27076 14532 27086
rect 14476 26982 14532 27020
rect 14588 26290 14644 27132
rect 15596 27188 15652 27198
rect 15596 27094 15652 27132
rect 15764 27020 15820 27030
rect 15932 27020 15988 27244
rect 15764 27018 15988 27020
rect 15764 26966 15766 27018
rect 15818 26966 15988 27018
rect 15764 26964 15988 26966
rect 16044 27074 16100 27086
rect 16044 27022 16046 27074
rect 16098 27022 16100 27074
rect 15764 26954 15820 26964
rect 16044 26908 16100 27022
rect 16044 26852 16324 26908
rect 14588 26238 14590 26290
rect 14642 26238 14644 26290
rect 14588 26226 14644 26238
rect 14084 25674 14140 25686
rect 14084 25622 14086 25674
rect 14138 25622 14140 25674
rect 14084 25620 14140 25622
rect 14084 25564 14420 25620
rect 13804 25506 13972 25508
rect 13804 25454 13806 25506
rect 13858 25454 13972 25506
rect 14364 25506 14420 25564
rect 13804 25452 13972 25454
rect 13524 24946 13580 25452
rect 13804 25442 13860 25452
rect 14252 25450 14308 25462
rect 14252 25398 14254 25450
rect 14306 25398 14308 25450
rect 14364 25454 14366 25506
rect 14418 25454 14420 25506
rect 14364 25442 14420 25454
rect 15148 25506 15204 25518
rect 15148 25454 15150 25506
rect 15202 25454 15204 25506
rect 13636 25284 13692 25294
rect 13636 25282 14084 25284
rect 13636 25230 13638 25282
rect 13690 25230 14084 25282
rect 13636 25228 14084 25230
rect 13636 25218 13692 25228
rect 13524 24894 13526 24946
rect 13578 24894 13580 24946
rect 13524 24882 13580 24894
rect 13356 24670 13358 24722
rect 13410 24670 13412 24722
rect 13356 24658 13412 24670
rect 14028 24722 14084 25228
rect 14028 24670 14030 24722
rect 14082 24670 14084 24722
rect 14028 24658 14084 24670
rect 14252 23940 14308 25398
rect 15148 25060 15204 25454
rect 15148 24994 15204 25004
rect 14812 24610 14868 24622
rect 14812 24558 14814 24610
rect 14866 24558 14868 24610
rect 14812 24052 14868 24558
rect 15708 24276 15764 24286
rect 14812 23986 14868 23996
rect 15596 24052 15652 24062
rect 15596 23958 15652 23996
rect 14252 23874 14308 23884
rect 15708 23940 15764 24220
rect 15708 23871 15710 23884
rect 15762 23871 15764 23884
rect 16044 23940 16100 23950
rect 16268 23940 16324 26852
rect 16492 26402 16548 27244
rect 16604 27074 16660 27244
rect 18844 27234 18900 27244
rect 16604 27022 16606 27074
rect 16658 27022 16660 27074
rect 16604 27010 16660 27022
rect 19068 27188 19124 27198
rect 16772 26908 16828 26918
rect 16772 26906 16884 26908
rect 16772 26854 16774 26906
rect 16826 26854 16884 26906
rect 16772 26842 16884 26854
rect 18564 26852 18620 26862
rect 16492 26350 16494 26402
rect 16546 26350 16548 26402
rect 16492 26338 16548 26350
rect 16604 25060 16660 25070
rect 16604 24052 16660 25004
rect 16828 24724 16884 26842
rect 18172 26850 18620 26852
rect 18172 26798 18566 26850
rect 18618 26798 18620 26850
rect 18172 26796 18620 26798
rect 18172 26331 18228 26796
rect 18564 26786 18620 26796
rect 18116 26319 18228 26331
rect 17276 26290 17332 26302
rect 17276 26238 17278 26290
rect 17330 26238 17332 26290
rect 17052 25620 17108 25630
rect 17276 25620 17332 26238
rect 17836 26292 17892 26302
rect 18116 26292 18118 26319
rect 17836 26198 17892 26236
rect 18060 26267 18118 26292
rect 18170 26267 18228 26319
rect 18060 26236 18228 26267
rect 18732 26292 18788 26302
rect 16828 24658 16884 24668
rect 16940 25618 17332 25620
rect 16940 25566 17054 25618
rect 17106 25566 17332 25618
rect 16940 25564 17332 25566
rect 17444 26066 17500 26078
rect 18060 26068 18116 26236
rect 18732 26198 18788 26236
rect 19068 26290 19124 27132
rect 19292 26908 19348 32508
rect 19404 32498 19460 32508
rect 19628 32562 19684 32574
rect 19628 32510 19630 32562
rect 19682 32510 19684 32562
rect 19628 31780 19684 32510
rect 19740 32562 19796 32732
rect 20076 32786 20244 32788
rect 20076 32734 20078 32786
rect 20130 32734 20244 32786
rect 20076 32732 20244 32734
rect 20076 32722 20132 32732
rect 19740 32510 19742 32562
rect 19794 32510 19796 32562
rect 19740 32498 19796 32510
rect 19628 30324 19684 31724
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20076 31014 20132 31026
rect 20076 30962 20078 31014
rect 20130 30962 20132 31014
rect 19908 30770 19964 30782
rect 19908 30718 19910 30770
rect 19962 30718 19964 30770
rect 19740 30324 19796 30334
rect 19628 30322 19796 30324
rect 19628 30270 19742 30322
rect 19794 30270 19796 30322
rect 19628 30268 19796 30270
rect 19740 30258 19796 30268
rect 19908 30212 19964 30718
rect 20076 30436 20132 30962
rect 20188 30996 20244 31006
rect 20188 30994 20356 30996
rect 20188 30942 20190 30994
rect 20242 30942 20356 30994
rect 20188 30940 20356 30942
rect 20188 30930 20244 30940
rect 20076 30370 20132 30380
rect 19908 30146 19964 30156
rect 20300 30210 20356 30940
rect 20300 30158 20302 30210
rect 20354 30158 20356 30210
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19740 29540 19796 29550
rect 19740 29446 19796 29484
rect 20300 29540 20356 30158
rect 20300 29474 20356 29484
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20412 27300 20468 33292
rect 20860 33282 20916 33292
rect 20748 33124 20804 33134
rect 20748 30996 20804 33068
rect 20860 32564 20916 32574
rect 21644 32564 21700 32574
rect 20860 32562 21252 32564
rect 20860 32510 20862 32562
rect 20914 32510 21252 32562
rect 20860 32508 21252 32510
rect 20860 32498 20916 32508
rect 21196 31778 21252 32508
rect 21644 32470 21700 32508
rect 21868 32228 21924 35196
rect 22876 32900 22932 35532
rect 23268 35364 23324 35532
rect 23268 35298 23324 35308
rect 23436 33572 23492 35644
rect 25116 35364 25172 38782
rect 25900 38836 25956 38846
rect 26012 38836 26068 40684
rect 26572 40628 26628 41090
rect 25900 38834 26068 38836
rect 25900 38782 25902 38834
rect 25954 38782 26068 38834
rect 25900 38780 26068 38782
rect 26124 40572 26628 40628
rect 25900 38770 25956 38780
rect 26124 38388 26180 40572
rect 27020 40292 27076 41132
rect 30156 41186 30212 41198
rect 30156 41134 30158 41186
rect 30210 41134 30212 41186
rect 28644 40964 28700 40974
rect 28644 40514 28700 40908
rect 28644 40462 28646 40514
rect 28698 40462 28700 40514
rect 28644 40450 28700 40462
rect 27804 40404 27860 40414
rect 28140 40404 28196 40414
rect 27804 40402 28196 40404
rect 27804 40350 27806 40402
rect 27858 40350 28142 40402
rect 28194 40350 28196 40402
rect 27804 40348 28196 40350
rect 27804 40338 27860 40348
rect 27020 40226 27076 40236
rect 27356 39732 27412 39742
rect 27356 39638 27412 39676
rect 27244 39618 27300 39630
rect 27244 39566 27246 39618
rect 27298 39566 27300 39618
rect 26796 39508 26852 39518
rect 27244 39508 27300 39566
rect 27468 39620 27524 39630
rect 27916 39618 27972 40348
rect 28140 40338 28196 40348
rect 28364 40402 28420 40414
rect 28364 40350 28366 40402
rect 28418 40350 28420 40402
rect 26796 39506 27412 39508
rect 26796 39454 26798 39506
rect 26850 39454 27412 39506
rect 26796 39452 27412 39454
rect 26796 39442 26852 39452
rect 26124 38332 26292 38388
rect 26236 38218 26292 38332
rect 26236 38166 26238 38218
rect 26290 38166 26292 38218
rect 26236 38154 26292 38166
rect 25676 38052 25732 38062
rect 25676 35700 25732 37996
rect 26236 38050 26292 38062
rect 26236 37998 26238 38050
rect 26290 37998 26292 38050
rect 26236 37828 26292 37998
rect 26460 38052 26516 38062
rect 26460 37958 26516 37996
rect 26964 38052 27020 38062
rect 26964 37958 27020 37996
rect 27244 38052 27300 38062
rect 27356 38052 27412 39452
rect 27468 38836 27524 39564
rect 27468 38668 27524 38780
rect 27692 39562 27748 39574
rect 27692 39510 27694 39562
rect 27746 39510 27748 39562
rect 27916 39566 27918 39618
rect 27970 39566 27972 39618
rect 27916 39554 27972 39566
rect 28364 40292 28420 40350
rect 27692 38724 27748 39510
rect 28028 38836 28084 38846
rect 27804 38724 27860 38734
rect 27692 38722 27860 38724
rect 27692 38670 27806 38722
rect 27858 38670 27860 38722
rect 27692 38668 27860 38670
rect 27468 38612 27636 38668
rect 27468 38052 27524 38062
rect 27356 38050 27524 38052
rect 27356 37998 27470 38050
rect 27522 37998 27524 38050
rect 27356 37996 27524 37998
rect 27244 37958 27300 37996
rect 27468 37940 27524 37996
rect 27580 38050 27636 38612
rect 27580 37998 27582 38050
rect 27634 37998 27636 38050
rect 27580 37986 27636 37998
rect 27804 38052 27860 38668
rect 27804 37986 27860 37996
rect 27468 37874 27524 37884
rect 26236 37156 26292 37772
rect 27580 37828 27636 37838
rect 26236 37090 26292 37100
rect 27132 37266 27188 37278
rect 27132 37214 27134 37266
rect 27186 37214 27188 37266
rect 26348 37044 26404 37054
rect 25676 35634 25732 35644
rect 25956 35924 26012 35934
rect 25956 35586 26012 35868
rect 26124 35700 26180 35710
rect 26124 35606 26180 35644
rect 26348 35698 26404 36988
rect 26852 37044 26908 37054
rect 26852 36950 26908 36988
rect 27132 36932 27188 37214
rect 27244 37266 27300 37278
rect 27244 37214 27246 37266
rect 27298 37214 27300 37266
rect 27244 36932 27300 37214
rect 27412 37268 27468 37278
rect 27412 37174 27468 37212
rect 27580 37266 27636 37772
rect 27580 37214 27582 37266
rect 27634 37214 27636 37266
rect 27580 37202 27636 37214
rect 28028 37266 28084 38780
rect 28364 38724 28420 40236
rect 28812 40404 28868 40414
rect 28812 40292 28868 40348
rect 29708 40402 29764 40414
rect 29708 40350 29710 40402
rect 29762 40350 29764 40402
rect 29204 40292 29260 40302
rect 28812 40290 29260 40292
rect 28812 40238 29206 40290
rect 29258 40238 29260 40290
rect 28812 40236 29260 40238
rect 28812 39844 28868 40236
rect 29204 40226 29260 40236
rect 28644 39788 28868 39844
rect 28644 39730 28700 39788
rect 28644 39678 28646 39730
rect 28698 39678 28700 39730
rect 28644 39666 28700 39678
rect 29708 39620 29764 40350
rect 30156 39620 30212 41134
rect 30492 40290 30548 41804
rect 31164 41794 31220 41804
rect 31276 41524 31332 41933
rect 31612 41972 31668 41982
rect 31612 41878 31668 41916
rect 32284 41956 32286 42008
rect 32338 41956 32340 42008
rect 32620 41972 32676 41982
rect 31164 41468 31332 41524
rect 30940 41300 30996 41310
rect 30940 41206 30996 41244
rect 31164 40628 31220 41468
rect 31164 40562 31220 40572
rect 32284 40516 32340 41956
rect 32284 40450 32340 40460
rect 32396 41970 32676 41972
rect 32396 41918 32622 41970
rect 32674 41918 32676 41970
rect 32396 41916 32676 41918
rect 32396 40514 32452 41916
rect 32620 41906 32676 41916
rect 32844 41970 32900 42028
rect 32844 41918 32846 41970
rect 32898 41918 32900 41970
rect 32844 41906 32900 41918
rect 33012 41914 33068 41926
rect 33012 41862 33014 41914
rect 33066 41862 33068 41914
rect 33012 41412 33068 41862
rect 33180 41524 33236 42028
rect 43036 41997 43092 42009
rect 33628 41972 33684 41982
rect 33628 41746 33684 41916
rect 36876 41970 36932 41982
rect 36876 41918 36878 41970
rect 36930 41918 36932 41970
rect 33628 41694 33630 41746
rect 33682 41694 33684 41746
rect 33180 41468 33460 41524
rect 32396 40462 32398 40514
rect 32450 40462 32452 40514
rect 32396 40404 32452 40462
rect 32396 40338 32452 40348
rect 32844 41356 33068 41412
rect 32844 41074 32900 41356
rect 33292 41300 33348 41310
rect 33292 41206 33348 41244
rect 33404 41171 33460 41468
rect 33404 41119 33406 41171
rect 33458 41119 33460 41171
rect 33628 41186 33684 41694
rect 34636 41748 34692 41758
rect 36596 41748 36652 41758
rect 34636 41746 35028 41748
rect 34636 41694 34638 41746
rect 34690 41694 35028 41746
rect 34636 41692 35028 41694
rect 34636 41682 34692 41692
rect 33628 41134 33630 41186
rect 33682 41134 33684 41186
rect 33628 41122 33684 41134
rect 33404 41107 33460 41119
rect 32844 41022 32846 41074
rect 32898 41022 32900 41074
rect 30492 40238 30494 40290
rect 30546 40238 30548 40290
rect 30492 40226 30548 40238
rect 30268 39620 30324 39630
rect 30156 39564 30268 39620
rect 28700 38836 28756 38846
rect 28700 38742 28756 38780
rect 29708 38836 29764 39564
rect 30268 39526 30324 39564
rect 31052 39618 31108 39630
rect 31052 39566 31054 39618
rect 31106 39566 31108 39618
rect 31052 39060 31108 39566
rect 32844 39620 32900 41022
rect 33180 40628 33236 40638
rect 33180 40514 33236 40572
rect 33180 40462 33182 40514
rect 33234 40462 33236 40514
rect 33180 40450 33236 40462
rect 33423 40516 33479 40526
rect 33423 40458 33479 40460
rect 33423 40406 33425 40458
rect 33477 40406 33479 40458
rect 33423 40394 33479 40406
rect 33628 40404 33684 40414
rect 33628 39956 33684 40348
rect 34300 40404 34356 40442
rect 34300 40338 34356 40348
rect 33628 39900 33908 39956
rect 32844 39554 32900 39564
rect 33740 39620 33796 39630
rect 33740 39526 33796 39564
rect 33852 39620 33908 39900
rect 34300 39786 34356 39798
rect 34300 39734 34302 39786
rect 34354 39734 34356 39786
rect 34188 39620 34244 39630
rect 33852 39618 34244 39620
rect 33852 39566 33854 39618
rect 33906 39566 34190 39618
rect 34242 39566 34244 39618
rect 33852 39564 34244 39566
rect 33852 39554 33908 39564
rect 34188 39554 34244 39564
rect 32956 39506 33012 39518
rect 33460 39508 33516 39518
rect 32956 39454 32958 39506
rect 33010 39454 33012 39506
rect 31052 38994 31108 39004
rect 32396 39060 32452 39070
rect 32396 38966 32452 39004
rect 32956 39060 33012 39454
rect 32956 38994 33012 39004
rect 33292 39506 33516 39508
rect 33292 39454 33462 39506
rect 33514 39454 33516 39506
rect 33292 39452 33516 39454
rect 29708 38770 29764 38780
rect 30380 38861 30436 38873
rect 30380 38809 30382 38861
rect 30434 38809 30436 38861
rect 31724 38836 31780 38846
rect 28364 38658 28420 38668
rect 29540 38724 29596 38734
rect 29540 38274 29596 38668
rect 29540 38222 29542 38274
rect 29594 38222 29596 38274
rect 29540 38210 29596 38222
rect 29036 38050 29092 38062
rect 29036 37998 29038 38050
rect 29090 37998 29092 38050
rect 29036 37940 29092 37998
rect 29260 38052 29316 38062
rect 29260 37958 29316 37996
rect 29036 37874 29092 37884
rect 28028 37214 28030 37266
rect 28082 37214 28084 37266
rect 28028 37202 28084 37214
rect 28812 37156 28868 37166
rect 28812 37154 29092 37156
rect 28812 37102 28814 37154
rect 28866 37102 29092 37154
rect 28812 37100 29092 37102
rect 28812 37090 28868 37100
rect 27244 36876 27636 36932
rect 27132 36866 27188 36876
rect 26908 36484 26964 36494
rect 27020 36484 27076 36494
rect 26908 36482 27020 36484
rect 26908 36430 26910 36482
rect 26962 36430 27020 36482
rect 26908 36428 27020 36430
rect 26908 36418 26964 36428
rect 26908 35924 26964 35934
rect 26628 35812 26684 35822
rect 26628 35718 26684 35756
rect 26348 35646 26350 35698
rect 26402 35646 26404 35698
rect 26348 35634 26404 35646
rect 26908 35698 26964 35868
rect 26908 35646 26910 35698
rect 26962 35646 26964 35698
rect 25956 35534 25958 35586
rect 26010 35534 26012 35586
rect 25116 35298 25172 35308
rect 25676 35364 25732 35374
rect 25676 34914 25732 35308
rect 25956 35364 26012 35534
rect 25956 35298 26012 35308
rect 26908 35364 26964 35646
rect 25676 34862 25678 34914
rect 25730 34862 25732 34914
rect 25676 34850 25732 34862
rect 26908 34354 26964 35308
rect 27020 34804 27076 36428
rect 27020 34738 27076 34748
rect 26908 34302 26910 34354
rect 26962 34302 26964 34354
rect 26908 34290 26964 34302
rect 24556 34132 24612 34142
rect 24556 34038 24612 34076
rect 24780 34130 24836 34142
rect 24780 34078 24782 34130
rect 24834 34078 24836 34130
rect 24276 33908 24332 33918
rect 24276 33906 24500 33908
rect 24276 33854 24278 33906
rect 24330 33854 24500 33906
rect 24276 33852 24500 33854
rect 24276 33842 24332 33852
rect 24220 33684 24276 33694
rect 23436 33516 23604 33572
rect 22988 33346 23044 33358
rect 23436 33348 23492 33358
rect 22988 33294 22990 33346
rect 23042 33294 23044 33346
rect 22988 33012 23044 33294
rect 23156 33346 23492 33348
rect 23156 33294 23438 33346
rect 23490 33294 23492 33346
rect 23156 33292 23492 33294
rect 23156 33178 23212 33292
rect 23436 33282 23492 33292
rect 23156 33126 23158 33178
rect 23210 33126 23212 33178
rect 23156 33114 23212 33126
rect 23548 33124 23604 33516
rect 24220 33458 24276 33628
rect 24220 33406 24222 33458
rect 24274 33406 24276 33458
rect 24220 33394 24276 33406
rect 24444 33348 24500 33852
rect 24780 33796 24836 34078
rect 25452 34132 25508 34142
rect 24780 33730 24836 33740
rect 25284 33906 25340 33918
rect 25284 33854 25286 33906
rect 25338 33854 25340 33906
rect 25284 33684 25340 33854
rect 25284 33618 25340 33628
rect 25452 33460 25508 34076
rect 24444 33282 24500 33292
rect 25340 33404 25452 33460
rect 23436 33068 23604 33124
rect 24668 33124 24724 33134
rect 25340 33124 25396 33404
rect 25452 33394 25508 33404
rect 26124 33460 26180 33470
rect 26124 33366 26180 33404
rect 22988 32956 23268 33012
rect 22876 32844 23156 32900
rect 21868 32172 22148 32228
rect 21196 31726 21198 31778
rect 21250 31726 21252 31778
rect 20972 30996 21028 31006
rect 20748 30994 21028 30996
rect 20748 30942 20974 30994
rect 21026 30942 21028 30994
rect 20748 30940 21028 30942
rect 20972 30930 21028 30940
rect 20636 30436 20692 30446
rect 20636 30342 20692 30380
rect 21196 30436 21252 31726
rect 21980 31780 22036 31790
rect 21980 31686 22036 31724
rect 21196 30210 21252 30380
rect 21980 30660 22036 30670
rect 21980 30322 22036 30604
rect 21980 30270 21982 30322
rect 22034 30270 22036 30322
rect 21980 30258 22036 30270
rect 21196 30158 21198 30210
rect 21250 30158 21252 30210
rect 21196 30146 21252 30158
rect 21644 30212 21700 30222
rect 21644 29426 21700 30156
rect 21644 29374 21646 29426
rect 21698 29374 21700 29426
rect 21644 29362 21700 29374
rect 22092 29092 22148 32172
rect 22876 30996 22932 31006
rect 22876 30902 22932 30940
rect 22428 29428 22484 29438
rect 22820 29428 22876 29438
rect 22316 29426 22876 29428
rect 22316 29374 22430 29426
rect 22482 29374 22822 29426
rect 22874 29374 22876 29426
rect 22316 29372 22876 29374
rect 22092 29036 22240 29092
rect 20860 28642 20916 28654
rect 20860 28590 20862 28642
rect 20914 28590 20916 28642
rect 20524 28420 20580 28430
rect 20524 28326 20580 28364
rect 20524 27300 20580 27310
rect 20412 27298 20580 27300
rect 20412 27246 20526 27298
rect 20578 27246 20580 27298
rect 20412 27244 20580 27246
rect 20300 27188 20356 27198
rect 19460 27076 19516 27086
rect 19852 27076 19908 27086
rect 19460 27074 19852 27076
rect 19460 27022 19462 27074
rect 19514 27022 19852 27074
rect 19460 27020 19852 27022
rect 19460 27010 19516 27020
rect 19852 26982 19908 27020
rect 20188 27074 20244 27086
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 19292 26852 19572 26908
rect 19068 26238 19070 26290
rect 19122 26238 19124 26290
rect 19068 26226 19124 26238
rect 17444 26014 17446 26066
rect 17498 26014 17500 26066
rect 16716 24610 16772 24622
rect 16716 24558 16718 24610
rect 16770 24558 16772 24610
rect 16716 24276 16772 24558
rect 16716 24210 16772 24220
rect 16828 24052 16884 24062
rect 16604 24050 16884 24052
rect 16604 23998 16830 24050
rect 16882 23998 16884 24050
rect 16604 23996 16884 23998
rect 16828 23986 16884 23996
rect 16044 23938 16268 23940
rect 16044 23886 16046 23938
rect 16098 23886 16268 23938
rect 16044 23884 16268 23886
rect 16044 23874 16100 23884
rect 15708 23846 15764 23871
rect 16268 23846 16324 23884
rect 16940 23923 16996 25564
rect 17052 25554 17108 25564
rect 17444 25506 17500 26014
rect 17444 25454 17446 25506
rect 17498 25454 17500 25506
rect 17444 25442 17500 25454
rect 17836 26012 18116 26068
rect 18284 26178 18340 26190
rect 18284 26126 18286 26178
rect 18338 26126 18340 26178
rect 17836 25396 17892 26012
rect 18172 25620 18228 25630
rect 18284 25620 18340 26126
rect 18172 25618 18340 25620
rect 18172 25566 18174 25618
rect 18226 25566 18340 25618
rect 18172 25564 18340 25566
rect 19404 26066 19460 26078
rect 19404 26014 19406 26066
rect 19458 26014 19460 26066
rect 18172 25554 18228 25564
rect 17836 25172 17892 25340
rect 17276 24724 17332 24734
rect 17276 24630 17332 24668
rect 16940 23871 16942 23923
rect 16994 23871 16996 23923
rect 16940 23859 16996 23871
rect 17164 23940 17220 23950
rect 17164 23846 17220 23884
rect 13692 23181 13748 23193
rect 13692 23129 13694 23181
rect 13746 23129 13748 23181
rect 13692 22820 13748 23129
rect 14476 23156 14532 23166
rect 14476 23062 14532 23100
rect 15708 23154 15764 23166
rect 15708 23102 15710 23154
rect 15762 23102 15764 23154
rect 14140 22932 14196 22942
rect 15148 22932 15204 22942
rect 14140 22930 14644 22932
rect 14140 22878 14142 22930
rect 14194 22878 14644 22930
rect 14140 22876 14644 22878
rect 14140 22866 14196 22876
rect 13692 22754 13748 22764
rect 13580 22372 13636 22382
rect 13580 22278 13636 22316
rect 14456 22314 14512 22326
rect 14456 22262 14458 22314
rect 14510 22262 14512 22314
rect 14456 21924 14512 22262
rect 13020 21868 13300 21924
rect 14456 21868 14532 21924
rect 10220 21534 10222 21586
rect 10274 21534 10276 21586
rect 10220 21522 10276 21534
rect 12348 21586 12628 21588
rect 12348 21534 12574 21586
rect 12626 21534 12628 21586
rect 12348 21532 12628 21534
rect 12124 21476 12180 21486
rect 8260 21354 8316 21366
rect 8876 21362 8932 21374
rect 8876 21310 8878 21362
rect 8930 21310 8932 21362
rect 8204 20804 8260 20814
rect 8204 20802 8372 20804
rect 8204 20750 8206 20802
rect 8258 20750 8372 20802
rect 8204 20748 8372 20750
rect 8204 20738 8260 20748
rect 8092 20132 8148 20636
rect 8092 20066 8148 20076
rect 8036 19908 8092 19918
rect 8036 19814 8092 19852
rect 8316 19906 8372 20748
rect 8764 20132 8820 20142
rect 8316 19854 8318 19906
rect 8370 19854 8372 19906
rect 8316 19842 8372 19854
rect 8428 20033 8484 20045
rect 8428 19981 8430 20033
rect 8482 19981 8484 20033
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 8428 19460 8484 19981
rect 8428 19394 8484 19404
rect 8764 20018 8820 20076
rect 8764 19966 8766 20018
rect 8818 19966 8820 20018
rect 8764 19348 8820 19966
rect 8764 19282 8820 19292
rect 8372 19236 8428 19246
rect 8372 19066 8428 19180
rect 8372 19014 8374 19066
rect 8426 19014 8428 19066
rect 8372 19002 8428 19014
rect 8540 19234 8596 19246
rect 8540 19182 8542 19234
rect 8594 19182 8596 19234
rect 8316 18564 8372 18574
rect 7980 18226 8036 18238
rect 7980 18174 7982 18226
rect 8034 18174 8036 18226
rect 7980 18116 8036 18174
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 7980 18050 8036 18060
rect 4476 17994 4740 18004
rect 8316 17778 8372 18508
rect 8316 17726 8318 17778
rect 8370 17726 8372 17778
rect 8316 17714 8372 17726
rect 8540 17780 8596 19182
rect 8876 18477 8932 21310
rect 8988 21364 9044 21374
rect 8988 20802 9044 21308
rect 9660 21028 9716 21420
rect 12012 21420 12124 21476
rect 9660 20972 9828 21028
rect 8988 20750 8990 20802
rect 9042 20750 9044 20802
rect 8988 19908 9044 20750
rect 9100 20804 9156 20814
rect 9100 20802 9716 20804
rect 9100 20750 9102 20802
rect 9154 20750 9716 20802
rect 9100 20748 9716 20750
rect 9100 20738 9156 20748
rect 8988 19842 9044 19852
rect 9436 20018 9492 20030
rect 9436 19966 9438 20018
rect 9490 19966 9492 20018
rect 9436 19236 9492 19966
rect 8876 18425 8878 18477
rect 8930 18425 8932 18477
rect 8876 18413 8932 18425
rect 9100 19206 9156 19218
rect 9100 19154 9102 19206
rect 9154 19154 9156 19206
rect 9660 19236 9716 20748
rect 9772 20580 9828 20972
rect 9884 20804 9940 20814
rect 12012 20804 12068 21420
rect 12124 21382 12180 21420
rect 12348 21252 12404 21532
rect 12572 21522 12628 21532
rect 9884 20802 10052 20804
rect 9884 20750 9886 20802
rect 9938 20750 10052 20802
rect 9884 20748 10052 20750
rect 9884 20738 9940 20748
rect 9772 20524 9940 20580
rect 9772 19460 9828 19470
rect 9772 19366 9828 19404
rect 9660 19180 9772 19236
rect 9436 19170 9492 19180
rect 9100 18116 9156 19154
rect 9716 18282 9772 19180
rect 9884 18450 9940 20524
rect 9996 18788 10052 20748
rect 12012 20738 12068 20748
rect 12124 21196 12628 21252
rect 11788 20690 11844 20702
rect 11788 20638 11790 20690
rect 11842 20638 11844 20690
rect 10220 20580 10276 20590
rect 10220 20018 10276 20524
rect 10220 19966 10222 20018
rect 10274 19966 10276 20018
rect 10220 19954 10276 19966
rect 11788 19684 11844 20638
rect 12124 20130 12180 21196
rect 12236 20914 12292 20926
rect 12236 20862 12238 20914
rect 12290 20862 12292 20914
rect 12236 20580 12292 20862
rect 12572 20802 12628 21196
rect 12236 20514 12292 20524
rect 12348 20758 12404 20770
rect 12348 20706 12350 20758
rect 12402 20706 12404 20758
rect 12572 20750 12574 20802
rect 12626 20750 12628 20802
rect 12572 20738 12628 20750
rect 12124 20078 12126 20130
rect 12178 20078 12180 20130
rect 12124 20066 12180 20078
rect 11676 19628 11844 19684
rect 11676 19572 11732 19628
rect 11452 19516 11732 19572
rect 11004 19460 11060 19470
rect 9996 18732 10164 18788
rect 9884 18398 9886 18450
rect 9938 18398 9940 18450
rect 9884 18386 9940 18398
rect 9716 18230 9718 18282
rect 9770 18230 9772 18282
rect 10108 18338 10164 18732
rect 10892 18564 10948 18574
rect 10220 18465 10276 18490
rect 10220 18452 10222 18465
rect 10274 18452 10276 18465
rect 10220 18386 10276 18396
rect 10444 18450 10500 18462
rect 10444 18398 10446 18450
rect 10498 18398 10500 18450
rect 10108 18286 10110 18338
rect 10162 18286 10164 18338
rect 10108 18274 10164 18286
rect 10444 18340 10500 18398
rect 9716 18218 9772 18230
rect 9100 18050 9156 18060
rect 10108 18116 10164 18126
rect 8540 17714 8596 17724
rect 7532 17668 7588 17678
rect 7532 17666 8260 17668
rect 7532 17614 7534 17666
rect 7586 17614 8260 17666
rect 7532 17612 8260 17614
rect 7532 17602 7588 17612
rect 8204 17118 8260 17612
rect 8932 17164 9380 17220
rect 8204 17106 8316 17118
rect 8204 17054 8262 17106
rect 8314 17054 8316 17106
rect 8204 17052 8316 17054
rect 8260 17042 8316 17052
rect 8932 17106 8988 17164
rect 8932 17054 8934 17106
rect 8986 17054 8988 17106
rect 8932 17042 8988 17054
rect 9100 16996 9156 17006
rect 8428 16882 8484 16894
rect 8428 16830 8430 16882
rect 8482 16830 8484 16882
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 8428 16212 8484 16830
rect 8092 16156 8484 16212
rect 8764 16884 8820 16894
rect 7868 16098 7924 16110
rect 7868 16046 7870 16098
rect 7922 16046 7924 16098
rect 7364 15540 7420 15550
rect 7868 15540 7924 16046
rect 7364 15538 7924 15540
rect 7364 15486 7366 15538
rect 7418 15486 7924 15538
rect 7364 15484 7924 15486
rect 7980 15764 8036 15774
rect 8092 15764 8148 16156
rect 8652 16100 8708 16110
rect 8036 15708 8148 15764
rect 8204 16098 8708 16100
rect 8204 16046 8654 16098
rect 8706 16046 8708 16098
rect 8204 16044 8708 16046
rect 7364 15474 7420 15484
rect 7532 15314 7588 15326
rect 7532 15262 7534 15314
rect 7586 15262 7588 15314
rect 7532 15148 7588 15262
rect 7868 15316 7924 15326
rect 7980 15316 8036 15708
rect 7868 15314 8036 15316
rect 7868 15262 7870 15314
rect 7922 15262 8036 15314
rect 7868 15260 8036 15262
rect 8092 15329 8148 15341
rect 8092 15277 8094 15329
rect 8146 15277 8148 15329
rect 7868 15250 7924 15260
rect 8092 15204 8148 15277
rect 7532 15092 7700 15148
rect 8092 15138 8148 15148
rect 8204 15202 8260 16044
rect 8652 16034 8708 16044
rect 8652 15316 8708 15326
rect 8764 15316 8820 16828
rect 9100 16882 9156 16940
rect 9100 16830 9102 16882
rect 9154 16830 9156 16882
rect 9100 16818 9156 16830
rect 9324 16884 9380 17164
rect 9436 16884 9492 16894
rect 9324 16882 9492 16884
rect 9324 16830 9438 16882
rect 9490 16830 9492 16882
rect 9324 16828 9492 16830
rect 9436 16818 9492 16828
rect 8652 15314 8820 15316
rect 8652 15262 8654 15314
rect 8706 15262 8820 15314
rect 8652 15260 8820 15262
rect 8876 16436 8932 16446
rect 8876 15358 8932 16380
rect 8876 15306 8878 15358
rect 8930 15306 8932 15358
rect 8652 15250 8708 15260
rect 8204 15150 8206 15202
rect 8258 15150 8260 15202
rect 8204 15138 8260 15150
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 7532 14756 7588 14766
rect 7532 13746 7588 14700
rect 7644 13860 7700 15092
rect 8428 14756 8484 14766
rect 7644 13794 7700 13804
rect 7756 14530 7812 14542
rect 7756 14478 7758 14530
rect 7810 14478 7812 14530
rect 7756 14420 7812 14478
rect 7532 13694 7534 13746
rect 7586 13694 7588 13746
rect 7532 13682 7588 13694
rect 7756 13746 7812 14364
rect 8428 14530 8484 14700
rect 8764 14644 8820 14654
rect 8764 14550 8820 14588
rect 8428 14478 8430 14530
rect 8482 14478 8484 14530
rect 7924 14308 7980 14318
rect 7924 14306 8036 14308
rect 7924 14254 7926 14306
rect 7978 14254 8036 14306
rect 7924 14242 8036 14254
rect 7756 13694 7758 13746
rect 7810 13694 7812 13746
rect 7756 13682 7812 13694
rect 7364 13522 7420 13534
rect 7364 13470 7366 13522
rect 7418 13470 7420 13522
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 7364 12964 7420 13470
rect 7980 13076 8036 14242
rect 8428 13972 8484 14478
rect 8428 13906 8484 13916
rect 8652 14486 8708 14498
rect 8652 14434 8654 14486
rect 8706 14434 8708 14486
rect 8540 13860 8596 13870
rect 8092 13761 8148 13773
rect 8092 13748 8094 13761
rect 8146 13748 8148 13761
rect 8092 13669 8148 13692
rect 8540 13746 8596 13804
rect 8540 13694 8542 13746
rect 8594 13694 8596 13746
rect 8204 13634 8260 13646
rect 8204 13582 8206 13634
rect 8258 13582 8260 13634
rect 8092 13076 8148 13086
rect 7980 13020 8092 13076
rect 8092 13010 8148 13020
rect 7364 12898 7420 12908
rect 8204 12180 8260 13582
rect 8540 13636 8596 13694
rect 8652 13748 8708 14434
rect 8876 13790 8932 15306
rect 8988 15876 9044 15886
rect 8988 15202 9044 15820
rect 8988 15150 8990 15202
rect 9042 15150 9044 15202
rect 8988 15138 9044 15150
rect 9100 15204 9156 15214
rect 8988 14532 9044 14542
rect 9100 14532 9156 15148
rect 8988 14530 9156 14532
rect 8988 14478 8990 14530
rect 9042 14478 9156 14530
rect 8988 14476 9156 14478
rect 10108 14502 10164 18060
rect 10220 17780 10276 17790
rect 10220 17686 10276 17724
rect 10444 16996 10500 18284
rect 10892 18338 10948 18508
rect 11004 18494 11060 19404
rect 11004 18442 11006 18494
rect 11058 18442 11060 18494
rect 11004 18430 11060 18442
rect 11228 18450 11284 18462
rect 10892 18286 10894 18338
rect 10946 18286 10948 18338
rect 10892 18274 10948 18286
rect 11228 18398 11230 18450
rect 11282 18398 11284 18450
rect 11228 17780 11284 18398
rect 11452 18340 11508 19516
rect 11676 19236 11732 19246
rect 11676 19142 11732 19180
rect 12012 18452 12068 18462
rect 12012 18358 12068 18396
rect 12348 18452 12404 20706
rect 13244 20244 13300 21868
rect 13448 21586 13504 21598
rect 13448 21534 13450 21586
rect 13502 21534 13504 21586
rect 13448 21140 13504 21534
rect 14252 21476 14308 21486
rect 14308 21420 14420 21476
rect 14252 21382 14308 21420
rect 13692 21364 13748 21374
rect 13692 21362 14196 21364
rect 13692 21310 13694 21362
rect 13746 21310 14196 21362
rect 13692 21308 14196 21310
rect 13692 21298 13748 21308
rect 14140 21252 14196 21308
rect 14140 21196 14308 21252
rect 13448 21074 13504 21084
rect 13580 20804 13636 20814
rect 13580 20710 13636 20748
rect 13356 20244 13412 20254
rect 13244 20242 13972 20244
rect 13244 20190 13358 20242
rect 13410 20190 13972 20242
rect 13244 20188 13972 20190
rect 13356 20178 13412 20188
rect 12552 19684 12608 19694
rect 12552 19234 12608 19628
rect 13804 19348 13860 19386
rect 13804 19282 13860 19292
rect 12552 19182 12554 19234
rect 12606 19182 12608 19234
rect 12552 19170 12608 19182
rect 12684 19236 12740 19246
rect 12348 18386 12404 18396
rect 11452 18274 11508 18284
rect 12684 17890 12740 19180
rect 13468 19236 13524 19246
rect 13468 19142 13524 19180
rect 13804 19178 13860 19190
rect 12796 19124 12852 19134
rect 12796 19030 12852 19068
rect 13804 19126 13806 19178
rect 13858 19126 13860 19178
rect 13804 19124 13860 19126
rect 13804 19058 13860 19068
rect 13916 18477 13972 20188
rect 14140 19236 14196 19246
rect 14252 19236 14308 21196
rect 14364 21028 14420 21420
rect 14476 21252 14532 21868
rect 14476 21186 14532 21196
rect 14364 20972 14512 21028
rect 14456 20802 14512 20972
rect 14456 20750 14458 20802
rect 14510 20750 14512 20802
rect 14456 20738 14512 20750
rect 14588 20468 14644 22876
rect 15148 22342 15204 22876
rect 15148 22290 15150 22342
rect 15202 22290 15204 22342
rect 15148 22278 15204 22290
rect 15372 22930 15428 22942
rect 15372 22878 15374 22930
rect 15426 22878 15428 22930
rect 14700 22260 14756 22270
rect 14700 22258 14980 22260
rect 14700 22206 14702 22258
rect 14754 22206 14980 22258
rect 14700 22204 14980 22206
rect 14700 22194 14756 22204
rect 14700 20692 14756 20702
rect 14700 20690 14868 20692
rect 14700 20638 14702 20690
rect 14754 20638 14868 20690
rect 14700 20636 14868 20638
rect 14700 20626 14756 20636
rect 14588 20412 14756 20468
rect 14700 20045 14756 20412
rect 14812 20132 14868 20636
rect 14812 20066 14868 20076
rect 14700 19993 14702 20045
rect 14754 19993 14756 20045
rect 14700 19981 14756 19993
rect 14140 19234 14308 19236
rect 14140 19182 14142 19234
rect 14194 19182 14308 19234
rect 14140 19180 14308 19182
rect 14476 19234 14532 19246
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 14140 19170 14196 19180
rect 13916 18425 13918 18477
rect 13970 18425 13972 18477
rect 13916 18413 13972 18425
rect 12684 17838 12686 17890
rect 12738 17838 12740 17890
rect 12684 17826 12740 17838
rect 14140 17892 14196 17902
rect 11228 17714 11284 17724
rect 11564 17668 11620 17678
rect 13468 17666 13524 17678
rect 11564 17574 11620 17612
rect 12440 17610 12496 17622
rect 12440 17558 12442 17610
rect 12494 17558 12496 17610
rect 12440 17444 12496 17558
rect 12440 17378 12496 17388
rect 13468 17614 13470 17666
rect 13522 17614 13524 17666
rect 10444 16930 10500 16940
rect 12796 17108 12852 17118
rect 12684 16909 12740 16921
rect 12124 16884 12180 16894
rect 12124 16790 12180 16828
rect 12684 16857 12686 16909
rect 12738 16857 12740 16909
rect 10220 16770 10276 16782
rect 10220 16718 10222 16770
rect 10274 16718 10276 16770
rect 10220 15876 10276 16718
rect 11452 16098 11508 16110
rect 11452 16046 11454 16098
rect 11506 16046 11508 16098
rect 10220 15810 10276 15820
rect 10556 15986 10612 15998
rect 10556 15934 10558 15986
rect 10610 15934 10612 15986
rect 10556 15876 10612 15934
rect 11116 15876 11172 15886
rect 10556 15810 10612 15820
rect 10668 15874 11172 15876
rect 10668 15822 11118 15874
rect 11170 15822 11172 15874
rect 10668 15820 11172 15822
rect 10668 15652 10724 15820
rect 11116 15810 11172 15820
rect 10220 15596 10724 15652
rect 10220 15341 10276 15596
rect 10220 15289 10222 15341
rect 10274 15289 10276 15341
rect 10220 15277 10276 15289
rect 11452 15204 11508 16046
rect 11676 16098 11732 16110
rect 11676 16046 11678 16098
rect 11730 16046 11732 16098
rect 11564 15540 11620 15550
rect 11564 15446 11620 15484
rect 11452 14754 11508 15148
rect 11452 14702 11454 14754
rect 11506 14702 11508 14754
rect 11452 14690 11508 14702
rect 8988 14466 9044 14476
rect 10108 14450 10110 14502
rect 10162 14450 10164 14502
rect 10108 14438 10164 14450
rect 11564 14644 11620 14654
rect 8876 13738 8878 13790
rect 8930 13738 8932 13790
rect 9660 13860 9716 13870
rect 9660 13766 9716 13804
rect 8876 13726 8932 13738
rect 11340 13748 11396 13758
rect 8652 13682 8708 13692
rect 8540 13570 8596 13580
rect 8988 13636 9044 13646
rect 8988 13634 9604 13636
rect 8988 13582 8990 13634
rect 9042 13582 9604 13634
rect 8988 13580 9604 13582
rect 8988 13570 9044 13580
rect 9548 13300 9604 13580
rect 9548 13244 9828 13300
rect 8988 13076 9044 13086
rect 8988 12962 9044 13020
rect 9772 13074 9828 13244
rect 9772 13022 9774 13074
rect 9826 13022 9828 13074
rect 9772 13010 9828 13022
rect 8988 12910 8990 12962
rect 9042 12910 9044 12962
rect 8988 12898 9044 12910
rect 9436 12964 9492 12974
rect 8204 12114 8260 12124
rect 9436 12178 9492 12908
rect 9436 12126 9438 12178
rect 9490 12126 9492 12178
rect 9436 12114 9492 12126
rect 10220 12180 10276 12190
rect 10220 12086 10276 12124
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 11340 11618 11396 13692
rect 11564 13746 11620 14588
rect 11564 13694 11566 13746
rect 11618 13694 11620 13746
rect 11564 13682 11620 13694
rect 11676 13636 11732 16046
rect 12552 16042 12608 16054
rect 12552 15990 12554 16042
rect 12606 15990 12608 16042
rect 12552 15652 12608 15990
rect 12552 15586 12608 15596
rect 11676 13074 11732 13580
rect 11676 13022 11678 13074
rect 11730 13022 11732 13074
rect 11676 13010 11732 13022
rect 12012 15540 12068 15550
rect 11340 11566 11342 11618
rect 11394 11566 11396 11618
rect 11340 11554 11396 11566
rect 12012 11366 12068 15484
rect 12684 15540 12740 16857
rect 12796 16322 12852 17052
rect 13244 16996 13300 17006
rect 12796 16270 12798 16322
rect 12850 16270 12852 16322
rect 12796 16258 12852 16270
rect 12908 16884 12964 16894
rect 12684 15474 12740 15484
rect 12908 15314 12964 16828
rect 13244 16100 13300 16940
rect 13468 16884 13524 17614
rect 13468 16818 13524 16828
rect 13580 16658 13636 16670
rect 13580 16606 13582 16658
rect 13634 16606 13636 16658
rect 13580 16548 13636 16606
rect 13580 16482 13636 16492
rect 13468 16100 13524 16110
rect 13244 16098 13524 16100
rect 13244 16046 13470 16098
rect 13522 16046 13524 16098
rect 13244 16044 13524 16046
rect 13468 16034 13524 16044
rect 13468 15876 13524 15886
rect 12908 15262 12910 15314
rect 12962 15262 12964 15314
rect 12908 15250 12964 15262
rect 13244 15314 13300 15326
rect 13244 15262 13246 15314
rect 13298 15262 13300 15314
rect 12740 15092 12796 15102
rect 12348 15090 12796 15092
rect 12348 15038 12742 15090
rect 12794 15038 12796 15090
rect 12348 15036 12796 15038
rect 12124 14420 12180 14430
rect 12124 12292 12180 14364
rect 12348 13746 12404 15036
rect 12740 15026 12796 15036
rect 12348 13694 12350 13746
rect 12402 13694 12404 13746
rect 12348 13682 12404 13694
rect 13132 13860 13188 13870
rect 13132 13746 13188 13804
rect 13132 13694 13134 13746
rect 13186 13694 13188 13746
rect 13132 13682 13188 13694
rect 13244 13748 13300 15262
rect 13468 14868 13524 15820
rect 14140 15764 14196 17836
rect 14344 17668 14400 17678
rect 14344 17574 14400 17612
rect 14476 17108 14532 19182
rect 14924 18506 14980 22204
rect 15372 21812 15428 22878
rect 15372 21746 15428 21756
rect 15708 21812 15764 23102
rect 16156 23156 16212 23166
rect 16156 22594 16212 23100
rect 16828 23156 16884 23166
rect 16828 23154 17556 23156
rect 16828 23102 16830 23154
rect 16882 23102 17556 23154
rect 16828 23100 17556 23102
rect 16828 23090 16884 23100
rect 16492 22932 16548 22942
rect 16156 22542 16158 22594
rect 16210 22542 16212 22594
rect 16156 22530 16212 22542
rect 16268 22930 16548 22932
rect 16268 22878 16494 22930
rect 16546 22878 16548 22930
rect 16268 22876 16548 22878
rect 15708 21746 15764 21756
rect 15932 21700 15988 21710
rect 15708 21140 15764 21150
rect 15596 21028 15652 21038
rect 15260 20692 15316 20702
rect 15260 20690 15428 20692
rect 15260 20638 15262 20690
rect 15314 20638 15428 20690
rect 15260 20636 15428 20638
rect 15260 20626 15316 20636
rect 15036 20132 15316 20188
rect 15036 20066 15092 20076
rect 14588 18450 14644 18462
rect 14588 18398 14590 18450
rect 14642 18398 14644 18450
rect 14924 18454 14926 18506
rect 14978 18454 14980 18506
rect 14924 18442 14980 18454
rect 15036 19234 15092 19246
rect 15036 19182 15038 19234
rect 15090 19182 15092 19234
rect 14588 17890 14644 18398
rect 14924 18340 14980 18350
rect 15036 18340 15092 19182
rect 15260 18450 15316 20132
rect 15372 19684 15428 20636
rect 15372 19618 15428 19628
rect 15260 18398 15262 18450
rect 15314 18398 15316 18450
rect 15260 18386 15316 18398
rect 15372 19178 15428 19190
rect 15372 19126 15374 19178
rect 15426 19126 15428 19178
rect 14924 18338 15092 18340
rect 14924 18286 14926 18338
rect 14978 18286 15092 18338
rect 14924 18284 15092 18286
rect 14924 18274 14980 18284
rect 14588 17838 14590 17890
rect 14642 17838 14644 17890
rect 14588 17826 14644 17838
rect 15372 17892 15428 19126
rect 15596 19066 15652 20972
rect 15708 19908 15764 21084
rect 15932 21140 15988 21644
rect 16156 21588 16212 21598
rect 16268 21588 16324 22876
rect 16492 22866 16548 22876
rect 17500 22930 17556 23100
rect 17500 22878 17502 22930
rect 17554 22878 17556 22930
rect 17500 22866 17556 22878
rect 16156 21586 16324 21588
rect 16156 21534 16158 21586
rect 16210 21534 16324 21586
rect 16156 21532 16324 21534
rect 16940 21586 16996 21598
rect 16940 21534 16942 21586
rect 16994 21534 16996 21586
rect 16156 21522 16212 21532
rect 15932 21074 15988 21084
rect 16940 21140 16996 21534
rect 16940 21074 16996 21084
rect 17612 21586 17668 21598
rect 17612 21534 17614 21586
rect 17666 21534 17668 21586
rect 17612 21028 17668 21534
rect 17612 20962 17668 20972
rect 17164 20804 17220 20814
rect 17164 20802 17668 20804
rect 17164 20750 17166 20802
rect 17218 20750 17668 20802
rect 17164 20748 17668 20750
rect 17164 20738 17220 20748
rect 17612 20242 17668 20748
rect 17836 20580 17892 25116
rect 19180 25284 19236 25294
rect 18060 24610 18116 24622
rect 18060 24558 18062 24610
rect 18114 24558 18116 24610
rect 18060 24052 18116 24558
rect 19180 24164 19236 25228
rect 18844 24108 19236 24164
rect 18060 23986 18116 23996
rect 18620 24052 18676 24062
rect 18620 23958 18676 23996
rect 18844 23940 18900 24108
rect 18788 23908 18900 23940
rect 18788 23856 18790 23908
rect 18842 23884 18900 23908
rect 18956 23940 19012 23950
rect 18842 23856 18844 23884
rect 18788 23844 18844 23856
rect 18956 23846 19012 23884
rect 19404 23940 19460 26014
rect 19516 24162 19572 26852
rect 20188 26740 20244 27022
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20188 26674 20244 26684
rect 19836 26618 20100 26628
rect 20300 26516 20356 27132
rect 20412 27076 20468 27086
rect 20412 26852 20468 27020
rect 20412 26786 20468 26796
rect 20524 26964 20580 27244
rect 20860 27300 20916 28590
rect 20860 27234 20916 27244
rect 21308 28642 21364 28654
rect 21308 28590 21310 28642
rect 21362 28590 21364 28642
rect 21308 27300 21364 28590
rect 22184 28642 22240 29036
rect 22184 28590 22186 28642
rect 22238 28590 22240 28642
rect 22184 28578 22240 28590
rect 22204 28420 22260 28430
rect 21420 27860 21476 27870
rect 21532 27860 21588 27870
rect 21420 27858 21532 27860
rect 21420 27806 21422 27858
rect 21474 27806 21532 27858
rect 21420 27804 21532 27806
rect 21420 27794 21476 27804
rect 21420 27300 21476 27310
rect 21308 27298 21476 27300
rect 21308 27246 21422 27298
rect 21474 27246 21476 27298
rect 21308 27244 21476 27246
rect 21308 27188 21364 27244
rect 21420 27234 21476 27244
rect 21308 27122 21364 27132
rect 20860 27076 20916 27086
rect 20860 26982 20916 27020
rect 20524 26628 20580 26908
rect 21532 26964 21588 27804
rect 22204 27858 22260 28364
rect 22204 27806 22206 27858
rect 22258 27806 22260 27858
rect 22204 27794 22260 27806
rect 22316 27636 22372 29372
rect 22428 29362 22484 29372
rect 22820 29362 22876 29372
rect 21980 27580 22372 27636
rect 22428 28530 22484 28542
rect 22428 28478 22430 28530
rect 22482 28478 22484 28530
rect 20076 26460 20356 26516
rect 20412 26572 20580 26628
rect 21420 26852 21476 26862
rect 19740 26292 19796 26302
rect 20076 26292 20132 26460
rect 19740 26290 20132 26292
rect 19740 26238 19742 26290
rect 19794 26238 20078 26290
rect 20130 26238 20132 26290
rect 20412 26334 20468 26572
rect 20412 26282 20414 26334
rect 20466 26282 20468 26334
rect 20412 26270 20468 26282
rect 20636 26516 20692 26526
rect 19740 26236 20132 26238
rect 19740 26226 19796 26236
rect 20076 26226 20132 26236
rect 20524 26178 20580 26190
rect 20524 26126 20526 26178
rect 20578 26126 20580 26178
rect 20188 25956 20244 25966
rect 20076 25396 20132 25406
rect 20076 25302 20132 25340
rect 20188 25284 20244 25900
rect 20524 25620 20580 26126
rect 20524 25554 20580 25564
rect 20636 25452 20692 26460
rect 20792 26328 20848 26340
rect 20792 26276 20794 26328
rect 20846 26276 20848 26328
rect 20792 25956 20848 26276
rect 20792 25890 20848 25900
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24948 20244 25228
rect 19964 24892 20244 24948
rect 20524 25396 20692 25452
rect 20748 25676 21252 25732
rect 19964 24834 20020 24892
rect 19964 24782 19966 24834
rect 20018 24782 20020 24834
rect 19964 24770 20020 24782
rect 19516 24110 19518 24162
rect 19570 24110 19572 24162
rect 19516 24098 19572 24110
rect 19404 23874 19460 23884
rect 19852 23940 19908 23950
rect 19852 23846 19908 23884
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 17948 23268 18004 23278
rect 20524 23268 20580 25396
rect 20748 25294 20804 25676
rect 20860 25508 20916 25518
rect 20860 25506 21140 25508
rect 20860 25454 20862 25506
rect 20914 25454 21140 25506
rect 20860 25452 21140 25454
rect 20860 25442 20916 25452
rect 20692 25282 20804 25294
rect 20692 25230 20694 25282
rect 20746 25230 20804 25282
rect 20692 25228 20804 25230
rect 20692 25218 20748 25228
rect 21084 23716 21140 25452
rect 21196 25506 21252 25676
rect 21196 25454 21198 25506
rect 21250 25454 21252 25506
rect 21196 25442 21252 25454
rect 21196 23940 21252 23950
rect 21196 23938 21364 23940
rect 21196 23886 21198 23938
rect 21250 23886 21364 23938
rect 21196 23884 21364 23886
rect 21196 23874 21252 23884
rect 21084 23660 21252 23716
rect 21084 23268 21140 23278
rect 20524 23212 20636 23268
rect 17948 21810 18004 23212
rect 20580 23210 20636 23212
rect 20580 23158 20582 23210
rect 20634 23158 20636 23210
rect 21084 23210 21140 23212
rect 20580 23146 20636 23158
rect 20860 23182 20916 23194
rect 20860 23130 20862 23182
rect 20914 23130 20916 23182
rect 21084 23158 21086 23210
rect 21138 23158 21140 23210
rect 21084 23146 21140 23158
rect 21196 23210 21252 23660
rect 21196 23158 21198 23210
rect 21250 23158 21252 23210
rect 21308 23268 21364 23884
rect 21308 23202 21364 23212
rect 21196 23156 21252 23158
rect 20860 23044 20916 23130
rect 21196 23080 21252 23100
rect 21420 23044 21476 26796
rect 21532 26290 21588 26908
rect 21756 27074 21812 27086
rect 21756 27022 21758 27074
rect 21810 27022 21812 27074
rect 21756 26516 21812 27022
rect 21980 26908 22036 27580
rect 22428 27524 22484 28478
rect 23100 28084 23156 32844
rect 23212 30884 23268 32956
rect 23324 30884 23380 30894
rect 23212 30828 23324 30884
rect 23212 29428 23268 29438
rect 23212 29202 23268 29372
rect 23212 29150 23214 29202
rect 23266 29150 23268 29202
rect 23212 28644 23268 29150
rect 23212 28578 23268 28588
rect 23100 28018 23156 28028
rect 23324 27524 23380 30828
rect 22428 27468 22932 27524
rect 22596 27300 22652 27310
rect 22596 27206 22652 27244
rect 22652 27076 22708 27086
rect 21756 26450 21812 26460
rect 21868 26852 22036 26908
rect 22148 26964 22204 27002
rect 22148 26898 22204 26908
rect 21532 26238 21534 26290
rect 21586 26238 21588 26290
rect 21532 26226 21588 26238
rect 21644 26122 21700 26134
rect 21644 26070 21646 26122
rect 21698 26070 21700 26122
rect 21644 24612 21700 26070
rect 21644 24546 21700 24556
rect 21644 23940 21700 23950
rect 21644 23268 21700 23884
rect 21868 23380 21924 26852
rect 22316 26516 22372 26526
rect 22316 26422 22372 26460
rect 22652 26290 22708 27020
rect 22876 27074 22932 27468
rect 22876 27022 22878 27074
rect 22930 27022 22932 27074
rect 22876 27010 22932 27022
rect 22988 27468 23380 27524
rect 22988 26908 23044 27468
rect 23436 27412 23492 33068
rect 24332 32564 24388 32574
rect 24332 32470 24388 32508
rect 24556 32562 24612 32574
rect 24556 32510 24558 32562
rect 24610 32510 24612 32562
rect 23548 32450 23604 32462
rect 23548 32398 23550 32450
rect 23602 32398 23604 32450
rect 23548 31780 23604 32398
rect 23884 31892 23940 31902
rect 24556 31892 24612 32510
rect 24668 32394 24724 33068
rect 25228 33068 25396 33124
rect 26572 33346 26628 33358
rect 26572 33294 26574 33346
rect 26626 33294 26628 33346
rect 26572 33124 26628 33294
rect 27448 33348 27504 33358
rect 27448 33254 27504 33292
rect 25004 33012 25060 33022
rect 24668 32342 24670 32394
rect 24722 32342 24724 32394
rect 24668 32330 24724 32342
rect 24892 32564 24948 32574
rect 23884 31890 24612 31892
rect 23884 31838 23886 31890
rect 23938 31838 24612 31890
rect 23884 31836 24612 31838
rect 24724 31892 24780 31902
rect 23884 31826 23940 31836
rect 24724 31798 24780 31836
rect 23548 31714 23604 31724
rect 23884 30212 23940 30222
rect 24220 30212 24276 30222
rect 23884 30118 23940 30156
rect 23996 30210 24276 30212
rect 23996 30158 24222 30210
rect 24274 30158 24276 30210
rect 23996 30156 24276 30158
rect 24892 30212 24948 32508
rect 25004 31722 25060 32956
rect 25228 32562 25284 33068
rect 26572 33058 26628 33068
rect 25228 32510 25230 32562
rect 25282 32510 25284 32562
rect 25228 32498 25284 32510
rect 25396 32730 25452 32742
rect 25396 32678 25398 32730
rect 25450 32678 25452 32730
rect 25396 32564 25452 32678
rect 25676 32564 25732 32574
rect 25396 32562 25732 32564
rect 25396 32510 25678 32562
rect 25730 32510 25732 32562
rect 25396 32508 25732 32510
rect 25676 32498 25732 32508
rect 26460 32452 26516 32462
rect 26460 32358 26516 32396
rect 27580 32116 27636 36876
rect 29036 36820 29092 37100
rect 29036 36764 29988 36820
rect 29932 36706 29988 36764
rect 29932 36654 29934 36706
rect 29986 36654 29988 36706
rect 29932 36642 29988 36654
rect 29036 36482 29092 36494
rect 27784 36426 27840 36438
rect 27784 36374 27786 36426
rect 27838 36374 27840 36426
rect 29036 36430 29038 36482
rect 29090 36430 29092 36482
rect 27784 35812 27840 36374
rect 28028 36372 28084 36382
rect 27916 36370 28084 36372
rect 27916 36318 28030 36370
rect 28082 36318 28084 36370
rect 27916 36316 28084 36318
rect 27784 35756 27860 35812
rect 27692 35700 27748 35710
rect 27692 35606 27748 35644
rect 27692 33572 27748 33582
rect 27804 33572 27860 35756
rect 27916 35588 27972 36316
rect 28028 36306 28084 36316
rect 29036 35812 29092 36430
rect 30268 36484 30324 36494
rect 30268 36390 30324 36428
rect 29036 35746 29092 35756
rect 29372 36258 29428 36270
rect 29372 36206 29374 36258
rect 29426 36206 29428 36258
rect 29372 35700 29428 36206
rect 29596 36148 29652 36158
rect 29596 35810 29652 36092
rect 29596 35758 29598 35810
rect 29650 35758 29652 35810
rect 29596 35746 29652 35758
rect 29372 35634 29428 35644
rect 27916 35522 27972 35532
rect 30268 35588 30324 35598
rect 27972 35364 28028 35374
rect 27972 35026 28028 35308
rect 27972 34974 27974 35026
rect 28026 34974 28028 35026
rect 27972 34962 28028 34974
rect 27692 33570 27860 33572
rect 27692 33518 27694 33570
rect 27746 33518 27860 33570
rect 27692 33516 27860 33518
rect 28028 34804 28084 34814
rect 27692 33506 27748 33516
rect 27580 32060 27748 32116
rect 27692 31892 27748 32060
rect 27692 31826 27748 31836
rect 27916 31892 27972 31902
rect 27916 31798 27972 31836
rect 25452 31780 25508 31790
rect 25788 31780 25844 31790
rect 25004 31670 25006 31722
rect 25058 31670 25060 31722
rect 25004 31444 25060 31670
rect 25004 31378 25060 31388
rect 25228 31722 25284 31734
rect 25228 31670 25230 31722
rect 25282 31670 25284 31722
rect 25452 31698 25454 31724
rect 25506 31698 25508 31724
rect 25620 31762 25732 31780
rect 25620 31710 25622 31762
rect 25674 31710 25732 31762
rect 25620 31698 25732 31710
rect 25452 31686 25508 31698
rect 25228 30884 25284 31670
rect 25564 31332 25620 31342
rect 25228 30818 25284 30828
rect 25452 30994 25508 31006
rect 25452 30942 25454 30994
rect 25506 30942 25508 30994
rect 25452 30884 25508 30942
rect 25452 30818 25508 30828
rect 25564 30222 25620 31276
rect 25676 30436 25732 31698
rect 25788 30994 25844 31724
rect 27804 31780 27860 31790
rect 26012 31668 26068 31678
rect 26012 31574 26068 31612
rect 26236 31556 26292 31566
rect 25788 30942 25790 30994
rect 25842 30942 25844 30994
rect 25788 30930 25844 30942
rect 26124 31021 26180 31033
rect 26124 30969 26126 31021
rect 26178 30969 26180 31021
rect 26124 30772 26180 30969
rect 26236 30882 26292 31500
rect 27244 31444 27300 31454
rect 27244 31033 27300 31388
rect 26460 30996 26516 31006
rect 26460 30994 26628 30996
rect 26460 30942 26462 30994
rect 26514 30942 26628 30994
rect 26460 30940 26628 30942
rect 26460 30930 26516 30940
rect 26236 30830 26238 30882
rect 26290 30830 26292 30882
rect 26236 30818 26292 30830
rect 26124 30706 26180 30716
rect 26348 30772 26404 30782
rect 25676 30380 25844 30436
rect 25004 30212 25060 30222
rect 24892 30210 25060 30212
rect 24892 30158 25006 30210
rect 25058 30158 25060 30210
rect 24892 30156 25060 30158
rect 23548 29988 23604 29998
rect 23548 29426 23604 29932
rect 23548 29374 23550 29426
rect 23602 29374 23604 29426
rect 23548 28756 23604 29374
rect 23884 29204 23940 29214
rect 23884 29110 23940 29148
rect 23548 28700 23940 28756
rect 23660 28532 23716 28542
rect 23100 27356 23492 27412
rect 23548 28420 23604 28430
rect 23100 27074 23156 27356
rect 23100 27022 23102 27074
rect 23154 27022 23156 27074
rect 23100 27010 23156 27022
rect 23548 26908 23604 28364
rect 23660 27186 23716 28476
rect 23660 27134 23662 27186
rect 23714 27134 23716 27186
rect 23660 27122 23716 27134
rect 23772 28418 23828 28430
rect 23772 28366 23774 28418
rect 23826 28366 23828 28418
rect 23772 27972 23828 28366
rect 23772 27076 23828 27916
rect 23772 27010 23828 27020
rect 23884 26908 23940 28700
rect 23996 27972 24052 30156
rect 24220 30146 24276 30156
rect 25004 30100 25060 30156
rect 25228 30212 25284 30222
rect 25228 30118 25284 30156
rect 25508 30210 25620 30222
rect 25508 30158 25510 30210
rect 25562 30158 25620 30210
rect 25508 30156 25620 30158
rect 25788 30212 25844 30380
rect 25508 30146 25564 30156
rect 24556 29988 24612 29998
rect 24556 29894 24612 29932
rect 24220 29428 24276 29466
rect 24220 29362 24276 29372
rect 24220 29204 24276 29214
rect 24108 28644 24164 28654
rect 24108 28550 24164 28588
rect 24220 28644 24276 29148
rect 25004 28868 25060 30044
rect 25788 29652 25844 30156
rect 26348 30210 26404 30716
rect 26348 30158 26350 30210
rect 26402 30158 26404 30210
rect 26348 30146 26404 30158
rect 26460 30212 26516 30222
rect 25900 29652 25956 29662
rect 25788 29650 25956 29652
rect 25788 29598 25902 29650
rect 25954 29598 25956 29650
rect 25788 29596 25956 29598
rect 25900 29586 25956 29596
rect 25564 29426 25620 29438
rect 25564 29374 25566 29426
rect 25618 29374 25620 29426
rect 25004 28802 25060 28812
rect 25116 29316 25172 29326
rect 24444 28644 24500 28654
rect 24556 28644 24612 28654
rect 24220 28642 24388 28644
rect 24220 28590 24222 28642
rect 24274 28590 24388 28642
rect 24220 28588 24388 28590
rect 24220 28578 24276 28588
rect 24108 27972 24164 27982
rect 23996 27970 24164 27972
rect 23996 27918 24110 27970
rect 24162 27918 24164 27970
rect 23996 27916 24164 27918
rect 24108 27906 24164 27916
rect 22988 26852 23156 26908
rect 23548 26852 23716 26908
rect 23884 26852 24276 26908
rect 22652 26238 22654 26290
rect 22706 26238 22708 26290
rect 22652 26226 22708 26238
rect 23100 26292 23156 26852
rect 23100 26198 23156 26236
rect 22932 26066 22988 26078
rect 22932 26014 22934 26066
rect 22986 26014 22988 26066
rect 22932 25844 22988 26014
rect 22092 25788 22988 25844
rect 21980 25620 22036 25630
rect 21980 25526 22036 25564
rect 21980 24052 22036 24062
rect 22092 24052 22148 25788
rect 23548 24612 23604 24622
rect 21980 24050 22148 24052
rect 21980 23998 21982 24050
rect 22034 23998 22148 24050
rect 21980 23996 22148 23998
rect 22204 24498 22260 24510
rect 22204 24446 22206 24498
rect 22258 24446 22260 24498
rect 21980 23986 22036 23996
rect 21868 23314 21924 23324
rect 20860 22978 20916 22988
rect 21308 22988 21476 23044
rect 21532 23044 21588 23054
rect 17948 21758 17950 21810
rect 18002 21758 18004 21810
rect 17948 21746 18004 21758
rect 18284 22930 18340 22942
rect 18284 22878 18286 22930
rect 18338 22878 18340 22930
rect 17948 21140 18004 21150
rect 17948 20802 18004 21084
rect 18284 21038 18340 22878
rect 20356 22930 20412 22942
rect 20356 22878 20358 22930
rect 20410 22878 20412 22930
rect 19628 22820 19684 22830
rect 19628 22594 19684 22764
rect 19628 22542 19630 22594
rect 19682 22542 19684 22594
rect 19628 22530 19684 22542
rect 19871 22820 19927 22830
rect 19871 22370 19927 22764
rect 20356 22820 20412 22878
rect 20356 22754 20412 22764
rect 19871 22318 19873 22370
rect 19925 22318 19927 22370
rect 19871 22306 19927 22318
rect 20748 22372 20804 22382
rect 20748 22278 20804 22316
rect 21084 22372 21140 22382
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 18396 21812 18452 21822
rect 18396 21586 18452 21756
rect 19292 21812 19348 21822
rect 19292 21718 19348 21756
rect 19628 21812 19684 21822
rect 18396 21534 18398 21586
rect 18450 21534 18452 21586
rect 18396 21522 18452 21534
rect 19628 21586 19684 21756
rect 19628 21534 19630 21586
rect 19682 21534 19684 21586
rect 19628 21522 19684 21534
rect 20207 21586 20263 21598
rect 20207 21534 20209 21586
rect 20261 21534 20263 21586
rect 18266 21026 18340 21038
rect 18266 20974 18268 21026
rect 18320 20974 18340 21026
rect 18266 20972 18340 20974
rect 18732 21362 18788 21374
rect 18732 21310 18734 21362
rect 18786 21310 18788 21362
rect 18266 20962 18322 20972
rect 17948 20750 17950 20802
rect 18002 20750 18004 20802
rect 17948 20738 18004 20750
rect 18508 20802 18564 20814
rect 18508 20750 18510 20802
rect 18562 20750 18564 20802
rect 18508 20580 18564 20750
rect 17836 20524 18004 20580
rect 17612 20190 17614 20242
rect 17666 20190 17668 20242
rect 17612 20178 17668 20190
rect 15820 20132 15876 20142
rect 15820 20038 15876 20076
rect 16492 20018 16548 20030
rect 15988 19962 16044 19974
rect 15988 19910 15990 19962
rect 16042 19910 16044 19962
rect 15708 19852 15876 19908
rect 15708 19348 15764 19358
rect 15708 19234 15764 19292
rect 15708 19182 15710 19234
rect 15762 19182 15764 19234
rect 15708 19170 15764 19182
rect 15596 19014 15598 19066
rect 15650 19014 15652 19066
rect 15596 19002 15652 19014
rect 15372 17826 15428 17836
rect 14476 17042 14532 17052
rect 15820 17666 15876 19852
rect 15988 19684 16044 19910
rect 15988 19618 16044 19628
rect 16492 19966 16494 20018
rect 16546 19966 16548 20018
rect 15820 17614 15822 17666
rect 15874 17614 15876 17666
rect 14344 16100 14400 16110
rect 14344 16006 14400 16044
rect 15372 16100 15428 16110
rect 15820 16100 15876 17614
rect 15372 16098 15876 16100
rect 15372 16046 15374 16098
rect 15426 16046 15876 16098
rect 15372 16044 15876 16046
rect 15932 19012 15988 19022
rect 15932 17108 15988 18956
rect 16492 19012 16548 19966
rect 16734 20020 16790 20030
rect 16734 19926 16790 19964
rect 17276 20020 17332 20030
rect 17276 19926 17332 19964
rect 16492 18946 16548 18956
rect 17108 19012 17164 19022
rect 17108 18918 17164 18956
rect 16940 18452 16996 18462
rect 17482 18452 17538 18462
rect 16940 18450 17538 18452
rect 16940 18398 16942 18450
rect 16994 18398 17484 18450
rect 17536 18398 17538 18450
rect 16940 18396 17538 18398
rect 16940 18386 16996 18396
rect 17482 18386 17538 18396
rect 17724 18450 17780 18462
rect 17724 18398 17726 18450
rect 17778 18398 17780 18450
rect 16604 18228 16660 18238
rect 16268 18226 16660 18228
rect 16268 18174 16606 18226
rect 16658 18174 16660 18226
rect 16268 18172 16660 18174
rect 16100 17108 16156 17118
rect 15932 17106 16156 17108
rect 15932 17054 16102 17106
rect 16154 17054 16156 17106
rect 15932 17052 16156 17054
rect 15372 16034 15428 16044
rect 14588 15988 14644 15998
rect 13580 15708 14196 15764
rect 14476 15986 14644 15988
rect 14476 15934 14590 15986
rect 14642 15934 14644 15986
rect 14476 15932 14644 15934
rect 13580 15202 13636 15708
rect 14476 15652 14532 15932
rect 14588 15922 14644 15932
rect 13916 15596 14532 15652
rect 13580 15150 13582 15202
rect 13634 15150 13636 15202
rect 13580 15138 13636 15150
rect 13692 15353 13748 15365
rect 13692 15301 13694 15353
rect 13746 15301 13748 15353
rect 13692 14980 13748 15301
rect 13916 15314 13972 15596
rect 13916 15262 13918 15314
rect 13970 15262 13972 15314
rect 13916 15250 13972 15262
rect 14252 15314 14308 15326
rect 14252 15262 14254 15314
rect 14306 15262 14308 15314
rect 14252 15148 14308 15262
rect 14812 15316 14868 15326
rect 15484 15316 15540 15326
rect 15932 15316 15988 17052
rect 16100 17042 16156 17052
rect 16156 16212 16212 16222
rect 16268 16212 16324 18172
rect 16604 18162 16660 18172
rect 17724 18116 17780 18398
rect 17780 18060 17892 18116
rect 17724 18050 17780 18060
rect 16604 17666 16660 17678
rect 16604 17614 16606 17666
rect 16658 17614 16660 17666
rect 16604 17106 16660 17614
rect 16604 17054 16606 17106
rect 16658 17054 16660 17106
rect 16604 17042 16660 17054
rect 16940 16884 16996 16894
rect 17482 16884 17538 16894
rect 16940 16882 17538 16884
rect 16940 16830 16942 16882
rect 16994 16830 17484 16882
rect 17536 16830 17538 16882
rect 16940 16828 17538 16830
rect 16940 16818 16996 16828
rect 17482 16818 17538 16828
rect 17724 16884 17780 16894
rect 17724 16790 17780 16828
rect 16156 16210 16324 16212
rect 16156 16158 16158 16210
rect 16210 16158 16324 16210
rect 16156 16156 16324 16158
rect 16156 16146 16212 16156
rect 15484 15314 15988 15316
rect 14812 15222 14868 15260
rect 14980 15258 15036 15270
rect 13692 14914 13748 14924
rect 14140 15092 14308 15148
rect 14980 15206 14982 15258
rect 15034 15206 15036 15258
rect 15484 15262 15486 15314
rect 15538 15262 15988 15314
rect 15484 15260 15988 15262
rect 16492 15316 16548 15326
rect 15484 15250 15540 15260
rect 13468 14802 13524 14812
rect 13468 14532 13524 14542
rect 13468 14438 13524 14476
rect 14140 13860 14196 15092
rect 14588 14980 14644 14990
rect 14588 14754 14644 14924
rect 14980 14756 15036 15206
rect 15726 15092 15782 15102
rect 14588 14702 14590 14754
rect 14642 14702 14644 14754
rect 14588 14690 14644 14702
rect 14700 14700 15036 14756
rect 15708 15090 15782 15092
rect 15708 15038 15728 15090
rect 15780 15038 15782 15090
rect 15708 15026 15782 15038
rect 16156 15092 16212 15102
rect 14344 14474 14400 14486
rect 14344 14422 14346 14474
rect 14398 14422 14400 14474
rect 14344 14420 14400 14422
rect 14344 14354 14400 14364
rect 14252 13860 14308 13870
rect 14140 13858 14308 13860
rect 14140 13806 14254 13858
rect 14306 13806 14308 13858
rect 14140 13804 14308 13806
rect 14252 13794 14308 13804
rect 13244 13682 13300 13692
rect 13804 13748 13860 13758
rect 13468 13300 13524 13310
rect 13468 12852 13524 13244
rect 13448 12796 13524 12852
rect 12124 12290 12628 12292
rect 12124 12238 12126 12290
rect 12178 12238 12628 12290
rect 12124 12236 12628 12238
rect 12124 12226 12180 12236
rect 12572 12178 12628 12236
rect 12572 12126 12574 12178
rect 12626 12126 12628 12178
rect 13448 12234 13504 12796
rect 13448 12182 13450 12234
rect 13502 12182 13504 12234
rect 13692 12292 13748 12302
rect 13804 12292 13860 13692
rect 14008 13746 14064 13758
rect 14008 13694 14010 13746
rect 14062 13694 14064 13746
rect 14008 13636 14064 13694
rect 14700 13636 14756 14700
rect 15596 14532 15652 14542
rect 15596 14438 15652 14476
rect 15708 14308 15764 15026
rect 15932 14644 15988 14654
rect 15932 14530 15988 14588
rect 15932 14478 15934 14530
rect 15986 14478 15988 14530
rect 15932 14466 15988 14478
rect 16044 14532 16100 14542
rect 15708 14242 15764 14252
rect 15596 13748 15652 13758
rect 15914 13748 15970 13758
rect 15596 13746 15970 13748
rect 15596 13694 15598 13746
rect 15650 13694 15916 13746
rect 15968 13694 15970 13746
rect 15596 13692 15970 13694
rect 15596 13682 15652 13692
rect 15914 13682 15970 13692
rect 16044 13748 16100 14476
rect 16044 13682 16100 13692
rect 16156 13746 16212 15036
rect 16492 13914 16548 15260
rect 16940 15316 16996 15326
rect 17482 15316 17538 15326
rect 16940 15314 17538 15316
rect 16940 15262 16942 15314
rect 16994 15262 17484 15314
rect 17536 15262 17538 15314
rect 16940 15260 17538 15262
rect 16940 15250 16996 15260
rect 17482 15250 17538 15260
rect 17724 15316 17780 15326
rect 17836 15316 17892 18060
rect 17724 15314 17892 15316
rect 17724 15262 17726 15314
rect 17778 15262 17892 15314
rect 17724 15260 17892 15262
rect 17724 15250 17780 15260
rect 16604 15090 16660 15102
rect 16604 15038 16606 15090
rect 16658 15038 16660 15090
rect 16604 14644 16660 15038
rect 16828 14644 16884 14654
rect 16604 14642 16884 14644
rect 16604 14590 16830 14642
rect 16882 14590 16884 14642
rect 16604 14588 16884 14590
rect 16828 14578 16884 14588
rect 16492 13862 16494 13914
rect 16546 13862 16548 13914
rect 16492 13850 16548 13862
rect 17164 14308 17220 14318
rect 16156 13694 16158 13746
rect 16210 13694 16212 13746
rect 17052 13748 17108 13758
rect 16156 13682 16212 13694
rect 16660 13690 16716 13702
rect 14008 13580 14756 13636
rect 16660 13638 16662 13690
rect 16714 13638 16716 13690
rect 13692 12290 13860 12292
rect 13692 12238 13694 12290
rect 13746 12238 13860 12290
rect 13692 12236 13860 12238
rect 14252 12290 14308 13580
rect 15260 13524 15316 13534
rect 16660 13524 16716 13638
rect 15260 13522 16436 13524
rect 15260 13470 15262 13522
rect 15314 13470 16436 13522
rect 15260 13468 16436 13470
rect 15260 13458 15316 13468
rect 14476 13412 14532 13422
rect 14476 13074 14532 13356
rect 14476 13022 14478 13074
rect 14530 13022 14532 13074
rect 14476 13010 14532 13022
rect 16380 13074 16436 13468
rect 16660 13458 16716 13468
rect 16380 13022 16382 13074
rect 16434 13022 16436 13074
rect 16380 13010 16436 13022
rect 14252 12238 14254 12290
rect 14306 12238 14308 12290
rect 13692 12226 13748 12236
rect 14252 12226 14308 12238
rect 17052 12964 17108 13692
rect 17164 13524 17220 14252
rect 17276 13748 17332 13758
rect 17276 13654 17332 13692
rect 17164 13468 17332 13524
rect 17164 12964 17220 12974
rect 17052 12962 17220 12964
rect 17052 12910 17166 12962
rect 17218 12910 17220 12962
rect 17052 12908 17220 12910
rect 13448 12170 13504 12182
rect 16156 12180 16212 12190
rect 12572 12114 12628 12126
rect 16156 12086 16212 12124
rect 16940 12180 16996 12190
rect 17052 12180 17108 12908
rect 17164 12898 17220 12908
rect 17276 12962 17332 13468
rect 17276 12910 17278 12962
rect 17330 12910 17332 12962
rect 17276 12898 17332 12910
rect 16940 12178 17108 12180
rect 16940 12126 16942 12178
rect 16994 12126 17108 12178
rect 16940 12124 17108 12126
rect 17612 12738 17668 12750
rect 17612 12686 17614 12738
rect 17666 12686 17668 12738
rect 17612 12180 17668 12686
rect 16940 12114 16996 12124
rect 17612 12114 17668 12124
rect 17948 11620 18004 20524
rect 18508 20514 18564 20524
rect 18396 20132 18452 20142
rect 18396 18562 18452 20076
rect 18732 20020 18788 21310
rect 19012 21364 19068 21374
rect 19964 21364 20020 21374
rect 19012 20858 19068 21308
rect 19012 20806 19014 20858
rect 19066 20806 19068 20858
rect 19012 20794 19068 20806
rect 19516 21362 20020 21364
rect 19516 21310 19966 21362
rect 20018 21310 20020 21362
rect 19516 21308 20020 21310
rect 19180 20690 19236 20702
rect 19180 20638 19182 20690
rect 19234 20638 19236 20690
rect 19180 20244 19236 20638
rect 19180 20178 19236 20188
rect 19292 20580 19348 20590
rect 19180 20020 19236 20030
rect 18732 20018 19236 20020
rect 18732 19966 19182 20018
rect 19234 19966 19236 20018
rect 18732 19964 19236 19966
rect 18396 18510 18398 18562
rect 18450 18510 18452 18562
rect 18228 18394 18284 18406
rect 18228 18342 18230 18394
rect 18282 18342 18284 18394
rect 18228 17892 18284 18342
rect 18060 17836 18284 17892
rect 18396 17892 18452 18510
rect 19068 18452 19124 19964
rect 19180 19954 19236 19964
rect 19068 18450 19236 18452
rect 19068 18398 19070 18450
rect 19122 18398 19236 18450
rect 19068 18396 19236 18398
rect 19068 18386 19124 18396
rect 18900 18338 18956 18350
rect 18900 18286 18902 18338
rect 18954 18286 18956 18338
rect 18900 18116 18956 18286
rect 18900 18050 18956 18060
rect 19068 17892 19124 17902
rect 18396 17890 19124 17892
rect 18396 17838 19070 17890
rect 19122 17838 19124 17890
rect 18396 17836 19124 17838
rect 18060 16100 18116 17836
rect 18172 17668 18228 17678
rect 18172 17332 18228 17612
rect 18172 17276 18284 17332
rect 18228 16938 18284 17276
rect 18228 16886 18230 16938
rect 18282 16886 18284 16938
rect 18396 16994 18452 17836
rect 19068 17826 19124 17836
rect 18508 17668 18564 17678
rect 18508 17574 18564 17612
rect 18396 16942 18398 16994
rect 18450 16942 18452 16994
rect 18396 16930 18452 16942
rect 18228 16874 18284 16886
rect 18956 16884 19012 16894
rect 18060 16006 18116 16044
rect 18228 15540 18284 15550
rect 18228 15370 18284 15484
rect 18228 15318 18230 15370
rect 18282 15318 18284 15370
rect 18732 15540 18788 15550
rect 18228 15306 18284 15318
rect 18396 15316 18452 15326
rect 18396 15222 18452 15260
rect 18060 15204 18116 15214
rect 18060 13746 18116 15148
rect 18060 13694 18062 13746
rect 18114 13694 18116 13746
rect 18060 13682 18116 13694
rect 18172 15092 18228 15102
rect 18172 13086 18228 15036
rect 18732 14642 18788 15484
rect 18844 15204 18900 15242
rect 18844 15138 18900 15148
rect 18956 14980 19012 16828
rect 19180 16884 19236 18396
rect 19180 16818 19236 16828
rect 18956 14914 19012 14924
rect 19180 15314 19236 15326
rect 19180 15262 19182 15314
rect 19234 15262 19236 15314
rect 19180 14868 19236 15262
rect 19292 15204 19348 20524
rect 19404 17668 19460 17678
rect 19404 17574 19460 17612
rect 19516 17444 19572 21308
rect 19964 21298 20020 21308
rect 20207 21028 20263 21534
rect 21084 21586 21140 22316
rect 21084 21534 21086 21586
rect 21138 21534 21140 21586
rect 21084 21522 21140 21534
rect 21308 21588 21364 22988
rect 21308 21252 21364 21532
rect 20207 20962 20263 20972
rect 21084 21196 21364 21252
rect 20860 20916 20916 20926
rect 20860 20802 20916 20860
rect 20860 20750 20862 20802
rect 20914 20750 20916 20802
rect 20860 20738 20916 20750
rect 19684 20580 19740 20590
rect 19684 20486 19740 20524
rect 20524 20578 20580 20590
rect 20524 20526 20526 20578
rect 20578 20526 20580 20578
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19964 20244 20020 20254
rect 19964 20018 20020 20188
rect 20524 20244 20580 20526
rect 20524 20178 20580 20188
rect 19964 19966 19966 20018
rect 20018 19966 20020 20018
rect 19964 19954 20020 19966
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19852 18564 19908 18574
rect 19852 18450 19908 18508
rect 19852 18398 19854 18450
rect 19906 18398 19908 18450
rect 19852 18386 19908 18398
rect 19292 15138 19348 15148
rect 19404 17388 19572 17444
rect 19628 18116 19684 18126
rect 21084 18116 21140 21196
rect 21402 20916 21458 20926
rect 21402 20822 21458 20860
rect 21532 20580 21588 22988
rect 21644 22372 21700 23212
rect 21756 23156 21812 23166
rect 21756 23062 21812 23100
rect 22204 22372 22260 24446
rect 22652 23604 22708 23614
rect 22652 22594 22708 23548
rect 22652 22542 22654 22594
rect 22706 22542 22708 22594
rect 22652 22530 22708 22542
rect 22316 22372 22372 22382
rect 22204 22370 22372 22372
rect 22204 22318 22318 22370
rect 22370 22318 22372 22370
rect 22204 22316 22372 22318
rect 21644 22306 21700 22316
rect 22316 22306 22372 22316
rect 23548 22342 23604 24556
rect 23548 22290 23550 22342
rect 23602 22290 23604 22342
rect 23548 22278 23604 22290
rect 21868 21252 21924 21262
rect 21644 20916 21700 20926
rect 21644 20802 21700 20860
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20738 21700 20750
rect 21756 20804 21812 20814
rect 21532 20524 21700 20580
rect 21476 19236 21532 19246
rect 21476 19142 21532 19180
rect 21308 19124 21364 19134
rect 21308 19030 21364 19068
rect 19180 14812 19330 14868
rect 19274 14754 19330 14812
rect 19274 14702 19276 14754
rect 19328 14702 19330 14754
rect 19274 14690 19330 14702
rect 18732 14590 18734 14642
rect 18786 14590 18788 14642
rect 18732 14578 18788 14590
rect 18172 13074 18284 13086
rect 18172 13022 18230 13074
rect 18282 13022 18284 13074
rect 18172 13020 18284 13022
rect 18228 13010 18284 13020
rect 19404 12205 19460 17388
rect 19516 15874 19572 15886
rect 19516 15822 19518 15874
rect 19570 15822 19572 15874
rect 19516 15428 19572 15822
rect 19516 15362 19572 15372
rect 19628 15214 19684 18060
rect 20748 18060 21140 18116
rect 20524 17442 20580 17454
rect 20524 17390 20526 17442
rect 20578 17390 20580 17442
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 19740 16884 19796 16894
rect 19740 16790 19796 16828
rect 19852 16098 19908 17052
rect 20524 16882 20580 17390
rect 20524 16830 20526 16882
rect 20578 16830 20580 16882
rect 20524 16818 20580 16830
rect 19852 16046 19854 16098
rect 19906 16046 19908 16098
rect 19852 16034 19908 16046
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19572 15202 19684 15214
rect 19572 15150 19574 15202
rect 19626 15150 19684 15202
rect 19572 15148 19684 15150
rect 19852 15316 19908 15326
rect 19572 15138 19628 15148
rect 19516 14980 19572 14990
rect 19516 14530 19572 14924
rect 19516 14478 19518 14530
rect 19570 14478 19572 14530
rect 19516 14466 19572 14478
rect 19628 14420 19684 14430
rect 19628 13972 19684 14364
rect 19852 14362 19908 15260
rect 19852 14310 19854 14362
rect 19906 14310 19908 14362
rect 20020 14474 20076 14486
rect 20020 14422 20022 14474
rect 20074 14422 20076 14474
rect 20020 14420 20076 14422
rect 20020 14354 20076 14364
rect 19852 14298 19908 14310
rect 20300 14308 20356 14318
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13916 20020 13972
rect 19964 13858 20020 13916
rect 19964 13806 19966 13858
rect 20018 13806 20020 13858
rect 19964 13794 20020 13806
rect 20300 12962 20356 14252
rect 20300 12910 20302 12962
rect 20354 12910 20356 12962
rect 20300 12898 20356 12910
rect 19964 12740 20020 12750
rect 19964 12738 20244 12740
rect 19964 12686 19966 12738
rect 20018 12686 20244 12738
rect 19964 12684 20244 12686
rect 19964 12674 20020 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20188 12404 20244 12684
rect 18732 12193 18788 12205
rect 18396 12178 18452 12190
rect 18732 12180 18734 12193
rect 18396 12126 18398 12178
rect 18450 12126 18452 12178
rect 17948 11564 18116 11620
rect 17948 11396 18004 11406
rect 12012 11314 12014 11366
rect 12066 11314 12068 11366
rect 12012 11302 12068 11314
rect 16828 11394 18004 11396
rect 16828 11342 17950 11394
rect 18002 11342 18004 11394
rect 16828 11340 18004 11342
rect 14028 11172 14084 11182
rect 14028 10610 14084 11116
rect 14028 10558 14030 10610
rect 14082 10558 14084 10610
rect 14028 10546 14084 10558
rect 16716 10612 16772 10622
rect 16716 10518 16772 10556
rect 14812 10500 14868 10510
rect 14812 10406 14868 10444
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 16828 9278 16884 11340
rect 17948 11330 18004 11340
rect 17108 11172 17164 11182
rect 17108 11078 17164 11116
rect 18060 11172 18116 11564
rect 18396 11508 18452 12126
rect 18620 12141 18734 12180
rect 18786 12141 18788 12193
rect 19404 12153 19406 12205
rect 19458 12153 19460 12205
rect 19404 12141 19460 12153
rect 20076 12348 20244 12404
rect 20748 12404 20804 18060
rect 21532 17780 21588 17790
rect 21644 17780 21700 20524
rect 21756 19236 21812 20748
rect 21868 20130 21924 21196
rect 22148 21252 22204 21262
rect 22148 20858 22204 21196
rect 22148 20806 22150 20858
rect 22202 20806 22204 20858
rect 22820 20916 22876 20926
rect 22820 20822 22876 20860
rect 22148 20794 22204 20806
rect 22316 20692 22372 20702
rect 21868 20078 21870 20130
rect 21922 20078 21924 20130
rect 21868 20066 21924 20078
rect 22092 20690 22372 20692
rect 22092 20638 22318 20690
rect 22370 20638 22372 20690
rect 22092 20636 22372 20638
rect 21756 18562 21812 19180
rect 21980 19348 22036 19358
rect 21980 19234 22036 19292
rect 21980 19182 21982 19234
rect 22034 19182 22036 19234
rect 21980 19170 22036 19182
rect 22092 19124 22148 20636
rect 22316 20626 22372 20636
rect 22204 20018 22260 20030
rect 22204 19966 22206 20018
rect 22258 19966 22260 20018
rect 22204 19470 22260 19966
rect 22540 19794 22596 19806
rect 22540 19742 22542 19794
rect 22594 19742 22596 19794
rect 22204 19458 22278 19470
rect 22204 19406 22224 19458
rect 22276 19406 22278 19458
rect 22204 19404 22278 19406
rect 22222 19394 22278 19404
rect 22204 19124 22260 19134
rect 22092 19068 22204 19124
rect 21756 18510 21758 18562
rect 21810 18510 21812 18562
rect 21756 18498 21812 18510
rect 22204 18450 22260 19068
rect 22540 18564 22596 19742
rect 23492 19796 23548 19806
rect 22820 19348 22876 19358
rect 22820 19254 22876 19292
rect 23492 19346 23548 19740
rect 23660 19684 23716 26852
rect 23884 26740 23940 26750
rect 23772 26292 23828 26302
rect 23772 25172 23828 26236
rect 23884 25618 23940 26684
rect 23884 25566 23886 25618
rect 23938 25566 23940 25618
rect 23884 25554 23940 25566
rect 23772 25116 23940 25172
rect 23772 24749 23828 24761
rect 23772 24697 23774 24749
rect 23826 24697 23828 24749
rect 23772 22596 23828 24697
rect 23884 24050 23940 25116
rect 23884 23998 23886 24050
rect 23938 23998 23940 24050
rect 23884 23986 23940 23998
rect 23996 24500 24052 24510
rect 23996 23181 24052 24444
rect 24220 23492 24276 26852
rect 24332 24724 24388 28588
rect 24500 28642 24612 28644
rect 24500 28590 24558 28642
rect 24610 28590 24612 28642
rect 24500 28588 24612 28590
rect 24444 26908 24500 28588
rect 24556 28578 24612 28588
rect 24724 27860 24780 27870
rect 24724 27766 24780 27804
rect 25116 27412 25172 29260
rect 25564 28868 25620 29374
rect 25564 28802 25620 28812
rect 25900 28868 25956 28878
rect 25900 28866 26404 28868
rect 25900 28814 25902 28866
rect 25954 28814 26404 28866
rect 25900 28812 26404 28814
rect 25900 28802 25956 28812
rect 25564 28644 25620 28654
rect 25564 28642 25732 28644
rect 25564 28590 25566 28642
rect 25618 28590 25732 28642
rect 25564 28588 25732 28590
rect 25564 28578 25620 28588
rect 25228 28420 25284 28430
rect 25228 28418 25508 28420
rect 25228 28366 25230 28418
rect 25282 28366 25508 28418
rect 25228 28364 25508 28366
rect 25228 28354 25284 28364
rect 25116 27346 25172 27356
rect 25452 27188 25508 28364
rect 25564 27972 25620 27982
rect 25564 27858 25620 27916
rect 25564 27806 25566 27858
rect 25618 27806 25620 27858
rect 25564 27524 25620 27806
rect 25564 27458 25620 27468
rect 25676 27412 25732 28588
rect 25676 27346 25732 27356
rect 26236 28642 26292 28654
rect 26236 28590 26238 28642
rect 26290 28590 26292 28642
rect 25564 27188 25620 27198
rect 25452 27186 25620 27188
rect 25452 27134 25566 27186
rect 25618 27134 25620 27186
rect 25452 27132 25620 27134
rect 25564 27122 25620 27132
rect 26012 26964 26068 26974
rect 24444 26852 24724 26908
rect 24332 24668 24612 24724
rect 24444 24498 24500 24510
rect 24444 24446 24446 24498
rect 24498 24446 24500 24498
rect 24444 24052 24500 24446
rect 24444 23986 24500 23996
rect 24220 23426 24276 23436
rect 24556 23938 24612 24668
rect 24556 23886 24558 23938
rect 24610 23886 24612 23938
rect 23996 23129 23998 23181
rect 24050 23129 24052 23181
rect 23996 23117 24052 23129
rect 23772 22530 23828 22540
rect 24444 22596 24500 22606
rect 24444 22502 24500 22540
rect 24556 21812 24612 23886
rect 24556 21746 24612 21756
rect 24108 21588 24164 21598
rect 24108 21494 24164 21532
rect 24332 21588 24388 21598
rect 24332 21494 24388 21532
rect 24668 21476 24724 26852
rect 25116 26852 25172 26862
rect 25116 26290 25172 26796
rect 25116 26238 25118 26290
rect 25170 26238 25172 26290
rect 25116 26226 25172 26238
rect 25452 26292 25508 26302
rect 26012 26292 26068 26908
rect 26236 26458 26292 28590
rect 26348 27858 26404 28812
rect 26460 28642 26516 30156
rect 26572 30100 26628 30940
rect 26796 30994 26852 31006
rect 26796 30942 26798 30994
rect 26850 30942 26852 30994
rect 26796 30212 26852 30942
rect 27244 30981 27246 31033
rect 27298 30981 27300 31033
rect 27132 30884 27188 30894
rect 27132 30790 27188 30828
rect 27244 30436 27300 30981
rect 26796 30146 26852 30156
rect 27132 30380 27300 30436
rect 27468 30996 27524 31006
rect 27804 30996 27860 31724
rect 28028 31556 28084 34748
rect 28252 34244 28308 34254
rect 28252 34157 28308 34188
rect 28252 34105 28254 34157
rect 28306 34105 28308 34157
rect 28252 34093 28308 34105
rect 28588 33514 28644 33526
rect 28476 33460 28532 33470
rect 28028 31490 28084 31500
rect 28140 33346 28196 33358
rect 28140 33294 28142 33346
rect 28194 33294 28196 33346
rect 26572 30034 26628 30044
rect 26684 29986 26740 29998
rect 26684 29934 26686 29986
rect 26738 29934 26740 29986
rect 26684 29650 26740 29934
rect 26684 29598 26686 29650
rect 26738 29598 26740 29650
rect 26684 29586 26740 29598
rect 27132 29652 27188 30380
rect 27244 30212 27300 30222
rect 27468 30212 27524 30940
rect 27692 30994 27860 30996
rect 27692 30942 27806 30994
rect 27858 30942 27860 30994
rect 27692 30940 27860 30942
rect 27692 30212 27748 30940
rect 27804 30930 27860 30940
rect 28140 31108 28196 33294
rect 28476 33346 28532 33404
rect 28476 33294 28478 33346
rect 28530 33294 28532 33346
rect 28476 33282 28532 33294
rect 28588 33462 28590 33514
rect 28642 33462 28644 33514
rect 28588 33348 28644 33462
rect 29484 33348 29540 33358
rect 28588 33282 28644 33292
rect 29092 33290 29148 33302
rect 29092 33238 29094 33290
rect 29146 33238 29148 33290
rect 29092 32900 29148 33238
rect 29260 33290 29316 33302
rect 29260 33238 29262 33290
rect 29314 33238 29316 33290
rect 29484 33255 29486 33292
rect 29538 33255 29540 33292
rect 29484 33243 29540 33255
rect 30044 33348 30100 33358
rect 30044 33254 30100 33292
rect 29260 33124 29316 33238
rect 29260 33058 29316 33068
rect 29092 32844 29428 32900
rect 28364 32564 28420 32574
rect 28364 32470 28420 32508
rect 28588 32564 28644 32574
rect 27916 30772 27972 30782
rect 27916 30660 27972 30716
rect 28140 30660 28196 31052
rect 27916 30604 28196 30660
rect 28476 30996 28532 31006
rect 28588 30996 28644 32508
rect 29036 32564 29092 32574
rect 28868 32452 28924 32462
rect 28868 32394 28924 32396
rect 28868 32342 28870 32394
rect 28922 32342 28924 32394
rect 28868 32330 28924 32342
rect 28700 31778 28756 31790
rect 28700 31726 28702 31778
rect 28754 31726 28756 31778
rect 28700 31556 28756 31726
rect 29036 31778 29092 32508
rect 29036 31726 29038 31778
rect 29090 31726 29092 31778
rect 29036 31714 29092 31726
rect 29204 31556 29260 31566
rect 28700 31554 29260 31556
rect 28700 31502 29206 31554
rect 29258 31502 29260 31554
rect 28700 31500 29260 31502
rect 29204 31490 29260 31500
rect 29372 31556 29428 32844
rect 30268 32116 30324 35532
rect 30380 34244 30436 38809
rect 31612 38834 31780 38836
rect 31612 38782 31726 38834
rect 31778 38782 31780 38834
rect 31612 38780 31780 38782
rect 31444 38724 31500 38734
rect 31444 38630 31500 38668
rect 31332 38276 31388 38286
rect 31612 38276 31668 38780
rect 31724 38770 31780 38780
rect 31948 38836 32004 38846
rect 31948 38742 32004 38780
rect 32060 38834 32116 38846
rect 32060 38782 32062 38834
rect 32114 38782 32116 38834
rect 32060 38724 32116 38782
rect 33124 38836 33180 38846
rect 33124 38742 33180 38780
rect 32060 38658 32116 38668
rect 31332 38274 31668 38276
rect 31332 38222 31334 38274
rect 31386 38222 31668 38274
rect 31332 38220 31668 38222
rect 31332 38210 31388 38220
rect 30828 38164 30884 38174
rect 30828 38050 30884 38108
rect 31836 38164 31892 38174
rect 31836 38070 31892 38108
rect 30828 37998 30830 38050
rect 30882 37998 30884 38050
rect 30828 37986 30884 37998
rect 31052 38050 31108 38062
rect 31052 37998 31054 38050
rect 31106 37998 31108 38050
rect 31052 37716 31108 37998
rect 31052 37650 31108 37660
rect 32172 38050 32228 38062
rect 32172 37998 32174 38050
rect 32226 37998 32228 38050
rect 32172 37492 32228 37998
rect 30716 37436 31668 37492
rect 30716 37378 30772 37436
rect 30716 37326 30718 37378
rect 30770 37326 30772 37378
rect 30716 37314 30772 37326
rect 30828 37268 30884 37278
rect 31500 37268 31556 37278
rect 30884 37266 31556 37268
rect 30884 37214 31502 37266
rect 31554 37214 31556 37266
rect 30884 37212 31556 37214
rect 30828 37202 30884 37212
rect 30716 37156 30772 37166
rect 30548 36484 30604 36494
rect 30548 36390 30604 36428
rect 30716 35922 30772 37100
rect 31500 37156 31556 37212
rect 31612 37268 31668 37436
rect 32172 37426 32228 37436
rect 33180 37604 33236 37614
rect 31836 37268 31892 37278
rect 32060 37268 32116 37278
rect 31612 37266 31892 37268
rect 31612 37214 31614 37266
rect 31666 37214 31838 37266
rect 31890 37214 31892 37266
rect 31612 37212 31892 37214
rect 31612 37202 31668 37212
rect 31836 37202 31892 37212
rect 31948 37266 32564 37268
rect 31948 37214 32062 37266
rect 32114 37214 32564 37266
rect 31948 37212 32564 37214
rect 31500 37090 31556 37100
rect 31220 37044 31276 37054
rect 30828 37042 31276 37044
rect 30828 36990 31222 37042
rect 31274 36990 31276 37042
rect 30828 36988 31276 36990
rect 30828 36482 30884 36988
rect 31220 36978 31276 36988
rect 30828 36430 30830 36482
rect 30882 36430 30884 36482
rect 30828 36418 30884 36430
rect 31052 36484 31108 36494
rect 31052 36390 31108 36428
rect 31668 36484 31724 36494
rect 31668 36390 31724 36428
rect 31948 36482 32004 37212
rect 32060 37202 32116 37212
rect 32508 37156 32564 37212
rect 33180 37266 33236 37548
rect 33180 37214 33182 37266
rect 33234 37214 33236 37266
rect 33180 37202 33236 37214
rect 32508 37100 33124 37156
rect 33068 37098 33124 37100
rect 32340 37044 32396 37054
rect 33068 37046 33070 37098
rect 33122 37046 33124 37098
rect 33068 37034 33124 37046
rect 32340 36950 32396 36988
rect 33068 36932 33124 36942
rect 31948 36430 31950 36482
rect 32002 36430 32004 36482
rect 31948 36418 32004 36430
rect 32172 36482 32228 36494
rect 32172 36430 32174 36482
rect 32226 36430 32228 36482
rect 30716 35870 30718 35922
rect 30770 35870 30772 35922
rect 30716 35700 30772 35870
rect 32172 35924 32228 36430
rect 32956 36482 33012 36494
rect 32956 36430 32958 36482
rect 33010 36430 33012 36482
rect 32956 36148 33012 36430
rect 32956 36082 33012 36092
rect 31836 35812 31892 35822
rect 30716 35634 30772 35644
rect 31052 35698 31108 35710
rect 31836 35700 31892 35756
rect 31052 35646 31054 35698
rect 31106 35646 31108 35698
rect 31052 35588 31108 35646
rect 31612 35698 31892 35700
rect 31612 35646 31838 35698
rect 31890 35646 31892 35698
rect 31612 35644 31892 35646
rect 31052 35522 31108 35532
rect 31500 35588 31556 35598
rect 31500 35494 31556 35532
rect 31612 35138 31668 35644
rect 31836 35634 31892 35644
rect 32060 35700 32116 35710
rect 32060 35606 32116 35644
rect 32172 35588 32228 35868
rect 33068 35812 33124 36876
rect 32396 35700 32452 35710
rect 32396 35606 32452 35644
rect 33068 35698 33124 35756
rect 33068 35646 33070 35698
rect 33122 35646 33124 35698
rect 33068 35634 33124 35646
rect 33180 36820 33236 36830
rect 33292 36820 33348 39452
rect 33460 39442 33516 39452
rect 33628 39060 33684 39070
rect 33404 38834 33460 38846
rect 33404 38782 33406 38834
rect 33458 38782 33460 38834
rect 33404 38276 33460 38782
rect 33628 38834 33684 39004
rect 33628 38782 33630 38834
rect 33682 38782 33684 38834
rect 33628 38770 33684 38782
rect 33404 37044 33460 38220
rect 34188 38276 34244 38286
rect 34188 38218 34244 38220
rect 34188 38166 34190 38218
rect 34242 38166 34244 38218
rect 34188 38154 34244 38166
rect 34300 38050 34356 39734
rect 34524 39620 34580 39630
rect 34524 39526 34580 39564
rect 34972 39620 35028 41692
rect 36540 41746 36652 41748
rect 36540 41694 36598 41746
rect 36650 41694 36652 41746
rect 36540 41682 36652 41694
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35420 41412 35476 41422
rect 35420 41410 35924 41412
rect 35420 41358 35422 41410
rect 35474 41358 35924 41410
rect 35420 41356 35924 41358
rect 35420 41346 35476 41356
rect 35756 41188 35812 41198
rect 35644 41186 35812 41188
rect 35644 41134 35758 41186
rect 35810 41134 35812 41186
rect 35644 41132 35812 41134
rect 34972 39058 35028 39564
rect 34972 39006 34974 39058
rect 35026 39006 35028 39058
rect 34972 38994 35028 39006
rect 35084 40402 35140 40414
rect 35084 40350 35086 40402
rect 35138 40350 35140 40402
rect 35084 38836 35140 40350
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35644 39450 35700 41132
rect 35756 41122 35812 41132
rect 35756 40516 35812 40526
rect 35756 39618 35812 40460
rect 35868 40402 35924 41356
rect 35868 40350 35870 40402
rect 35922 40350 35924 40402
rect 35868 40338 35924 40350
rect 35980 41298 36036 41310
rect 35980 41246 35982 41298
rect 36034 41246 36036 41298
rect 35756 39566 35758 39618
rect 35810 39566 35812 39618
rect 35756 39554 35812 39566
rect 35980 39579 36036 41246
rect 36428 41188 36484 41198
rect 36092 41171 36260 41188
rect 36092 41119 36094 41171
rect 36146 41132 36260 41171
rect 36146 41119 36148 41132
rect 36092 41107 36148 41119
rect 35980 39527 35982 39579
rect 36034 39527 36036 39579
rect 35980 39515 36036 39527
rect 36092 40964 36148 40974
rect 35644 39398 35646 39450
rect 35698 39398 35700 39450
rect 35644 39386 35700 39398
rect 34300 37998 34302 38050
rect 34354 37998 34356 38050
rect 33628 37828 33684 37838
rect 33516 37268 33572 37278
rect 33516 37174 33572 37212
rect 33404 36988 33572 37044
rect 33236 36764 33348 36820
rect 33180 35698 33236 36764
rect 33516 36482 33572 36988
rect 33516 36430 33518 36482
rect 33570 36430 33572 36482
rect 33516 36372 33572 36430
rect 33628 36484 33684 37772
rect 33852 37266 33908 37278
rect 33852 37214 33854 37266
rect 33906 37214 33908 37266
rect 33852 37044 33908 37214
rect 34188 37268 34244 37278
rect 34300 37268 34356 37998
rect 34636 38050 34692 38062
rect 34636 37998 34638 38050
rect 34690 37998 34692 38050
rect 34636 37940 34692 37998
rect 34636 37874 34692 37884
rect 34860 37604 34916 37614
rect 34860 37490 34916 37548
rect 34860 37438 34862 37490
rect 34914 37438 34916 37490
rect 34860 37426 34916 37438
rect 34524 37268 34580 37278
rect 34188 37266 34580 37268
rect 34188 37214 34190 37266
rect 34242 37214 34526 37266
rect 34578 37214 34580 37266
rect 34188 37212 34580 37214
rect 34188 37202 34244 37212
rect 34524 37202 34580 37212
rect 33852 36978 33908 36988
rect 34300 37098 34356 37110
rect 34300 37046 34302 37098
rect 34354 37046 34356 37098
rect 34300 37044 34356 37046
rect 34300 36978 34356 36988
rect 33740 36708 33796 36718
rect 33740 36650 33796 36652
rect 33740 36598 33742 36650
rect 33794 36598 33796 36650
rect 34860 36708 34916 36718
rect 33740 36586 33796 36598
rect 34300 36596 34356 36606
rect 34132 36484 34188 36494
rect 33628 36482 34188 36484
rect 33628 36430 34134 36482
rect 34186 36430 34188 36482
rect 33628 36428 34188 36430
rect 34132 36418 34188 36428
rect 33516 36306 33572 36316
rect 33180 35646 33182 35698
rect 33234 35646 33236 35698
rect 33180 35634 33236 35646
rect 33852 36260 33908 36270
rect 33460 35588 33516 35598
rect 32172 35522 32228 35532
rect 32508 35530 32564 35542
rect 31612 35086 31614 35138
rect 31666 35086 31668 35138
rect 31612 35074 31668 35086
rect 32396 35476 32452 35486
rect 32396 35026 32452 35420
rect 32508 35478 32510 35530
rect 32562 35478 32564 35530
rect 33460 35494 33516 35532
rect 32508 35140 32564 35478
rect 33852 35252 33908 36204
rect 34300 35810 34356 36540
rect 34524 36596 34580 36606
rect 34412 36482 34468 36494
rect 34412 36430 34414 36482
rect 34466 36430 34468 36482
rect 34412 36260 34468 36430
rect 34524 36482 34580 36540
rect 34524 36430 34526 36482
rect 34578 36430 34580 36482
rect 34860 36482 34916 36652
rect 34524 36418 34580 36430
rect 34692 36426 34748 36438
rect 34692 36374 34694 36426
rect 34746 36374 34748 36426
rect 34860 36430 34862 36482
rect 34914 36430 34916 36482
rect 34860 36418 34916 36430
rect 35084 36596 35140 38780
rect 35308 38834 35364 38846
rect 35308 38782 35310 38834
rect 35362 38782 35364 38834
rect 35308 38668 35364 38782
rect 35420 38836 35476 38846
rect 36092 38836 36148 40908
rect 36204 40628 36260 41132
rect 36428 41094 36484 41132
rect 36540 40740 36596 41682
rect 36540 40674 36596 40684
rect 36204 40562 36260 40572
rect 36876 40628 36932 41918
rect 37100 41970 37156 41982
rect 37100 41918 37102 41970
rect 37154 41918 37156 41970
rect 36876 40562 36932 40572
rect 36988 41186 37044 41198
rect 36988 41134 36990 41186
rect 37042 41134 37044 41186
rect 36988 39844 37044 41134
rect 37100 41188 37156 41918
rect 43036 41945 43038 41997
rect 43090 41945 43092 41997
rect 37436 41748 37492 41758
rect 37100 41122 37156 41132
rect 37324 41746 37492 41748
rect 37324 41694 37438 41746
rect 37490 41694 37492 41746
rect 37324 41692 37492 41694
rect 37324 41171 37380 41692
rect 37436 41682 37492 41692
rect 38332 41746 38388 41758
rect 38332 41694 38334 41746
rect 38386 41694 38388 41746
rect 37324 41119 37326 41171
rect 37378 41119 37380 41171
rect 37324 41107 37380 41119
rect 37436 41298 37492 41310
rect 37436 41246 37438 41298
rect 37490 41246 37492 41298
rect 36988 39788 37156 39844
rect 36316 39620 36372 39630
rect 36316 39526 36372 39564
rect 36988 39620 37044 39630
rect 36988 39526 37044 39564
rect 37100 39060 37156 39788
rect 37436 39579 37492 41246
rect 37660 41188 37716 41198
rect 37436 39527 37438 39579
rect 37490 39527 37492 39579
rect 37436 39515 37492 39527
rect 37548 41186 37716 41188
rect 37548 41134 37662 41186
rect 37714 41134 37716 41186
rect 37548 41132 37716 41134
rect 37548 39450 37604 41132
rect 37660 41122 37716 41132
rect 37772 41188 37828 41198
rect 37772 40514 37828 41132
rect 37996 40964 38052 40974
rect 37996 40870 38052 40908
rect 37772 40462 37774 40514
rect 37826 40462 37828 40514
rect 37772 40450 37828 40462
rect 37660 40404 37716 40414
rect 38108 40404 38164 40414
rect 38332 40404 38388 41694
rect 42028 41158 42084 41170
rect 40796 41130 40852 41142
rect 39788 41076 39844 41086
rect 37660 39618 37716 40348
rect 37660 39566 37662 39618
rect 37714 39566 37716 39618
rect 37660 39554 37716 39566
rect 37996 40402 38164 40404
rect 37996 40350 38110 40402
rect 38162 40350 38164 40402
rect 37996 40348 38164 40350
rect 37548 39398 37550 39450
rect 37602 39398 37604 39450
rect 37548 39386 37604 39398
rect 37996 39060 38052 40348
rect 38108 40338 38164 40348
rect 38220 40402 38388 40404
rect 38220 40350 38334 40402
rect 38386 40350 38388 40402
rect 38220 40348 38388 40350
rect 37100 39004 38052 39060
rect 36204 38836 36260 38846
rect 36092 38834 36260 38836
rect 36092 38782 36206 38834
rect 36258 38782 36260 38834
rect 36092 38780 36260 38782
rect 35420 38742 35476 38780
rect 36204 38770 36260 38780
rect 35308 38612 35588 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35532 37044 35588 38612
rect 36540 38052 36596 38062
rect 36540 37958 36596 37996
rect 37100 37940 37156 37950
rect 37324 37940 37380 39004
rect 38108 38948 38164 38958
rect 38220 38948 38276 40348
rect 38332 40338 38388 40348
rect 38612 40404 38668 40414
rect 38612 40310 38668 40348
rect 39788 40402 39844 41020
rect 40516 41076 40572 41086
rect 40516 40982 40572 41020
rect 40796 41078 40798 41130
rect 40850 41078 40852 41130
rect 40796 40628 40852 41078
rect 41020 41130 41076 41142
rect 41020 41078 41022 41130
rect 41074 41078 41076 41130
rect 40796 40572 40964 40628
rect 39788 40350 39790 40402
rect 39842 40350 39844 40402
rect 39788 40338 39844 40350
rect 39900 40404 39956 40414
rect 40460 40404 40516 40414
rect 39452 40178 39508 40190
rect 39452 40126 39454 40178
rect 39506 40126 39508 40178
rect 39452 39732 39508 40126
rect 39452 39666 39508 39676
rect 39564 39620 39620 39630
rect 39900 39620 39956 40348
rect 40292 40402 40516 40404
rect 40292 40350 40462 40402
rect 40514 40350 40516 40402
rect 40292 40348 40516 40350
rect 40124 40292 40180 40302
rect 40124 40198 40180 40236
rect 39452 39562 39508 39574
rect 39452 39510 39454 39562
rect 39506 39510 39508 39562
rect 39452 39060 39508 39510
rect 39452 38994 39508 39004
rect 39564 39538 39566 39564
rect 39618 39538 39620 39564
rect 38108 38946 38276 38948
rect 38108 38894 38110 38946
rect 38162 38894 38276 38946
rect 38108 38892 38276 38894
rect 38108 38882 38164 38892
rect 39564 38890 39620 39538
rect 39788 39590 39956 39620
rect 39788 39538 39790 39590
rect 39842 39564 39956 39590
rect 39842 39538 39844 39564
rect 39788 39526 39844 39538
rect 39452 38869 39508 38881
rect 39452 38836 39454 38869
rect 39506 38836 39508 38869
rect 39452 38770 39508 38780
rect 39564 38838 39566 38890
rect 39618 38838 39620 38890
rect 39340 38612 39396 38622
rect 37436 38052 37492 38062
rect 37436 37958 37492 37996
rect 38668 38052 38724 38062
rect 38668 37958 38724 37996
rect 36988 37884 37100 37940
rect 37156 37884 37380 37940
rect 35868 37828 35924 37838
rect 35868 37268 35924 37772
rect 36372 37828 36428 37838
rect 36372 37734 36428 37772
rect 35868 37174 35924 37212
rect 36092 37281 36148 37293
rect 36092 37229 36094 37281
rect 36146 37229 36148 37281
rect 36652 37281 36708 37293
rect 35532 36978 35588 36988
rect 36092 37044 36148 37229
rect 36540 37268 36596 37278
rect 36204 37156 36260 37166
rect 36204 37062 36260 37100
rect 36540 37154 36596 37212
rect 36540 37102 36542 37154
rect 36594 37102 36596 37154
rect 36540 37090 36596 37102
rect 36652 37229 36654 37281
rect 36706 37229 36708 37281
rect 36092 36978 36148 36988
rect 36652 37044 36708 37229
rect 36988 37266 37044 37884
rect 37100 37846 37156 37884
rect 36988 37214 36990 37266
rect 37042 37214 37044 37266
rect 36988 37202 37044 37214
rect 37212 37266 37268 37278
rect 37212 37214 37214 37266
rect 37266 37214 37268 37266
rect 37212 37156 37268 37214
rect 37212 37090 37268 37100
rect 37436 37268 37492 37278
rect 36652 36978 36708 36988
rect 36988 37044 37044 37054
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 34468 36204 34580 36260
rect 34412 36194 34468 36204
rect 34300 35758 34302 35810
rect 34354 35758 34356 35810
rect 34300 35746 34356 35758
rect 34412 35924 34468 35934
rect 33964 35698 34020 35710
rect 33964 35646 33966 35698
rect 34018 35646 34020 35698
rect 34412 35698 34468 35868
rect 33964 35588 34020 35646
rect 33964 35522 34020 35532
rect 34132 35642 34188 35654
rect 34132 35590 34134 35642
rect 34186 35590 34188 35642
rect 34412 35646 34414 35698
rect 34466 35646 34468 35698
rect 34412 35634 34468 35646
rect 34132 35476 34188 35590
rect 34132 35410 34188 35420
rect 33852 35196 34244 35252
rect 32508 35084 33236 35140
rect 32396 34974 32398 35026
rect 32450 34974 32452 35026
rect 32396 34962 32452 34974
rect 31948 34914 32004 34926
rect 31948 34862 31950 34914
rect 32002 34862 32004 34914
rect 30380 34178 30436 34188
rect 30492 34692 30548 34702
rect 30492 32340 30548 34636
rect 31220 34692 31276 34702
rect 31220 34598 31276 34636
rect 31948 34692 32004 34862
rect 31948 34626 32004 34636
rect 33068 34916 33124 34926
rect 32172 34244 32228 34254
rect 31948 34130 32004 34142
rect 31948 34078 31950 34130
rect 32002 34078 32004 34130
rect 31500 33460 31556 33470
rect 31276 33348 31332 33358
rect 31276 33254 31332 33292
rect 31500 33331 31556 33404
rect 31500 33279 31502 33331
rect 31554 33279 31556 33331
rect 30716 32732 31108 32788
rect 30492 32274 30548 32284
rect 30604 32564 30660 32574
rect 30604 32228 30660 32508
rect 30716 32562 30772 32732
rect 31052 32676 31108 32732
rect 30716 32510 30718 32562
rect 30770 32510 30772 32562
rect 30716 32498 30772 32510
rect 30902 32599 30958 32611
rect 30902 32547 30904 32599
rect 30956 32547 30958 32599
rect 30604 32162 30660 32172
rect 30044 32060 30324 32116
rect 30902 32116 30958 32547
rect 31052 32340 31108 32620
rect 31052 32284 31200 32340
rect 30902 32060 30996 32116
rect 29652 31946 29708 31958
rect 29652 31894 29654 31946
rect 29706 31894 29708 31946
rect 29652 31892 29708 31894
rect 29652 31826 29708 31836
rect 29484 31780 29540 31790
rect 29484 31686 29540 31724
rect 29372 31490 29428 31500
rect 28980 31220 29036 31230
rect 28980 31106 29036 31164
rect 28980 31054 28982 31106
rect 29034 31054 29036 31106
rect 28980 31042 29036 31054
rect 29596 31108 29652 31118
rect 29596 31014 29652 31052
rect 28700 30996 28756 31006
rect 28588 30994 28756 30996
rect 28588 30942 28702 30994
rect 28754 30942 28756 30994
rect 28588 30940 28756 30942
rect 27916 30212 27972 30604
rect 28084 30436 28140 30446
rect 28084 30342 28140 30380
rect 27244 30123 27246 30156
rect 27298 30123 27300 30156
rect 27244 30111 27300 30123
rect 27412 30175 27524 30212
rect 27412 30123 27414 30175
rect 27466 30156 27524 30175
rect 27636 30175 27748 30212
rect 27466 30123 27468 30156
rect 27412 30111 27468 30123
rect 27636 30123 27638 30175
rect 27690 30156 27748 30175
rect 27860 30175 27972 30212
rect 27690 30123 27692 30156
rect 27636 30111 27692 30123
rect 27860 30123 27862 30175
rect 27914 30156 27972 30175
rect 27914 30123 27916 30156
rect 27860 30111 27916 30123
rect 27244 29652 27300 29662
rect 27132 29650 27300 29652
rect 27132 29598 27246 29650
rect 27298 29598 27300 29650
rect 27132 29596 27300 29598
rect 26460 28590 26462 28642
rect 26514 28590 26516 28642
rect 26460 28578 26516 28590
rect 26796 28644 26852 28667
rect 26796 28575 26798 28588
rect 26850 28575 26852 28588
rect 27244 28642 27300 29596
rect 27244 28590 27246 28642
rect 27298 28590 27300 28642
rect 27244 28578 27300 28590
rect 27580 28644 27636 28654
rect 26796 28563 26852 28575
rect 27580 28575 27582 28588
rect 27634 28575 27636 28588
rect 26572 28474 26628 28486
rect 26348 27806 26350 27858
rect 26402 27806 26404 27858
rect 26348 27794 26404 27806
rect 26460 28420 26516 28430
rect 26348 27524 26404 27534
rect 26348 27076 26404 27468
rect 26348 26982 26404 27020
rect 26236 26406 26238 26458
rect 26290 26406 26292 26458
rect 26236 26394 26292 26406
rect 25452 26290 26068 26292
rect 25452 26238 25454 26290
rect 25506 26238 26014 26290
rect 26066 26238 26068 26290
rect 25452 26236 26068 26238
rect 25452 26226 25508 26236
rect 25564 25506 25620 26236
rect 26012 26226 26068 26236
rect 26348 26329 26404 26341
rect 26348 26277 26350 26329
rect 26402 26277 26404 26329
rect 25564 25454 25566 25506
rect 25618 25454 25620 25506
rect 26124 25506 26180 25518
rect 25564 25442 25620 25454
rect 25900 25450 25956 25462
rect 25900 25398 25902 25450
rect 25954 25398 25956 25450
rect 25564 25338 25620 25350
rect 24780 25284 24836 25294
rect 24780 24722 24836 25228
rect 25564 25286 25566 25338
rect 25618 25286 25620 25338
rect 25564 25284 25620 25286
rect 25564 25218 25620 25228
rect 25900 25172 25956 25398
rect 26124 25454 26126 25506
rect 26178 25454 26180 25506
rect 26124 25284 26180 25454
rect 26124 25218 26180 25228
rect 25900 25106 25956 25116
rect 24780 24670 24782 24722
rect 24834 24670 24836 24722
rect 24780 24658 24836 24670
rect 25452 24749 25508 24761
rect 25452 24697 25454 24749
rect 25506 24697 25508 24749
rect 25340 24052 25396 24062
rect 25340 23958 25396 23996
rect 25452 23604 25508 24697
rect 26348 24276 26404 26277
rect 26460 26292 26516 28364
rect 26572 28422 26574 28474
rect 26626 28422 26628 28474
rect 26572 27524 26628 28422
rect 27356 28474 27412 28486
rect 27356 28422 27358 28474
rect 27410 28422 27412 28474
rect 27356 28420 27412 28422
rect 27356 28354 27412 28364
rect 26572 27458 26628 27468
rect 27244 27524 27300 27534
rect 26684 27412 26740 27422
rect 26572 27074 26628 27086
rect 26572 27022 26574 27074
rect 26626 27022 26628 27074
rect 26572 26964 26628 27022
rect 26572 26516 26628 26908
rect 26684 26906 26740 27356
rect 27020 27076 27076 27086
rect 26684 26854 26686 26906
rect 26738 26854 26740 26906
rect 26684 26842 26740 26854
rect 26908 27018 26964 27030
rect 26908 26966 26910 27018
rect 26962 26966 26964 27018
rect 26572 26460 26740 26516
rect 26572 26292 26628 26302
rect 26460 26290 26628 26292
rect 26460 26238 26574 26290
rect 26626 26238 26628 26290
rect 26460 26236 26628 26238
rect 26572 26226 26628 26236
rect 26684 25506 26740 26460
rect 26908 25620 26964 26966
rect 27020 26290 27076 27020
rect 27244 27074 27300 27468
rect 27244 27022 27246 27074
rect 27298 27022 27300 27074
rect 27244 27010 27300 27022
rect 27356 27300 27412 27310
rect 27020 26238 27022 26290
rect 27074 26238 27076 26290
rect 27020 26226 27076 26238
rect 26908 25564 27188 25620
rect 26684 25454 26686 25506
rect 26738 25454 26740 25506
rect 26684 25442 26740 25454
rect 27020 25450 27076 25462
rect 27020 25398 27022 25450
rect 27074 25398 27076 25450
rect 27020 25396 27076 25398
rect 26908 25340 27076 25396
rect 26460 24500 26516 24510
rect 26460 24406 26516 24444
rect 26348 24220 26516 24276
rect 26460 23716 26516 24220
rect 25452 23538 25508 23548
rect 26124 23660 26516 23716
rect 26908 23716 26964 25340
rect 27132 25284 27188 25564
rect 27356 25506 27412 27244
rect 27356 25454 27358 25506
rect 27410 25454 27412 25506
rect 27356 25442 27412 25454
rect 27468 25508 27524 25518
rect 25116 23154 25172 23166
rect 25116 23102 25118 23154
rect 25170 23102 25172 23154
rect 25116 21476 25172 23102
rect 25900 23044 25956 23054
rect 25900 22950 25956 22988
rect 25452 22596 25508 22606
rect 25452 21613 25508 22540
rect 26124 22484 26180 23660
rect 26908 23650 26964 23660
rect 27020 25228 27188 25284
rect 27468 25338 27524 25452
rect 27468 25286 27470 25338
rect 27522 25286 27524 25338
rect 27468 25274 27524 25286
rect 26236 22484 26292 22494
rect 26124 22482 26292 22484
rect 26124 22430 26238 22482
rect 26290 22430 26292 22482
rect 26124 22428 26292 22430
rect 26236 22418 26292 22428
rect 26684 22372 26740 22382
rect 26348 22326 26404 22338
rect 26348 22274 26350 22326
rect 26402 22274 26404 22326
rect 26348 21924 26404 22274
rect 26348 21858 26404 21868
rect 25452 21561 25454 21613
rect 25506 21561 25508 21613
rect 25452 21549 25508 21561
rect 26460 21588 26516 21598
rect 25228 21476 25284 21486
rect 24668 21420 24892 21476
rect 25116 21420 25228 21476
rect 23828 21364 23884 21374
rect 23828 21362 24724 21364
rect 23828 21310 23830 21362
rect 23882 21310 24724 21362
rect 23828 21308 24724 21310
rect 23828 21298 23884 21308
rect 24668 20802 24724 21308
rect 24668 20750 24670 20802
rect 24722 20750 24724 20802
rect 24668 20738 24724 20750
rect 24836 20858 24892 21420
rect 24836 20806 24838 20858
rect 24890 20806 24892 20858
rect 24836 20580 24892 20806
rect 25116 20804 25172 20814
rect 25116 20710 25172 20748
rect 23660 19618 23716 19628
rect 23772 20524 24892 20580
rect 25004 20690 25060 20702
rect 25004 20638 25006 20690
rect 25058 20638 25060 20690
rect 23492 19294 23494 19346
rect 23546 19294 23548 19346
rect 23492 19282 23548 19294
rect 23772 19236 23828 20524
rect 24276 20020 24332 20030
rect 24276 19926 24332 19964
rect 24724 19906 24780 19918
rect 24724 19854 24726 19906
rect 24778 19854 24780 19906
rect 22540 18498 22596 18508
rect 23660 19234 23828 19236
rect 23660 19182 23774 19234
rect 23826 19182 23828 19234
rect 23660 19180 23828 19182
rect 22204 18398 22206 18450
rect 22258 18398 22260 18450
rect 22876 18452 22932 18462
rect 23660 18452 23716 19180
rect 23772 19170 23828 19180
rect 23996 19796 24052 19806
rect 22204 18004 22260 18398
rect 22092 17948 22204 18004
rect 21868 17780 21924 17790
rect 21644 17778 21924 17780
rect 21644 17726 21870 17778
rect 21922 17726 21924 17778
rect 21644 17724 21924 17726
rect 20860 17668 20916 17678
rect 20860 17574 20916 17612
rect 21532 17666 21588 17724
rect 21868 17714 21924 17724
rect 21532 17614 21534 17666
rect 21586 17614 21588 17666
rect 21532 17108 21588 17614
rect 21924 17610 21980 17622
rect 21924 17558 21926 17610
rect 21978 17558 21980 17610
rect 21924 17556 21980 17558
rect 22092 17556 22148 17948
rect 22204 17938 22260 17948
rect 22372 18394 22428 18406
rect 22372 18342 22374 18394
rect 22426 18342 22428 18394
rect 22876 18358 22932 18396
rect 23548 18396 23716 18452
rect 23996 18452 24052 19740
rect 24724 19796 24780 19854
rect 24724 19730 24780 19740
rect 24220 19684 24276 19694
rect 22372 17780 22428 18342
rect 23118 18226 23174 18238
rect 23118 18174 23120 18226
rect 23172 18174 23174 18226
rect 22372 17724 22484 17780
rect 21924 17500 22148 17556
rect 22204 17666 22260 17678
rect 22204 17614 22206 17666
rect 22258 17614 22260 17666
rect 22204 17556 22260 17614
rect 22204 17490 22260 17500
rect 21532 17042 21588 17052
rect 22428 17444 22484 17724
rect 23118 17668 23174 18174
rect 23118 17602 23174 17612
rect 22428 16994 22484 17388
rect 23548 17108 23604 18396
rect 23996 18358 24052 18396
rect 24108 19348 24164 19358
rect 23754 18340 23810 18350
rect 23754 18246 23810 18284
rect 24108 17892 24164 19292
rect 23660 17834 23716 17846
rect 23660 17782 23662 17834
rect 23714 17782 23716 17834
rect 23660 17780 23716 17782
rect 23660 17714 23716 17724
rect 23996 17836 24164 17892
rect 23772 17668 23828 17678
rect 23772 17666 23940 17668
rect 23772 17614 23774 17666
rect 23826 17614 23940 17666
rect 23772 17612 23940 17614
rect 23772 17602 23828 17612
rect 22428 16942 22430 16994
rect 22482 16942 22484 16994
rect 22428 16930 22484 16942
rect 23324 17052 23604 17108
rect 23100 16658 23156 16670
rect 23100 16606 23102 16658
rect 23154 16606 23156 16658
rect 23100 16212 23156 16606
rect 23100 16146 23156 16156
rect 22876 16100 22932 16110
rect 22876 16006 22932 16044
rect 23324 16100 23380 17052
rect 23436 16884 23492 16894
rect 23754 16884 23810 16894
rect 23436 16882 23810 16884
rect 23436 16830 23438 16882
rect 23490 16830 23756 16882
rect 23808 16830 23810 16882
rect 23436 16828 23810 16830
rect 23436 16818 23492 16828
rect 23754 16818 23810 16828
rect 23884 16324 23940 17612
rect 23996 16884 24052 17836
rect 24108 17668 24164 17678
rect 24108 17574 24164 17612
rect 23996 16790 24052 16828
rect 24220 16772 24276 19628
rect 25004 19572 25060 20638
rect 25228 20244 25284 21420
rect 26460 21474 26516 21532
rect 26460 21422 26462 21474
rect 26514 21422 26516 21474
rect 25396 21028 25452 21038
rect 25396 20934 25452 20972
rect 26460 20804 26516 21422
rect 26684 20916 26740 22316
rect 26684 20850 26740 20860
rect 26796 21924 26852 21934
rect 26572 20804 26628 20814
rect 26460 20802 26628 20804
rect 26460 20750 26574 20802
rect 26626 20750 26628 20802
rect 26460 20748 26628 20750
rect 26572 20738 26628 20748
rect 26796 20692 26852 21868
rect 26908 20916 26964 20926
rect 27020 20916 27076 25228
rect 27468 25172 27524 25182
rect 27244 23828 27300 23838
rect 27244 23734 27300 23772
rect 27468 22820 27524 25116
rect 27468 22754 27524 22764
rect 27468 22370 27524 22382
rect 27468 22318 27470 22370
rect 27522 22318 27524 22370
rect 27132 22148 27188 22158
rect 27132 22146 27300 22148
rect 27132 22094 27134 22146
rect 27186 22094 27300 22146
rect 27132 22092 27300 22094
rect 27132 22082 27188 22092
rect 26908 20914 27076 20916
rect 26908 20862 26910 20914
rect 26962 20862 27076 20914
rect 26908 20860 27076 20862
rect 26908 20850 26964 20860
rect 27244 20802 27300 22092
rect 27020 20758 27076 20770
rect 27020 20706 27022 20758
rect 27074 20706 27076 20758
rect 27020 20692 27076 20706
rect 26796 20636 27076 20692
rect 27244 20750 27246 20802
rect 27298 20750 27300 20802
rect 26908 20580 26964 20636
rect 26852 20524 26964 20580
rect 26348 20468 26404 20478
rect 25340 20244 25396 20254
rect 25228 20242 25396 20244
rect 25228 20190 25342 20242
rect 25394 20190 25396 20242
rect 25228 20188 25396 20190
rect 25340 20178 25396 20188
rect 24332 19516 25060 19572
rect 25676 20018 25732 20030
rect 25676 19966 25678 20018
rect 25730 19966 25732 20018
rect 24332 17892 24388 19516
rect 24556 19236 24612 19246
rect 24556 19234 24836 19236
rect 24556 19182 24558 19234
rect 24610 19182 24836 19234
rect 24556 19180 24836 19182
rect 24556 19170 24612 19180
rect 24668 18450 24724 18462
rect 24500 18394 24556 18406
rect 24500 18342 24502 18394
rect 24554 18342 24556 18394
rect 24500 18228 24556 18342
rect 24500 18162 24556 18172
rect 24668 18398 24670 18450
rect 24722 18398 24724 18450
rect 24332 17826 24388 17836
rect 24444 18004 24500 18014
rect 24444 17834 24500 17948
rect 24444 17782 24446 17834
rect 24498 17782 24500 17834
rect 24444 17770 24500 17782
rect 24556 17780 24612 17790
rect 24556 17666 24612 17724
rect 24556 17614 24558 17666
rect 24610 17614 24612 17666
rect 24556 17602 24612 17614
rect 24500 17108 24556 17118
rect 24500 16938 24556 17052
rect 24500 16886 24502 16938
rect 24554 16886 24556 16938
rect 24500 16874 24556 16886
rect 24668 16882 24724 18398
rect 24780 18452 24836 19180
rect 24780 18386 24836 18396
rect 25116 18450 25172 18462
rect 25116 18398 25118 18450
rect 25170 18398 25172 18450
rect 25116 18340 25172 18398
rect 25452 18452 25508 18462
rect 25452 18358 25508 18396
rect 25116 18274 25172 18284
rect 25452 17892 25508 17902
rect 25340 17780 25396 17790
rect 25228 17778 25396 17780
rect 25228 17726 25342 17778
rect 25394 17726 25396 17778
rect 25228 17724 25396 17726
rect 24220 16706 24276 16716
rect 24668 16830 24670 16882
rect 24722 16830 24724 16882
rect 24668 16548 24724 16830
rect 24668 16482 24724 16492
rect 24892 17666 24948 17678
rect 24892 17614 24894 17666
rect 24946 17614 24948 17666
rect 23884 16258 23940 16268
rect 24892 16324 24948 17614
rect 24892 16258 24948 16268
rect 23660 16212 23716 16222
rect 23660 16118 23716 16156
rect 23324 16034 23380 16044
rect 23772 15540 23828 15550
rect 23772 15426 23828 15484
rect 24276 15540 24332 15550
rect 24276 15446 24332 15484
rect 23772 15374 23774 15426
rect 23826 15374 23828 15426
rect 23772 15362 23828 15374
rect 21756 15316 21812 15326
rect 21756 15222 21812 15260
rect 22540 15316 22596 15326
rect 22858 15316 22914 15326
rect 22540 15314 22914 15316
rect 22540 15262 22542 15314
rect 22594 15262 22860 15314
rect 22912 15262 22914 15314
rect 22540 15260 22914 15262
rect 22540 15250 22596 15260
rect 22858 15250 22914 15260
rect 23100 15314 23156 15326
rect 23100 15262 23102 15314
rect 23154 15262 23156 15314
rect 21420 15202 21476 15214
rect 21420 15150 21422 15202
rect 21474 15150 21476 15202
rect 21196 14644 21252 14654
rect 21196 12962 21252 14588
rect 21420 14644 21476 15150
rect 23100 15204 23156 15262
rect 22204 15092 22260 15102
rect 21420 14578 21476 14588
rect 21980 15090 22260 15092
rect 21980 15038 22206 15090
rect 22258 15038 22260 15090
rect 21980 15036 22260 15038
rect 21420 14502 21476 14514
rect 21420 14450 21422 14502
rect 21474 14450 21476 14502
rect 21308 13972 21364 13982
rect 21308 13858 21364 13916
rect 21308 13806 21310 13858
rect 21362 13806 21364 13858
rect 21308 13794 21364 13806
rect 21196 12910 21198 12962
rect 21250 12910 21252 12962
rect 21196 12898 21252 12910
rect 18620 12124 18788 12141
rect 18620 11620 18676 12124
rect 18844 12068 18900 12078
rect 18620 11554 18676 11564
rect 18732 12066 18900 12068
rect 18732 12014 18846 12066
rect 18898 12014 18900 12066
rect 18732 12012 18900 12014
rect 18396 11442 18452 11452
rect 18732 11506 18788 12012
rect 18844 12002 18900 12012
rect 18732 11454 18734 11506
rect 18786 11454 18788 11506
rect 18732 11442 18788 11454
rect 19852 11620 19908 11630
rect 19852 11172 19908 11564
rect 20076 11284 20132 12348
rect 20748 12338 20804 12348
rect 21420 12178 21476 14450
rect 21420 12126 21422 12178
rect 21474 12126 21476 12178
rect 21420 11844 21476 12126
rect 21868 13748 21924 13758
rect 21868 12178 21924 13692
rect 21980 13074 22036 15036
rect 22204 15026 22260 15036
rect 22988 15092 23156 15148
rect 23604 15258 23660 15270
rect 23604 15206 23606 15258
rect 23658 15206 23660 15258
rect 23604 15148 23660 15206
rect 24444 15204 24500 15214
rect 23604 15092 23828 15148
rect 22988 14980 23044 15092
rect 22988 14914 23044 14924
rect 22652 14308 22708 14318
rect 22652 14214 22708 14252
rect 21980 13022 21982 13074
rect 22034 13022 22036 13074
rect 21980 13010 22036 13022
rect 23100 13972 23156 13982
rect 23100 12404 23156 13916
rect 23212 13636 23268 13646
rect 23212 13542 23268 13580
rect 21868 12126 21870 12178
rect 21922 12126 21924 12178
rect 21868 12114 21924 12126
rect 22876 12348 23156 12404
rect 23772 12852 23828 15092
rect 24444 14530 24500 15148
rect 24444 14478 24446 14530
rect 24498 14478 24500 14530
rect 25116 14532 25172 14542
rect 25228 14532 25284 17724
rect 25340 17714 25396 17724
rect 25452 17666 25508 17836
rect 25452 17614 25454 17666
rect 25506 17614 25508 17666
rect 25452 17602 25508 17614
rect 25452 17108 25508 17118
rect 25340 16884 25396 16894
rect 25340 15550 25396 16828
rect 25452 16212 25508 17052
rect 25564 16212 25620 16222
rect 25452 16210 25620 16212
rect 25452 16158 25566 16210
rect 25618 16158 25620 16210
rect 25452 16156 25620 16158
rect 25564 16146 25620 16156
rect 25340 15538 25452 15550
rect 25340 15486 25398 15538
rect 25450 15486 25452 15538
rect 25340 15484 25452 15486
rect 25396 15474 25452 15484
rect 25676 15148 25732 19966
rect 26348 20020 26404 20412
rect 26852 20130 26908 20524
rect 27244 20356 27300 20750
rect 26852 20078 26854 20130
rect 26906 20078 26908 20130
rect 26852 20066 26908 20078
rect 27020 20300 27300 20356
rect 27356 20804 27412 20814
rect 26348 19926 26404 19964
rect 27020 20020 27076 20300
rect 27020 19954 27076 19964
rect 27132 20132 27188 20142
rect 27132 20018 27188 20076
rect 27356 20020 27412 20748
rect 27468 20468 27524 22318
rect 27580 22316 27636 28575
rect 28028 28308 28084 28318
rect 27804 27242 27860 27254
rect 27804 27190 27806 27242
rect 27858 27190 27860 27242
rect 27804 27188 27860 27190
rect 27804 27122 27860 27132
rect 28028 27074 28084 28252
rect 28252 27972 28308 27982
rect 28476 27972 28532 30940
rect 28700 30930 28756 30940
rect 29260 30996 29316 31006
rect 29260 30902 29316 30940
rect 30044 30660 30100 32060
rect 30268 31778 30324 31790
rect 30268 31726 30270 31778
rect 30322 31726 30324 31778
rect 30268 31668 30324 31726
rect 30268 31602 30324 31612
rect 30940 31444 30996 32060
rect 30324 31388 30996 31444
rect 31144 31722 31200 32284
rect 31144 31670 31146 31722
rect 31198 31670 31200 31722
rect 31276 32338 31332 32350
rect 31276 32286 31278 32338
rect 31330 32286 31332 32338
rect 31276 31780 31332 32286
rect 31276 31714 31332 31724
rect 31388 31780 31444 31790
rect 31500 31780 31556 33279
rect 31388 31778 31556 31780
rect 31388 31726 31390 31778
rect 31442 31726 31556 31778
rect 31388 31724 31556 31726
rect 31612 33458 31668 33470
rect 31612 33406 31614 33458
rect 31666 33406 31668 33458
rect 31612 32340 31668 33406
rect 31948 33348 32004 34078
rect 31948 33282 32004 33292
rect 32172 33346 32228 34188
rect 33068 34242 33124 34860
rect 33180 34692 33236 35084
rect 33180 34636 33262 34692
rect 33068 34190 33070 34242
rect 33122 34190 33124 34242
rect 33068 34178 33124 34190
rect 33206 34170 33262 34636
rect 34188 34186 34244 35196
rect 34300 34916 34356 34926
rect 34300 34822 34356 34860
rect 32284 34130 32340 34142
rect 32284 34078 32286 34130
rect 32338 34078 32340 34130
rect 33206 34118 33208 34170
rect 33260 34118 33262 34170
rect 33206 34106 33262 34118
rect 33516 34163 33572 34175
rect 33516 34132 33518 34163
rect 33570 34132 33572 34163
rect 32284 33460 32340 34078
rect 33516 34066 33572 34076
rect 33852 34166 33908 34178
rect 33852 34114 33854 34166
rect 33906 34114 33908 34166
rect 34188 34134 34190 34186
rect 34242 34134 34244 34186
rect 34188 34122 34244 34134
rect 32396 33962 32452 33974
rect 32396 33910 32398 33962
rect 32450 33910 32452 33962
rect 32396 33572 32452 33910
rect 32396 33506 32452 33516
rect 32284 33394 32340 33404
rect 32172 33294 32174 33346
rect 32226 33294 32228 33346
rect 32172 33282 32228 33294
rect 31836 32676 31892 32686
rect 31724 32564 31780 32574
rect 31724 32470 31780 32508
rect 31836 32562 31892 32620
rect 31836 32510 31838 32562
rect 31890 32510 31892 32562
rect 31836 32498 31892 32510
rect 31982 32599 32038 32611
rect 31982 32547 31984 32599
rect 32036 32547 32038 32599
rect 31982 32340 32038 32547
rect 33404 32562 33460 32574
rect 33404 32510 33406 32562
rect 33458 32510 33460 32562
rect 31612 32284 31982 32340
rect 31388 31714 31444 31724
rect 30324 31218 30380 31388
rect 30324 31166 30326 31218
rect 30378 31166 30380 31218
rect 30324 31154 30380 31166
rect 31144 31220 31200 31670
rect 31144 31154 31200 31164
rect 30492 31108 30548 31118
rect 30156 30994 30212 31006
rect 30156 30942 30158 30994
rect 30210 30942 30212 30994
rect 30156 30884 30212 30942
rect 30156 30818 30212 30828
rect 30044 30604 30324 30660
rect 28252 27970 28532 27972
rect 28252 27918 28254 27970
rect 28306 27918 28532 27970
rect 28252 27916 28532 27918
rect 28812 28644 28868 28654
rect 28252 27906 28308 27916
rect 28812 27902 28868 28588
rect 29820 28532 29876 28542
rect 28812 27850 28814 27902
rect 28866 27850 28868 27902
rect 28812 27838 28868 27850
rect 29148 28420 29204 28430
rect 29148 27858 29204 28364
rect 29148 27806 29150 27858
rect 29202 27806 29204 27858
rect 28700 27746 28756 27758
rect 28700 27694 28702 27746
rect 28754 27694 28756 27746
rect 28700 27300 28756 27694
rect 28700 27234 28756 27244
rect 28028 27022 28030 27074
rect 28082 27022 28084 27074
rect 28028 27010 28084 27022
rect 28588 27074 28644 27086
rect 28588 27022 28590 27074
rect 28642 27022 28644 27074
rect 28588 26516 28644 27022
rect 29148 26964 29204 27806
rect 29820 27858 29876 28476
rect 30268 28308 30324 30604
rect 30268 28242 30324 28252
rect 29820 27806 29822 27858
rect 29874 27806 29876 27858
rect 29820 27794 29876 27806
rect 29652 27634 29708 27646
rect 29652 27582 29654 27634
rect 29706 27582 29708 27634
rect 29652 27188 29708 27582
rect 29652 27122 29708 27132
rect 30268 27188 30324 27198
rect 30268 27094 30324 27132
rect 29484 27074 29540 27086
rect 29484 27022 29486 27074
rect 29538 27022 29540 27074
rect 29484 26908 29540 27022
rect 29148 26898 29204 26908
rect 28588 26450 28644 26460
rect 29372 26852 29540 26908
rect 29708 26964 29764 26974
rect 27804 26180 27860 26190
rect 27804 26178 28084 26180
rect 27804 26126 27806 26178
rect 27858 26126 28084 26178
rect 27804 26124 28084 26126
rect 27804 26114 27860 26124
rect 28028 25732 28084 26124
rect 29372 26068 29428 26852
rect 28140 25732 28196 25742
rect 28028 25730 28196 25732
rect 28028 25678 28142 25730
rect 28194 25678 28196 25730
rect 28028 25676 28196 25678
rect 28140 25666 28196 25676
rect 27804 25508 27860 25518
rect 27804 25414 27860 25452
rect 28476 25284 28532 25294
rect 28140 24722 28196 24734
rect 28364 24724 28420 24734
rect 28140 24670 28142 24722
rect 28194 24670 28196 24722
rect 27692 23828 27748 23838
rect 28140 23828 28196 24670
rect 27748 23772 28196 23828
rect 28252 24722 28420 24724
rect 28252 24670 28366 24722
rect 28418 24670 28420 24722
rect 28252 24668 28420 24670
rect 27692 23044 27748 23772
rect 28252 23604 28308 24668
rect 28364 24658 28420 24668
rect 28140 23548 28308 23604
rect 27804 23268 27860 23278
rect 28140 23268 28196 23548
rect 27804 23266 28196 23268
rect 27804 23214 27806 23266
rect 27858 23214 28196 23266
rect 27804 23212 28196 23214
rect 27804 23202 27860 23212
rect 28140 23154 28196 23212
rect 28140 23102 28142 23154
rect 28194 23102 28196 23154
rect 28140 23090 28196 23102
rect 28308 23044 28364 23054
rect 27692 22988 27972 23044
rect 27692 22820 27748 22830
rect 27692 22482 27748 22764
rect 27692 22430 27694 22482
rect 27746 22430 27748 22482
rect 27692 22418 27748 22430
rect 27916 22372 27972 22988
rect 28308 22986 28364 22988
rect 28308 22934 28310 22986
rect 28362 22934 28364 22986
rect 28308 22922 28364 22934
rect 28028 22372 28084 22382
rect 27916 22370 28084 22372
rect 27748 22340 27804 22352
rect 27748 22316 27750 22340
rect 27580 22288 27750 22316
rect 27802 22316 27804 22340
rect 27916 22318 28030 22370
rect 28082 22318 28084 22370
rect 27916 22316 28084 22318
rect 27802 22288 27860 22316
rect 28028 22306 28084 22316
rect 27580 22260 27860 22288
rect 27804 21700 27860 22260
rect 28364 21924 28420 21934
rect 27804 21644 28196 21700
rect 28140 20914 28196 21644
rect 28364 21630 28420 21868
rect 28476 21754 28532 25228
rect 28644 24836 28700 24846
rect 28644 24742 28700 24780
rect 29260 24722 29316 24734
rect 29260 24670 29262 24722
rect 29314 24670 29316 24722
rect 29148 24500 29204 24510
rect 28700 24052 28756 24062
rect 28700 23938 28756 23996
rect 28700 23886 28702 23938
rect 28754 23886 28756 23938
rect 28700 23210 28756 23886
rect 29148 23910 29204 24444
rect 29260 24052 29316 24670
rect 29372 24722 29428 26012
rect 29372 24670 29374 24722
rect 29426 24670 29428 24722
rect 29372 24658 29428 24670
rect 29484 26516 29540 26526
rect 29260 23986 29316 23996
rect 29148 23858 29150 23910
rect 29202 23858 29204 23910
rect 29148 23846 29204 23858
rect 29484 23828 29540 26460
rect 29708 26402 29764 26908
rect 29708 26350 29710 26402
rect 29762 26350 29764 26402
rect 29708 26338 29764 26350
rect 29932 25508 29988 25518
rect 29764 25506 29988 25508
rect 29764 25454 29934 25506
rect 29986 25454 29988 25506
rect 29764 25452 29988 25454
rect 29764 25396 29820 25452
rect 29932 25442 29988 25452
rect 29764 25302 29820 25340
rect 29652 24500 29708 24510
rect 29652 24498 29764 24500
rect 29652 24446 29654 24498
rect 29706 24446 29764 24498
rect 29652 24434 29764 24446
rect 29260 23772 29540 23828
rect 29148 23716 29204 23726
rect 28700 23158 28702 23210
rect 28754 23158 28756 23210
rect 28700 23146 28756 23158
rect 28812 23380 28868 23390
rect 28812 23182 28868 23324
rect 28812 23130 28814 23182
rect 28866 23130 28868 23182
rect 28812 22932 28868 23130
rect 28812 22866 28868 22876
rect 29036 23182 29092 23194
rect 29036 23130 29038 23182
rect 29090 23130 29092 23182
rect 28476 21702 28478 21754
rect 28530 21702 28532 21754
rect 28476 21690 28532 21702
rect 28588 22372 28644 22382
rect 28588 22158 28644 22316
rect 28588 22146 28700 22158
rect 28588 22094 28646 22146
rect 28698 22094 28700 22146
rect 28588 22082 28700 22094
rect 28364 21578 28366 21630
rect 28418 21578 28420 21630
rect 28364 21566 28420 21578
rect 28140 20862 28142 20914
rect 28194 20862 28196 20914
rect 28140 20850 28196 20862
rect 27692 20804 27748 20814
rect 28588 20804 28644 22082
rect 28700 21700 28756 21710
rect 28700 21588 28756 21644
rect 28700 21586 28868 21588
rect 28700 21534 28702 21586
rect 28754 21534 28868 21586
rect 28700 21532 28868 21534
rect 28700 21522 28756 21532
rect 27692 20710 27748 20748
rect 28028 20758 28084 20770
rect 27468 20402 27524 20412
rect 28028 20706 28030 20758
rect 28082 20706 28084 20758
rect 28028 20132 28084 20706
rect 28476 20748 28644 20804
rect 28476 20244 28532 20748
rect 28644 20578 28700 20590
rect 28644 20526 28646 20578
rect 28698 20526 28700 20578
rect 28644 20468 28700 20526
rect 28644 20402 28700 20412
rect 28028 20066 28084 20076
rect 28364 20186 28420 20198
rect 28476 20188 28644 20244
rect 28364 20134 28366 20186
rect 28418 20134 28420 20186
rect 27132 19966 27134 20018
rect 27186 19966 27188 20018
rect 27132 19954 27188 19966
rect 27244 20018 27412 20020
rect 27244 19966 27358 20018
rect 27410 19966 27412 20018
rect 27244 19964 27412 19966
rect 26012 19796 26068 19806
rect 27244 19796 27300 19964
rect 27356 19954 27412 19964
rect 27468 20018 27524 20030
rect 27468 19966 27470 20018
rect 27522 19966 27524 20018
rect 26012 19794 26292 19796
rect 26012 19742 26014 19794
rect 26066 19742 26292 19794
rect 26012 19740 26292 19742
rect 26012 19730 26068 19740
rect 25788 18340 25844 18350
rect 25788 17780 25844 18284
rect 25788 16882 25844 17724
rect 25788 16830 25790 16882
rect 25842 16830 25844 16882
rect 25788 16818 25844 16830
rect 26012 17892 26068 17902
rect 26012 16884 26068 17836
rect 26012 16790 26068 16828
rect 26124 17668 26180 17678
rect 25900 16770 25956 16782
rect 25900 16718 25902 16770
rect 25954 16718 25956 16770
rect 25900 15540 25956 16718
rect 25116 14530 25284 14532
rect 24444 14466 24500 14478
rect 24948 14474 25004 14486
rect 24202 14420 24258 14430
rect 24948 14422 24950 14474
rect 25002 14422 25004 14474
rect 25116 14478 25118 14530
rect 25170 14478 25284 14530
rect 25116 14476 25284 14478
rect 25116 14466 25172 14476
rect 24202 14418 24276 14420
rect 24202 14366 24204 14418
rect 24256 14366 24276 14418
rect 24202 14354 24276 14366
rect 23996 13748 24052 13758
rect 23996 13654 24052 13692
rect 24108 13748 24164 13758
rect 24220 13748 24276 14354
rect 24948 13972 25004 14422
rect 24948 13906 25004 13916
rect 24108 13746 24276 13748
rect 24108 13694 24110 13746
rect 24162 13694 24276 13746
rect 24108 13692 24276 13694
rect 24108 13682 24164 13692
rect 24444 13636 24500 13646
rect 24444 13542 24500 13580
rect 23884 12852 23940 12862
rect 23772 12850 23940 12852
rect 23772 12798 23886 12850
rect 23938 12798 23940 12850
rect 23772 12796 23940 12798
rect 22652 12066 22708 12078
rect 22652 12014 22654 12066
rect 22706 12014 22708 12066
rect 21420 11788 21924 11844
rect 20636 11508 20692 11518
rect 20636 11414 20692 11452
rect 21644 11366 21700 11378
rect 21644 11314 21646 11366
rect 21698 11314 21700 11366
rect 20076 11228 20244 11284
rect 18060 11106 18116 11116
rect 19628 11116 19908 11172
rect 17500 10625 17556 10637
rect 17500 10573 17502 10625
rect 17554 10573 17556 10625
rect 17388 10500 17444 10510
rect 17388 10406 17444 10444
rect 16940 9940 16996 9950
rect 17500 9940 17556 10573
rect 16940 9938 17556 9940
rect 16940 9886 16942 9938
rect 16994 9886 17556 9938
rect 16940 9884 17556 9886
rect 17836 10612 17892 10622
rect 16940 9874 16996 9884
rect 16772 9266 16884 9278
rect 16772 9214 16774 9266
rect 16826 9214 16884 9266
rect 16772 9212 16884 9214
rect 16940 9604 16996 9614
rect 16772 9202 16828 9212
rect 16324 9044 16380 9054
rect 16324 8874 16380 8988
rect 16324 8822 16326 8874
rect 16378 8822 16380 8874
rect 16492 9042 16548 9054
rect 16492 8990 16494 9042
rect 16546 8990 16548 9042
rect 16492 8932 16548 8990
rect 16940 9042 16996 9548
rect 16940 8990 16942 9042
rect 16994 8990 16996 9042
rect 16940 8978 16996 8990
rect 16492 8866 16548 8876
rect 16324 8810 16380 8822
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 16492 8260 16548 8270
rect 16492 8258 16828 8260
rect 16492 8206 16494 8258
rect 16546 8206 16828 8258
rect 16492 8204 16828 8206
rect 16492 8194 16548 8204
rect 16772 7698 16828 8204
rect 17052 8148 17108 9884
rect 17836 9604 17892 10556
rect 18956 10610 19012 10622
rect 18956 10558 18958 10610
rect 19010 10558 19012 10610
rect 18620 10386 18676 10398
rect 18620 10334 18622 10386
rect 18674 10334 18676 10386
rect 17948 10052 18004 10062
rect 17948 9798 18004 9996
rect 17948 9746 17950 9798
rect 18002 9746 18004 9798
rect 18620 9828 18676 10334
rect 18620 9762 18676 9772
rect 18732 10052 18788 10062
rect 17948 9734 18004 9746
rect 17836 9538 17892 9548
rect 17948 9156 18004 9166
rect 17948 9042 18004 9100
rect 17948 8990 17950 9042
rect 18002 8990 18004 9042
rect 17948 8978 18004 8990
rect 18340 9071 18396 9083
rect 18340 9019 18342 9071
rect 18394 9044 18396 9071
rect 18394 9019 18452 9044
rect 18340 8988 18452 9019
rect 18172 8932 18228 8942
rect 18060 8930 18228 8932
rect 18060 8878 18174 8930
rect 18226 8878 18228 8930
rect 18060 8876 18228 8878
rect 17780 8820 17836 8830
rect 17780 8726 17836 8764
rect 18060 8596 18116 8876
rect 18172 8866 18228 8876
rect 17276 8540 18116 8596
rect 17276 8370 17332 8540
rect 17276 8318 17278 8370
rect 17330 8318 17332 8370
rect 17276 8306 17332 8318
rect 18396 8372 18452 8988
rect 18620 9042 18676 9054
rect 18620 8990 18622 9042
rect 18674 8990 18676 9042
rect 18620 8932 18676 8990
rect 18620 8708 18676 8876
rect 18620 8642 18676 8652
rect 18396 8316 18564 8372
rect 17052 8092 17556 8148
rect 16772 7646 16774 7698
rect 16826 7646 16828 7698
rect 16772 7634 16828 7646
rect 17500 7518 17556 8092
rect 16940 7476 16996 7486
rect 17500 7466 17502 7518
rect 17554 7466 17556 7518
rect 18508 7489 18564 8316
rect 18732 8260 18788 9996
rect 18956 9268 19012 10558
rect 18956 9202 19012 9212
rect 19292 10498 19348 10510
rect 19292 10446 19294 10498
rect 19346 10446 19348 10498
rect 19292 9716 19348 10446
rect 19292 9156 19348 9660
rect 19628 9156 19684 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10836 20244 11228
rect 20076 10780 20244 10836
rect 20076 10276 20132 10780
rect 21196 10498 21252 10510
rect 21196 10446 21198 10498
rect 21250 10446 21252 10498
rect 20076 10220 20468 10276
rect 19740 9940 19796 9950
rect 19740 9846 19796 9884
rect 20412 9798 20468 10220
rect 20412 9746 20414 9798
rect 20466 9746 20468 9798
rect 20412 9734 20468 9746
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 9100 19908 9156
rect 19292 9090 19348 9100
rect 18844 9044 18900 9054
rect 18844 8950 18900 8988
rect 19628 8932 19684 8942
rect 17500 7454 17556 7466
rect 17724 7476 17780 7486
rect 16940 7382 16996 7420
rect 17388 7362 17444 7374
rect 17388 7310 17390 7362
rect 17442 7310 17444 7362
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 17388 7028 17444 7310
rect 4476 7018 4740 7028
rect 16828 6972 17444 7028
rect 15820 6692 15876 6702
rect 15820 6690 16380 6692
rect 15820 6638 15822 6690
rect 15874 6638 16380 6690
rect 15820 6636 16380 6638
rect 15820 6626 15876 6636
rect 16324 6130 16380 6636
rect 16324 6078 16326 6130
rect 16378 6078 16380 6130
rect 16324 6066 16380 6078
rect 16604 6690 16660 6702
rect 16604 6638 16606 6690
rect 16658 6638 16660 6690
rect 15148 5908 15204 5918
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 15148 5234 15204 5852
rect 16492 5908 16548 5918
rect 16492 5814 16548 5852
rect 16604 5796 16660 6638
rect 16828 6244 16884 6972
rect 16828 6188 17108 6244
rect 16940 6020 16996 6030
rect 16940 5906 16996 5964
rect 16940 5854 16942 5906
rect 16994 5854 16996 5906
rect 16940 5842 16996 5854
rect 16604 5730 16660 5740
rect 16772 5684 16828 5694
rect 16772 5590 16828 5628
rect 15148 5182 15150 5234
rect 15202 5182 15204 5234
rect 15148 5170 15204 5182
rect 17052 5234 17108 6188
rect 17724 6132 17780 7420
rect 17612 6020 17668 6030
rect 17500 5921 17556 5933
rect 17500 5869 17502 5921
rect 17554 5869 17556 5921
rect 17388 5796 17444 5806
rect 17388 5702 17444 5740
rect 17052 5182 17054 5234
rect 17106 5182 17108 5234
rect 17052 5170 17108 5182
rect 17500 5012 17556 5869
rect 17500 4946 17556 4956
rect 17612 4338 17668 5964
rect 17724 5906 17780 6076
rect 17724 5854 17726 5906
rect 17778 5854 17780 5906
rect 17724 5842 17780 5854
rect 17836 7474 17892 7486
rect 17836 7422 17838 7474
rect 17890 7422 17892 7474
rect 17836 5908 17892 7422
rect 18508 7437 18510 7489
rect 18562 7437 18564 7489
rect 18508 6916 18564 7437
rect 18620 8204 18788 8260
rect 18956 8930 19684 8932
rect 18956 8878 19630 8930
rect 19682 8878 19684 8930
rect 18956 8876 19684 8878
rect 18620 7028 18676 8204
rect 18956 8148 19012 8876
rect 19628 8866 19684 8876
rect 19740 8932 19796 8942
rect 19180 8708 19236 8718
rect 18732 8092 19012 8148
rect 19068 8372 19124 8382
rect 18732 7642 18788 8092
rect 18732 7590 18734 7642
rect 18786 7590 18788 7642
rect 18732 7578 18788 7590
rect 18844 7924 18900 7934
rect 18844 7474 18900 7868
rect 18844 7422 18846 7474
rect 18898 7422 18900 7474
rect 18844 7410 18900 7422
rect 19068 7474 19124 8316
rect 19068 7422 19070 7474
rect 19122 7422 19124 7474
rect 19068 7410 19124 7422
rect 19180 8146 19236 8652
rect 19740 8258 19796 8876
rect 19740 8206 19742 8258
rect 19794 8206 19796 8258
rect 19740 8194 19796 8206
rect 19852 8260 19908 9100
rect 20076 8708 20132 8718
rect 20076 8370 20132 8652
rect 21196 8708 21252 10446
rect 21644 9940 21700 11314
rect 21868 10388 21924 11788
rect 22316 11620 22372 11630
rect 22316 11526 22372 11564
rect 22428 11508 22484 11518
rect 21980 10612 22036 10622
rect 22428 10612 22484 11452
rect 22652 10836 22708 12014
rect 22876 10948 22932 12348
rect 23660 11844 23716 11854
rect 23660 11284 23716 11788
rect 23640 11228 23716 11284
rect 22876 10892 23492 10948
rect 22652 10770 22708 10780
rect 22764 10612 22820 10622
rect 21980 10610 22316 10612
rect 21980 10558 21982 10610
rect 22034 10558 22316 10610
rect 21980 10556 22316 10558
rect 21980 10546 22036 10556
rect 22260 10442 22316 10556
rect 22428 10610 22820 10612
rect 22428 10558 22430 10610
rect 22482 10558 22766 10610
rect 22818 10558 22820 10610
rect 22428 10556 22820 10558
rect 22428 10546 22484 10556
rect 22764 10546 22820 10556
rect 22260 10390 22262 10442
rect 22314 10390 22316 10442
rect 21868 10332 22036 10388
rect 22260 10378 22316 10390
rect 21308 9828 21364 9838
rect 21308 9746 21310 9772
rect 21362 9746 21364 9772
rect 21308 9734 21364 9746
rect 21196 8642 21252 8652
rect 21532 8930 21588 8942
rect 21532 8878 21534 8930
rect 21586 8878 21588 8930
rect 20076 8318 20078 8370
rect 20130 8318 20132 8370
rect 20076 8306 20132 8318
rect 20300 8260 20356 8270
rect 19852 8228 19964 8260
rect 19852 8204 19910 8228
rect 19908 8176 19910 8204
rect 19962 8176 19964 8228
rect 19908 8164 19964 8176
rect 20188 8258 20356 8260
rect 20188 8206 20302 8258
rect 20354 8206 20356 8258
rect 20188 8204 20356 8206
rect 19180 8094 19182 8146
rect 19234 8094 19236 8146
rect 18956 7364 19012 7374
rect 18620 6972 18900 7028
rect 18508 6850 18564 6860
rect 18620 6804 18676 6814
rect 18508 6580 18564 6590
rect 18396 6578 18564 6580
rect 18396 6526 18510 6578
rect 18562 6526 18564 6578
rect 18396 6524 18564 6526
rect 18396 6132 18452 6524
rect 18508 6514 18564 6524
rect 18396 6066 18452 6076
rect 18620 6244 18676 6748
rect 18620 6020 18676 6188
rect 18508 5964 18676 6020
rect 18508 5950 18564 5964
rect 17836 5842 17892 5852
rect 18284 5906 18340 5918
rect 18284 5854 18286 5906
rect 18338 5854 18340 5906
rect 18508 5898 18510 5950
rect 18562 5898 18564 5950
rect 18508 5886 18564 5898
rect 17836 5684 17892 5694
rect 17836 5122 17892 5628
rect 18284 5236 18340 5854
rect 18620 5796 18676 5806
rect 18620 5702 18676 5740
rect 18284 5170 18340 5180
rect 17836 5070 17838 5122
rect 17890 5070 17892 5122
rect 17836 5058 17892 5070
rect 17948 5122 18004 5134
rect 17948 5070 17950 5122
rect 18002 5070 18004 5122
rect 17948 4564 18004 5070
rect 17612 4286 17614 4338
rect 17666 4286 17668 4338
rect 17612 4274 17668 4286
rect 17836 4508 18004 4564
rect 18060 5124 18116 5134
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17332 3780 17388 3790
rect 17836 3780 17892 4508
rect 17948 4353 18004 4378
rect 17948 4340 17950 4353
rect 18002 4340 18004 4353
rect 17948 4274 18004 4284
rect 18060 4226 18116 5068
rect 18732 5124 18788 5134
rect 18732 5030 18788 5068
rect 18284 5012 18340 5022
rect 18284 4340 18340 4956
rect 18844 4564 18900 6972
rect 18956 6690 19012 7308
rect 18956 6638 18958 6690
rect 19010 6638 19012 6690
rect 18956 5906 19012 6638
rect 19068 6692 19124 6702
rect 19180 6692 19236 8094
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20188 7700 20244 8204
rect 20300 8194 20356 8204
rect 21532 8260 21588 8878
rect 21532 8194 21588 8204
rect 20636 8036 20692 8046
rect 20636 8034 21588 8036
rect 20636 7982 20638 8034
rect 20690 7982 21588 8034
rect 20636 7980 21588 7982
rect 20636 7970 20692 7980
rect 20076 7644 20244 7700
rect 19852 7364 19908 7374
rect 19124 6636 19236 6692
rect 19292 7362 19908 7364
rect 19292 7310 19854 7362
rect 19906 7310 19908 7362
rect 19292 7308 19908 7310
rect 19068 6626 19124 6636
rect 19292 6580 19348 7308
rect 19852 7298 19908 7308
rect 20076 7140 20132 7644
rect 20076 7084 20244 7140
rect 19516 6690 19572 6702
rect 19516 6638 19518 6690
rect 19570 6638 19572 6690
rect 19292 6524 19460 6580
rect 19124 6468 19180 6478
rect 19124 6466 19236 6468
rect 19124 6414 19126 6466
rect 19178 6414 19236 6466
rect 19124 6402 19236 6414
rect 18956 5854 18958 5906
rect 19010 5854 19012 5906
rect 18956 5842 19012 5854
rect 19180 5572 19236 6402
rect 19292 6244 19348 6254
rect 19292 5950 19348 6188
rect 19292 5898 19294 5950
rect 19346 5898 19348 5950
rect 19292 5886 19348 5898
rect 19404 5794 19460 6524
rect 19516 5908 19572 6638
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19516 5842 19572 5852
rect 19628 5906 19684 5918
rect 19628 5854 19630 5906
rect 19682 5854 19684 5906
rect 19404 5742 19406 5794
rect 19458 5742 19460 5794
rect 19404 5730 19460 5742
rect 19628 5572 19684 5854
rect 19180 5516 19684 5572
rect 20188 5012 20244 7084
rect 20636 6692 20692 6702
rect 20392 6634 20448 6646
rect 20392 6582 20394 6634
rect 20446 6582 20448 6634
rect 20636 6598 20692 6636
rect 20392 6580 20448 6582
rect 20392 6514 20448 6524
rect 20636 6020 20692 6030
rect 20412 5796 20468 5806
rect 20412 5702 20468 5740
rect 20636 5234 20692 5964
rect 21532 5348 21588 7980
rect 21644 6662 21700 9884
rect 21980 9069 22036 10332
rect 23436 10164 23492 10892
rect 23640 10666 23696 11228
rect 23640 10614 23642 10666
rect 23694 10614 23696 10666
rect 23640 10602 23696 10614
rect 23772 10500 23828 12796
rect 23884 12786 23940 12796
rect 25228 12292 25284 14476
rect 25564 15092 25732 15148
rect 25788 15316 25844 15326
rect 25340 12740 25396 12750
rect 25340 12646 25396 12684
rect 25228 12198 25284 12236
rect 25396 12122 25452 12134
rect 24556 12066 24612 12078
rect 24556 12014 24558 12066
rect 24610 12014 24612 12066
rect 24556 11844 24612 12014
rect 25396 12070 25398 12122
rect 25450 12070 25452 12122
rect 24556 11778 24612 11788
rect 24780 11956 24836 11966
rect 24668 11506 24724 11518
rect 24668 11454 24670 11506
rect 24722 11454 24724 11506
rect 24332 11396 24388 11406
rect 23884 11394 24388 11396
rect 23884 11342 24334 11394
rect 24386 11342 24388 11394
rect 23884 11340 24388 11342
rect 23884 10722 23940 11340
rect 24332 11330 24388 11340
rect 24556 11338 24612 11350
rect 24556 11286 24558 11338
rect 24610 11286 24612 11338
rect 24444 10836 24500 10846
rect 24444 10742 24500 10780
rect 23884 10670 23886 10722
rect 23938 10670 23940 10722
rect 23884 10658 23940 10670
rect 23212 10108 23492 10164
rect 23660 10444 23828 10500
rect 22316 10052 22372 10062
rect 22316 9958 22372 9996
rect 21980 9017 21982 9069
rect 22034 9017 22036 9069
rect 21980 9005 22036 9017
rect 23212 8148 23268 10108
rect 23436 9940 23492 9950
rect 23324 9268 23380 9278
rect 23324 9174 23380 9212
rect 23192 8092 23268 8148
rect 23324 8148 23380 8158
rect 22092 8034 22148 8046
rect 22092 7982 22094 8034
rect 22146 7982 22148 8034
rect 21756 7364 21812 7374
rect 21756 7270 21812 7308
rect 22092 6804 22148 7982
rect 23192 7530 23248 8092
rect 22316 7476 22372 7514
rect 23192 7478 23194 7530
rect 23246 7478 23248 7530
rect 23192 7466 23248 7478
rect 22316 7410 22372 7420
rect 22316 6916 22372 6926
rect 22316 6822 22372 6860
rect 22092 6738 22148 6748
rect 21644 6610 21646 6662
rect 21698 6610 21700 6662
rect 21644 6598 21700 6610
rect 20636 5182 20638 5234
rect 20690 5182 20692 5234
rect 20636 5170 20692 5182
rect 21196 5292 21588 5348
rect 22316 5908 22372 5918
rect 22316 5794 22372 5852
rect 23212 5908 23268 5918
rect 23324 5908 23380 8092
rect 23436 7586 23492 9884
rect 23436 7534 23438 7586
rect 23490 7534 23492 7586
rect 23436 7522 23492 7534
rect 23660 6580 23716 10444
rect 24556 10276 24612 11286
rect 24668 10276 24724 11454
rect 24780 10610 24836 11900
rect 25396 11844 25452 12070
rect 25396 11778 25452 11788
rect 25340 11620 25396 11630
rect 24780 10558 24782 10610
rect 24834 10558 24836 10610
rect 24780 10546 24836 10558
rect 24892 11394 24948 11406
rect 24892 11342 24894 11394
rect 24946 11342 24948 11394
rect 24668 10220 24836 10276
rect 24556 10210 24612 10220
rect 24780 10164 24836 10220
rect 24780 10098 24836 10108
rect 24892 9940 24948 11342
rect 25340 10724 25396 11564
rect 24780 9884 24948 9940
rect 25004 10722 25396 10724
rect 25004 10670 25342 10722
rect 25394 10670 25396 10722
rect 25004 10668 25396 10670
rect 24108 9826 24164 9838
rect 24108 9774 24110 9826
rect 24162 9774 24164 9826
rect 24108 9716 24164 9774
rect 24108 9650 24164 9660
rect 24780 8484 24836 9884
rect 25004 9838 25060 10668
rect 25340 10658 25396 10668
rect 24984 9826 25060 9838
rect 24984 9774 24986 9826
rect 25038 9774 25060 9826
rect 24984 9772 25060 9774
rect 25452 10052 25508 10062
rect 24984 9762 25040 9772
rect 25228 9714 25284 9726
rect 25228 9662 25230 9714
rect 25282 9662 25284 9714
rect 25228 9268 25284 9662
rect 24780 8418 24836 8428
rect 25116 9212 25284 9268
rect 23996 8260 24052 8270
rect 24108 8260 24164 8270
rect 23660 6514 23716 6524
rect 23772 8230 23828 8242
rect 23772 8178 23774 8230
rect 23826 8178 23828 8230
rect 24052 8258 24164 8260
rect 24052 8206 24110 8258
rect 24162 8206 24164 8258
rect 24052 8204 24164 8206
rect 23996 8194 24052 8204
rect 24108 8194 24164 8204
rect 24220 8260 24276 8270
rect 23772 6244 23828 8178
rect 24220 6802 24276 8204
rect 24984 8260 25040 8270
rect 24984 8166 25040 8204
rect 24220 6750 24222 6802
rect 24274 6750 24276 6802
rect 24220 6738 24276 6750
rect 24108 6690 24164 6702
rect 24108 6638 24110 6690
rect 24162 6638 24164 6690
rect 24108 6580 24164 6638
rect 24444 6692 24500 6702
rect 24780 6692 24836 6702
rect 24444 6611 24446 6636
rect 24498 6611 24500 6636
rect 24444 6598 24500 6611
rect 24556 6690 24836 6692
rect 24556 6638 24782 6690
rect 24834 6638 24836 6690
rect 24556 6636 24836 6638
rect 24108 6514 24164 6524
rect 24444 6468 24500 6478
rect 23772 6188 24164 6244
rect 23212 5906 23380 5908
rect 23212 5854 23214 5906
rect 23266 5854 23380 5906
rect 23212 5852 23380 5854
rect 23436 5908 23492 5946
rect 23212 5842 23268 5852
rect 23436 5842 23492 5852
rect 22316 5742 22318 5794
rect 22370 5742 22372 5794
rect 20188 4946 20244 4956
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18844 4508 19908 4564
rect 18060 4174 18062 4226
rect 18114 4174 18116 4226
rect 18060 4162 18116 4174
rect 18172 4338 18340 4340
rect 18172 4286 18286 4338
rect 18338 4286 18340 4338
rect 18172 4284 18340 4286
rect 17332 3778 17892 3780
rect 17332 3726 17334 3778
rect 17386 3726 17892 3778
rect 17332 3724 17892 3726
rect 17332 3714 17388 3724
rect 17500 3556 17556 3566
rect 17500 3462 17556 3500
rect 18172 3554 18228 4284
rect 18284 4274 18340 4284
rect 18172 3502 18174 3554
rect 18226 3502 18228 3554
rect 18172 3490 18228 3502
rect 19516 4226 19572 4238
rect 19516 4174 19518 4226
rect 19570 4174 19572 4226
rect 19516 4116 19572 4174
rect 19516 3556 19572 4060
rect 19516 3490 19572 3500
rect 19852 3526 19908 4508
rect 21196 4004 21252 5292
rect 22316 5236 22372 5742
rect 22876 5684 22932 5694
rect 22316 5170 22372 5180
rect 22540 5682 22932 5684
rect 22540 5630 22878 5682
rect 22930 5630 22932 5682
rect 22540 5628 22932 5630
rect 22540 5234 22596 5628
rect 22876 5618 22932 5628
rect 22540 5182 22542 5234
rect 22594 5182 22596 5234
rect 22540 5170 22596 5182
rect 21532 5124 21588 5134
rect 21532 5030 21588 5068
rect 21756 5124 21812 5134
rect 21756 5030 21812 5068
rect 21364 4900 21420 4910
rect 21364 4806 21420 4844
rect 22204 4900 22260 4910
rect 22204 4338 22260 4844
rect 22876 4564 22932 4574
rect 22204 4286 22206 4338
rect 22258 4286 22260 4338
rect 22204 4274 22260 4286
rect 22540 4353 22596 4365
rect 22540 4340 22542 4353
rect 22594 4340 22596 4353
rect 21420 4228 21476 4238
rect 21420 4134 21476 4172
rect 22428 4228 22484 4238
rect 22428 4134 22484 4172
rect 19852 3474 19854 3526
rect 19906 3474 19908 3526
rect 19852 3462 19908 3474
rect 21084 3948 21252 4004
rect 21084 3526 21140 3948
rect 22540 3780 22596 4284
rect 22876 4338 22932 4508
rect 22876 4286 22878 4338
rect 22930 4286 22932 4338
rect 22876 4116 22932 4286
rect 22876 4050 22932 4060
rect 22540 3714 22596 3724
rect 21084 3474 21086 3526
rect 21138 3474 21140 3526
rect 21084 3462 21140 3474
rect 22988 3556 23044 3566
rect 22988 3462 23044 3500
rect 24108 3556 24164 6188
rect 24312 5908 24368 5918
rect 24312 5906 24388 5908
rect 24312 5854 24314 5906
rect 24366 5854 24388 5906
rect 24312 5842 24388 5854
rect 24332 4452 24388 5842
rect 24444 5234 24500 6412
rect 24556 6018 24612 6636
rect 24780 6626 24836 6636
rect 25116 6690 25172 9212
rect 25340 9044 25396 9054
rect 25452 9044 25508 9996
rect 25564 9210 25620 15092
rect 25676 12964 25732 12974
rect 25788 12964 25844 15260
rect 25676 12962 25844 12964
rect 25676 12910 25678 12962
rect 25730 12910 25844 12962
rect 25676 12908 25844 12910
rect 25676 12898 25732 12908
rect 25900 12404 25956 15484
rect 26012 16660 26068 16670
rect 26012 15204 26068 16604
rect 26124 16324 26180 17612
rect 26236 16660 26292 19740
rect 26964 19740 27300 19796
rect 26964 19458 27020 19740
rect 27468 19460 27524 19966
rect 28140 20020 28196 20030
rect 27636 19796 27692 19806
rect 27636 19794 27860 19796
rect 27636 19742 27638 19794
rect 27690 19742 27860 19794
rect 27636 19740 27860 19742
rect 27636 19730 27692 19740
rect 26964 19406 26966 19458
rect 27018 19406 27020 19458
rect 26964 19394 27020 19406
rect 27356 19404 27524 19460
rect 26908 19236 26964 19246
rect 26460 19122 26516 19134
rect 26460 19070 26462 19122
rect 26514 19070 26516 19122
rect 26460 18228 26516 19070
rect 26908 18676 26964 19180
rect 26796 18620 26964 18676
rect 27244 19234 27300 19246
rect 27244 19182 27246 19234
rect 27298 19182 27300 19234
rect 26572 18452 26628 18462
rect 26572 18358 26628 18396
rect 26796 18340 26852 18620
rect 27020 18452 27076 18462
rect 27244 18452 27300 19182
rect 27020 18450 27300 18452
rect 27020 18398 27022 18450
rect 27074 18398 27300 18450
rect 27020 18396 27300 18398
rect 27020 18386 27076 18396
rect 26796 18246 26852 18284
rect 26460 18162 26516 18172
rect 27244 18228 27300 18396
rect 27244 18162 27300 18172
rect 27356 18452 27412 19404
rect 27468 19236 27524 19246
rect 27804 19236 27860 19740
rect 27468 19234 27860 19236
rect 27468 19182 27470 19234
rect 27522 19182 27806 19234
rect 27858 19182 27860 19234
rect 27468 19180 27860 19182
rect 27468 19170 27524 19180
rect 27804 19170 27860 19180
rect 28028 19190 28084 19202
rect 28028 19138 28030 19190
rect 28082 19138 28084 19190
rect 27916 19066 27972 19078
rect 27916 19014 27918 19066
rect 27970 19014 27972 19066
rect 26236 16594 26292 16604
rect 26572 18116 26628 18126
rect 26292 16324 26348 16334
rect 26124 16322 26348 16324
rect 26124 16270 26294 16322
rect 26346 16270 26348 16322
rect 26124 16268 26348 16270
rect 26292 16258 26348 16268
rect 26572 16098 26628 18060
rect 27132 18004 27188 18014
rect 27020 17556 27076 17566
rect 26908 16884 26964 16894
rect 26908 16790 26964 16828
rect 26908 16660 26964 16670
rect 26572 16046 26574 16098
rect 26626 16046 26628 16098
rect 26572 16034 26628 16046
rect 26796 16100 26852 16110
rect 26796 16006 26852 16044
rect 26908 16100 26964 16604
rect 27020 16266 27076 17500
rect 27020 16214 27022 16266
rect 27074 16214 27076 16266
rect 27020 16202 27076 16214
rect 26908 16034 26964 16044
rect 27132 16098 27188 17948
rect 27244 17668 27300 17678
rect 27356 17668 27412 18396
rect 27804 18450 27860 18462
rect 27804 18398 27806 18450
rect 27858 18398 27860 18450
rect 27804 18340 27860 18398
rect 27804 18274 27860 18284
rect 27244 17666 27412 17668
rect 27244 17614 27246 17666
rect 27298 17614 27412 17666
rect 27580 18116 27636 18126
rect 27580 17778 27636 18060
rect 27916 18004 27972 19014
rect 28028 18676 28084 19138
rect 28140 18900 28196 19964
rect 28140 18834 28196 18844
rect 28252 20018 28308 20030
rect 28252 19966 28254 20018
rect 28306 19966 28308 20018
rect 28028 18620 28196 18676
rect 27916 17938 27972 17948
rect 28028 18489 28084 18501
rect 28028 18437 28030 18489
rect 28082 18437 28084 18489
rect 27580 17726 27582 17778
rect 27634 17726 27636 17778
rect 27244 17612 27412 17614
rect 27244 17108 27300 17612
rect 27244 17042 27300 17052
rect 27468 17610 27524 17622
rect 27468 17558 27470 17610
rect 27522 17558 27524 17610
rect 27468 17006 27524 17558
rect 27465 16996 27524 17006
rect 27521 16940 27524 16996
rect 27465 16921 27521 16940
rect 27244 16882 27300 16894
rect 27244 16830 27246 16882
rect 27298 16830 27300 16882
rect 27465 16869 27467 16921
rect 27519 16869 27521 16921
rect 27465 16857 27521 16869
rect 27244 16212 27300 16830
rect 27580 16772 27636 17726
rect 27916 17666 27972 17678
rect 27916 17614 27918 17666
rect 27970 17614 27972 17666
rect 27916 17108 27972 17614
rect 27916 17042 27972 17052
rect 28028 16996 28084 18437
rect 28140 18228 28196 18620
rect 28252 18564 28308 19966
rect 28364 19684 28420 20134
rect 28364 19618 28420 19628
rect 28588 19236 28644 20188
rect 28476 19180 28644 19236
rect 28700 20057 28756 20069
rect 28700 20005 28702 20057
rect 28754 20005 28756 20057
rect 28700 19236 28756 20005
rect 28812 19460 28868 21532
rect 28924 20132 28980 20142
rect 28924 20018 28980 20076
rect 28924 19966 28926 20018
rect 28978 19966 28980 20018
rect 28924 19954 28980 19966
rect 29036 20020 29092 23130
rect 29148 22482 29204 23660
rect 29260 23210 29316 23772
rect 29260 23158 29262 23210
rect 29314 23158 29316 23210
rect 29260 23146 29316 23158
rect 29372 23156 29428 23166
rect 29148 22430 29150 22482
rect 29202 22430 29204 22482
rect 29148 22418 29204 22430
rect 29260 22326 29316 22338
rect 29260 22274 29262 22326
rect 29314 22274 29316 22326
rect 29260 21924 29316 22274
rect 29260 21858 29316 21868
rect 29204 21700 29260 21710
rect 29372 21700 29428 23100
rect 29540 22930 29596 22942
rect 29540 22878 29542 22930
rect 29594 22878 29596 22930
rect 29540 22596 29596 22878
rect 29540 22530 29596 22540
rect 29596 22370 29652 22382
rect 29596 22318 29598 22370
rect 29650 22318 29652 22370
rect 29596 22036 29652 22318
rect 29708 22148 29764 24434
rect 30492 24276 30548 31052
rect 31612 31050 31668 32284
rect 31982 32246 32038 32284
rect 32396 32338 32452 32350
rect 32396 32286 32398 32338
rect 32450 32286 32452 32338
rect 32396 32116 32452 32286
rect 32396 32050 32452 32060
rect 32956 32340 33012 32350
rect 31836 31778 31892 31790
rect 31836 31726 31838 31778
rect 31890 31726 31892 31778
rect 30604 30994 30660 31006
rect 30604 30942 30606 30994
rect 30658 30942 30660 30994
rect 30604 30884 30660 30942
rect 30604 30818 30660 30828
rect 30828 30994 30884 31006
rect 30828 30942 30830 30994
rect 30882 30942 30884 30994
rect 30828 30884 30884 30942
rect 31108 30996 31164 31006
rect 31612 30998 31614 31050
rect 31666 30998 31668 31050
rect 31612 30986 31668 30998
rect 31724 31108 31780 31118
rect 31724 31050 31780 31052
rect 31724 30998 31726 31050
rect 31778 30998 31780 31050
rect 31724 30986 31780 30998
rect 31108 30902 31164 30940
rect 30828 30436 30884 30828
rect 31836 30884 31892 31726
rect 31948 31780 32004 31790
rect 31948 31050 32004 31724
rect 32172 31780 32228 31790
rect 32172 31686 32228 31724
rect 32732 31778 32788 31790
rect 32732 31726 32734 31778
rect 32786 31726 32788 31778
rect 31948 30998 31950 31050
rect 32002 30998 32004 31050
rect 32732 31108 32788 31726
rect 32956 31778 33012 32284
rect 33404 32340 33460 32510
rect 33404 32274 33460 32284
rect 33572 32340 33628 32350
rect 33572 32338 33684 32340
rect 33572 32286 33574 32338
rect 33626 32286 33684 32338
rect 33572 32274 33684 32286
rect 33180 31892 33236 31902
rect 33628 31892 33684 32274
rect 33852 32004 33908 34114
rect 34524 33796 34580 36204
rect 34692 36036 34748 36374
rect 34692 35970 34748 35980
rect 34692 35812 34748 35822
rect 34692 35718 34748 35756
rect 34972 35698 35028 35710
rect 34972 35646 34974 35698
rect 35026 35646 35028 35698
rect 34972 35476 35028 35646
rect 34972 35410 35028 35420
rect 35084 34914 35140 36540
rect 35196 36372 35252 36382
rect 35196 35698 35252 36316
rect 35196 35646 35198 35698
rect 35250 35646 35252 35698
rect 35196 35634 35252 35646
rect 35476 35700 35532 35710
rect 36988 35700 37044 36988
rect 35476 35606 35532 35644
rect 36876 35644 37044 35700
rect 37212 36454 37268 36466
rect 37212 36402 37214 36454
rect 37266 36402 37268 36454
rect 35532 35476 35588 35486
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35084 34862 35086 34914
rect 35138 34862 35140 34914
rect 35084 34850 35140 34862
rect 34636 34132 34692 34142
rect 34636 33962 34692 34076
rect 34636 33910 34638 33962
rect 34690 33910 34692 33962
rect 34636 33898 34692 33910
rect 34748 34130 34804 34142
rect 34748 34078 34750 34130
rect 34802 34078 34804 34130
rect 34748 33796 34804 34078
rect 35084 34130 35140 34142
rect 35084 34078 35086 34130
rect 35138 34078 35140 34130
rect 35084 33908 35140 34078
rect 35308 34132 35364 34142
rect 35532 34132 35588 35420
rect 35924 35476 35980 35486
rect 35756 35140 35812 35150
rect 35308 34130 35588 34132
rect 35308 34078 35310 34130
rect 35362 34078 35588 34130
rect 35308 34076 35588 34078
rect 35644 34914 35700 34926
rect 35644 34862 35646 34914
rect 35698 34862 35700 34914
rect 35308 34066 35364 34076
rect 35084 33842 35140 33852
rect 35644 33906 35700 34862
rect 35756 34914 35812 35084
rect 35756 34862 35758 34914
rect 35810 34862 35812 34914
rect 35756 34850 35812 34862
rect 35924 34914 35980 35420
rect 36876 35252 36932 35644
rect 37044 35476 37100 35486
rect 37044 35382 37100 35420
rect 36876 35196 37044 35252
rect 36316 35028 36372 35038
rect 36316 35026 36708 35028
rect 36316 34974 36318 35026
rect 36370 34974 36708 35026
rect 36316 34972 36708 34974
rect 36316 34962 36372 34972
rect 35924 34862 35926 34914
rect 35978 34862 35980 34914
rect 35924 34850 35980 34862
rect 36484 33908 36540 33918
rect 35644 33854 35646 33906
rect 35698 33854 35700 33906
rect 34188 33740 34804 33796
rect 35196 33740 35460 33750
rect 34020 32676 34076 32686
rect 34020 32582 34076 32620
rect 34076 32004 34132 32014
rect 33852 32002 34132 32004
rect 33852 31950 34078 32002
rect 34130 31950 34132 32002
rect 33852 31948 34132 31950
rect 34076 31938 34132 31948
rect 33740 31892 33796 31902
rect 33180 31890 33460 31892
rect 33180 31838 33182 31890
rect 33234 31838 33460 31890
rect 33180 31836 33460 31838
rect 33628 31836 33740 31892
rect 33180 31826 33236 31836
rect 32956 31726 32958 31778
rect 33010 31726 33012 31778
rect 32956 31714 33012 31726
rect 33404 31778 33460 31836
rect 33740 31826 33796 31836
rect 33404 31726 33406 31778
rect 33458 31726 33460 31778
rect 33404 31714 33460 31726
rect 33516 31778 33572 31790
rect 33516 31726 33518 31778
rect 33570 31726 33572 31778
rect 32732 31042 32788 31052
rect 31948 30986 32004 30998
rect 32172 31022 32228 31034
rect 31836 30818 31892 30828
rect 32172 30970 32174 31022
rect 32226 30970 32228 31022
rect 32172 30884 32228 30970
rect 32172 30818 32228 30828
rect 32284 30996 32340 31006
rect 30828 30370 30884 30380
rect 31612 30212 31668 30222
rect 31612 29764 31668 30156
rect 32284 29764 32340 30940
rect 33068 30994 33124 31006
rect 33068 30942 33070 30994
rect 33122 30942 33124 30994
rect 32452 30772 32508 30782
rect 32452 30770 33012 30772
rect 32452 30718 32454 30770
rect 32506 30718 33012 30770
rect 32452 30716 33012 30718
rect 32452 30706 32508 30716
rect 32732 30436 32788 30446
rect 32732 30342 32788 30380
rect 32488 30154 32544 30166
rect 32488 30102 32490 30154
rect 32542 30102 32544 30154
rect 32488 29764 32544 30102
rect 32956 29988 33012 30716
rect 33068 30212 33124 30942
rect 33180 30996 33236 31006
rect 33180 30902 33236 30940
rect 33348 30996 33404 31006
rect 33348 30902 33404 30940
rect 33516 30436 33572 31726
rect 33684 31722 33740 31734
rect 33684 31670 33686 31722
rect 33738 31670 33740 31722
rect 33684 31108 33740 31670
rect 34188 31220 34244 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35084 33572 35140 33582
rect 34860 33346 34916 33358
rect 34412 33318 34468 33330
rect 34412 33266 34414 33318
rect 34466 33266 34468 33318
rect 34412 33124 34468 33266
rect 34860 33294 34862 33346
rect 34914 33294 34916 33346
rect 34412 33058 34468 33068
rect 34748 33236 34804 33246
rect 34580 32900 34636 32910
rect 34580 32618 34636 32844
rect 34300 32562 34356 32574
rect 34300 32510 34302 32562
rect 34354 32510 34356 32562
rect 34300 32340 34356 32510
rect 34300 32274 34356 32284
rect 34412 32562 34468 32574
rect 34412 32510 34414 32562
rect 34466 32510 34468 32562
rect 34580 32566 34582 32618
rect 34634 32566 34636 32618
rect 34580 32554 34636 32566
rect 34748 32618 34804 33180
rect 34748 32566 34750 32618
rect 34802 32566 34804 32618
rect 34748 32554 34804 32566
rect 34076 31164 34244 31220
rect 34300 32116 34356 32126
rect 33684 31052 33796 31108
rect 33740 30996 33796 31052
rect 33852 30996 33908 31006
rect 33740 30940 33852 30996
rect 33740 30772 33796 30782
rect 33740 30678 33796 30716
rect 33516 30370 33572 30380
rect 33852 30434 33908 30940
rect 33852 30382 33854 30434
rect 33906 30382 33908 30434
rect 33852 30370 33908 30382
rect 33068 30146 33124 30156
rect 33180 30210 33236 30222
rect 33180 30158 33182 30210
rect 33234 30158 33236 30210
rect 33180 29988 33236 30158
rect 32956 29932 33236 29988
rect 33292 30210 33348 30222
rect 33292 30158 33294 30210
rect 33346 30158 33348 30210
rect 31612 29708 32004 29764
rect 31276 29428 31332 29438
rect 31052 29426 31332 29428
rect 31052 29374 31278 29426
rect 31330 29374 31332 29426
rect 31052 29372 31332 29374
rect 31052 28810 31108 29372
rect 31276 29362 31332 29372
rect 31948 28878 32004 29708
rect 32284 29708 32544 29764
rect 32152 29428 32208 29438
rect 32284 29428 32340 29708
rect 33292 29652 33348 30158
rect 33460 30212 33516 30222
rect 34076 30212 34132 31164
rect 34188 30996 34244 31006
rect 34188 30902 34244 30940
rect 34300 30660 34356 32060
rect 34412 30826 34468 32510
rect 34860 32452 34916 33294
rect 34636 32396 34916 32452
rect 34972 33348 35028 33358
rect 34972 32562 35028 33292
rect 34972 32510 34974 32562
rect 35026 32510 35028 32562
rect 34636 32014 34692 32396
rect 34972 32340 35028 32510
rect 34580 32002 34692 32014
rect 34580 31950 34582 32002
rect 34634 31950 34692 32002
rect 34580 31948 34692 31950
rect 34748 32284 35028 32340
rect 34580 31938 34636 31948
rect 34412 30774 34414 30826
rect 34466 30774 34468 30826
rect 34412 30762 34468 30774
rect 34524 30994 34580 31006
rect 34524 30942 34526 30994
rect 34578 30942 34580 30994
rect 34524 30660 34580 30942
rect 34748 30996 34804 32284
rect 35084 32228 35140 33516
rect 35532 33346 35588 33358
rect 35532 33294 35534 33346
rect 35586 33294 35588 33346
rect 35196 33122 35252 33134
rect 35196 33070 35198 33122
rect 35250 33070 35252 33122
rect 35196 32452 35252 33070
rect 35532 32676 35588 33294
rect 35532 32610 35588 32620
rect 35644 32900 35700 33854
rect 35980 33906 36540 33908
rect 35980 33854 36486 33906
rect 36538 33854 36540 33906
rect 35980 33852 36540 33854
rect 35196 32386 35252 32396
rect 35644 32564 35700 32844
rect 35868 33122 35924 33134
rect 35868 33070 35870 33122
rect 35922 33070 35924 33122
rect 34972 32172 35140 32228
rect 35196 32172 35460 32182
rect 34860 31892 34916 31902
rect 34860 31778 34916 31836
rect 34860 31726 34862 31778
rect 34914 31726 34916 31778
rect 34860 31714 34916 31726
rect 34972 31778 35028 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35644 32116 35700 32508
rect 35756 32564 35812 32574
rect 35868 32564 35924 33070
rect 35756 32562 35924 32564
rect 35756 32510 35758 32562
rect 35810 32510 35924 32562
rect 35756 32508 35924 32510
rect 35756 32498 35812 32508
rect 35196 32106 35460 32116
rect 35532 32060 35700 32116
rect 35868 32340 35924 32350
rect 35532 32004 35588 32060
rect 34972 31726 34974 31778
rect 35026 31726 35028 31778
rect 35140 31948 35588 32004
rect 35756 32004 35812 32014
rect 35140 31834 35196 31948
rect 35140 31782 35142 31834
rect 35194 31782 35196 31834
rect 35140 31770 35196 31782
rect 35308 31780 35364 31790
rect 34972 31714 35028 31726
rect 35308 31686 35364 31724
rect 35532 31778 35588 31790
rect 35532 31726 35534 31778
rect 35586 31726 35588 31778
rect 34972 30996 35028 31006
rect 34748 30994 35028 30996
rect 34748 30942 34974 30994
rect 35026 30942 35028 30994
rect 34748 30940 35028 30942
rect 34972 30930 35028 30940
rect 35532 30996 35588 31726
rect 35644 31780 35700 31790
rect 35644 30996 35700 31724
rect 35756 31778 35812 31948
rect 35756 31726 35758 31778
rect 35810 31726 35812 31778
rect 35756 31714 35812 31726
rect 35868 31668 35924 32284
rect 35980 31892 36036 33852
rect 36484 33842 36540 33852
rect 36484 33124 36540 33134
rect 36484 32788 36540 33068
rect 36652 33012 36708 34972
rect 36988 34186 37044 35196
rect 37100 35028 37156 35038
rect 37100 34934 37156 34972
rect 37212 34356 37268 36402
rect 37212 34290 37268 34300
rect 37324 35726 37380 35738
rect 37324 35674 37326 35726
rect 37378 35674 37380 35726
rect 37324 35028 37380 35674
rect 36764 34158 36820 34170
rect 36764 34106 36766 34158
rect 36818 34106 36820 34158
rect 36764 33572 36820 34106
rect 36764 33506 36820 33516
rect 36988 34134 36990 34186
rect 37042 34134 37044 34186
rect 37324 34186 37380 34972
rect 36988 33460 37044 34134
rect 37212 34158 37268 34170
rect 37212 34132 37214 34158
rect 37266 34132 37268 34158
rect 37324 34134 37326 34186
rect 37378 34134 37380 34186
rect 37324 34122 37380 34134
rect 37436 34132 37492 37212
rect 37884 37268 37940 37278
rect 37884 37174 37940 37212
rect 38220 37268 38276 37278
rect 37548 37044 37604 37054
rect 37548 35754 37604 36988
rect 38220 37042 38276 37212
rect 39228 37268 39284 37278
rect 39228 37174 39284 37212
rect 38220 36990 38222 37042
rect 38274 36990 38276 37042
rect 38220 36820 38276 36990
rect 39340 37044 39396 38556
rect 39564 38388 39620 38838
rect 39788 38862 39844 38874
rect 39788 38810 39790 38862
rect 39842 38810 39844 38862
rect 39788 38612 39844 38810
rect 39788 38546 39844 38556
rect 39452 38332 39620 38388
rect 39900 38388 39956 39564
rect 40012 40180 40068 40190
rect 40012 39590 40068 40124
rect 40292 39842 40348 40348
rect 40460 40338 40516 40348
rect 40796 40402 40852 40414
rect 40796 40350 40798 40402
rect 40850 40350 40852 40402
rect 40292 39790 40294 39842
rect 40346 39790 40348 39842
rect 40292 39778 40348 39790
rect 40572 39620 40628 39630
rect 40796 39620 40852 40350
rect 40012 39538 40014 39590
rect 40066 39538 40068 39590
rect 40012 39526 40068 39538
rect 40460 39618 40852 39620
rect 40460 39566 40574 39618
rect 40626 39566 40852 39618
rect 40460 39564 40852 39566
rect 40012 38862 40068 38874
rect 40012 38810 40014 38862
rect 40066 38810 40068 38862
rect 40012 38724 40068 38810
rect 40012 38658 40068 38668
rect 40292 38612 40348 38622
rect 40292 38518 40348 38556
rect 39900 38332 40404 38388
rect 39452 37492 39508 38332
rect 40348 37828 40404 38332
rect 40236 37772 40404 37828
rect 39564 37492 39620 37502
rect 40236 37492 40292 37772
rect 39452 37490 39620 37492
rect 39452 37438 39566 37490
rect 39618 37438 39620 37490
rect 39452 37436 39620 37438
rect 39564 37426 39620 37436
rect 40124 37490 40292 37492
rect 40124 37438 40238 37490
rect 40290 37438 40292 37490
rect 40124 37436 40292 37438
rect 39340 36978 39396 36988
rect 39900 37266 39956 37278
rect 39900 37214 39902 37266
rect 39954 37214 39956 37266
rect 39900 37044 39956 37214
rect 39900 36978 39956 36988
rect 37548 35702 37550 35754
rect 37602 35702 37604 35754
rect 37548 35690 37604 35702
rect 37772 36764 38276 36820
rect 37772 35754 37828 36764
rect 37996 36596 38052 36606
rect 37996 36502 38052 36540
rect 39788 36372 39844 36382
rect 37772 35702 37774 35754
rect 37826 35702 37828 35754
rect 37772 35690 37828 35702
rect 37884 36148 37940 36158
rect 37884 35754 37940 36092
rect 37884 35702 37886 35754
rect 37938 35702 37940 35754
rect 37884 35690 37940 35702
rect 39788 35698 39844 36316
rect 40012 35812 40068 35822
rect 39788 35646 39790 35698
rect 39842 35646 39844 35698
rect 39788 35634 39844 35646
rect 39900 35698 39956 35710
rect 39900 35646 39902 35698
rect 39954 35646 39956 35698
rect 39452 35588 39508 35598
rect 39452 35494 39508 35532
rect 39900 35140 39956 35646
rect 39564 35084 39956 35140
rect 39004 34914 39060 34926
rect 39004 34862 39006 34914
rect 39058 34862 39060 34914
rect 37884 34244 37940 34254
rect 37884 34157 37940 34188
rect 37212 34066 37268 34076
rect 37492 34076 37716 34132
rect 37884 34105 37886 34157
rect 37938 34105 37940 34157
rect 37884 34093 37940 34105
rect 37436 34066 37492 34076
rect 36988 33394 37044 33404
rect 37324 33908 37380 33918
rect 37324 33318 37380 33852
rect 37324 33266 37326 33318
rect 37378 33266 37380 33318
rect 37044 33236 37100 33246
rect 37044 33142 37100 33180
rect 37324 33124 37380 33266
rect 37548 33460 37604 33470
rect 37548 33318 37604 33404
rect 37548 33266 37550 33318
rect 37602 33266 37604 33318
rect 37660 33348 37716 34076
rect 38892 33906 38948 33918
rect 38892 33854 38894 33906
rect 38946 33854 38948 33906
rect 38332 33684 38388 33694
rect 37884 33572 37940 33582
rect 37660 33311 37772 33348
rect 37660 33292 37718 33311
rect 37548 33254 37604 33266
rect 37716 33259 37718 33292
rect 37770 33259 37772 33311
rect 37716 33247 37772 33259
rect 37884 33290 37940 33516
rect 37884 33238 37886 33290
rect 37938 33238 37940 33290
rect 38108 33348 38164 33358
rect 38108 33254 38164 33292
rect 37324 33068 37716 33124
rect 36652 32946 36708 32956
rect 36484 32732 36932 32788
rect 35980 31826 36036 31836
rect 36036 31668 36092 31678
rect 35868 31666 36092 31668
rect 35868 31614 36038 31666
rect 36090 31614 36092 31666
rect 35868 31612 36092 31614
rect 36036 31602 36092 31612
rect 35756 30996 35812 31006
rect 35644 30994 35812 30996
rect 35644 30942 35758 30994
rect 35810 30942 35812 30994
rect 35644 30940 35812 30942
rect 35532 30930 35588 30940
rect 35756 30930 35812 30940
rect 36876 30660 36932 32732
rect 37660 32674 37716 33068
rect 37660 32622 37662 32674
rect 37714 32622 37716 32674
rect 37660 32610 37716 32622
rect 37660 31108 37716 31118
rect 37884 31108 37940 33238
rect 37996 33012 38052 33022
rect 37996 32562 38052 32956
rect 38332 32786 38388 33628
rect 38892 33348 38948 33854
rect 39004 33684 39060 34862
rect 39004 33618 39060 33628
rect 38892 33282 38948 33292
rect 39452 33348 39508 33358
rect 39452 33254 39508 33292
rect 38332 32734 38334 32786
rect 38386 32734 38388 32786
rect 38332 32722 38388 32734
rect 38836 32788 38892 32798
rect 38836 32694 38892 32732
rect 39564 32686 39620 35084
rect 39788 34916 39844 34926
rect 39900 34916 39956 34926
rect 39788 34914 39956 34916
rect 39788 34862 39790 34914
rect 39842 34862 39902 34914
rect 39954 34862 39956 34914
rect 39788 34860 39956 34862
rect 39788 34132 39844 34860
rect 39900 34850 39956 34860
rect 39788 33348 39844 34076
rect 39788 33282 39844 33292
rect 40012 33124 40068 35756
rect 39508 32674 39620 32686
rect 39508 32622 39510 32674
rect 39562 32622 39620 32674
rect 39508 32620 39620 32622
rect 39788 33068 40068 33124
rect 40124 34244 40180 37436
rect 40236 37426 40292 37436
rect 40460 36708 40516 39564
rect 40572 39554 40628 39564
rect 40908 39508 40964 40572
rect 41020 40404 41076 41078
rect 41020 40338 41076 40348
rect 41244 41130 41300 41142
rect 41244 41078 41246 41130
rect 41298 41078 41300 41130
rect 41244 39620 41300 41078
rect 41356 41130 41412 41142
rect 41356 41078 41358 41130
rect 41410 41078 41412 41130
rect 41356 40180 41412 41078
rect 42028 41106 42030 41158
rect 42082 41106 42084 41158
rect 42028 40628 42084 41106
rect 42028 40562 42084 40572
rect 42812 40628 42868 40638
rect 41580 40292 41636 40302
rect 41580 40198 41636 40236
rect 41356 40114 41412 40124
rect 41356 39732 41412 39742
rect 41356 39638 41412 39676
rect 41244 39554 41300 39564
rect 40572 39396 40628 39406
rect 40572 38162 40628 39340
rect 40908 38836 40964 39452
rect 40908 38770 40964 38780
rect 41356 38836 41412 38846
rect 41020 38724 41076 38734
rect 41020 38630 41076 38668
rect 40572 38110 40574 38162
rect 40626 38110 40628 38162
rect 40572 38098 40628 38110
rect 41356 38050 41412 38780
rect 41356 37998 41358 38050
rect 41410 37998 41412 38050
rect 40908 37268 40964 37278
rect 41356 37268 41412 37998
rect 41580 38724 41636 38734
rect 41580 38015 41636 38668
rect 41580 37963 41582 38015
rect 41634 37963 41636 38015
rect 41916 38500 41972 38510
rect 41916 38022 41972 38444
rect 41580 37951 41636 37963
rect 41692 37994 41748 38006
rect 41692 37942 41694 37994
rect 41746 37942 41748 37994
rect 41916 37970 41918 38022
rect 41970 37970 41972 38022
rect 42420 38052 42476 38062
rect 42700 38052 42756 38062
rect 42420 38050 42756 38052
rect 41916 37958 41972 37970
rect 42140 37994 42196 38006
rect 41692 37492 41748 37942
rect 42140 37942 42142 37994
rect 42194 37942 42196 37994
rect 42420 37998 42422 38050
rect 42474 37998 42702 38050
rect 42754 37998 42756 38050
rect 42420 37996 42756 37998
rect 42420 37986 42476 37996
rect 42700 37986 42756 37996
rect 42140 37492 42196 37942
rect 40908 37266 41412 37268
rect 40908 37214 40910 37266
rect 40962 37214 41412 37266
rect 40908 37212 41412 37214
rect 41468 37436 41748 37492
rect 41916 37436 42196 37492
rect 41468 37268 41524 37436
rect 40908 36708 40964 37212
rect 41468 36932 41524 37212
rect 41692 37268 41748 37278
rect 41692 37174 41748 37212
rect 40516 36652 40964 36708
rect 41244 36876 41524 36932
rect 41916 36932 41972 37436
rect 42028 36932 42084 36942
rect 41916 36876 42028 36932
rect 40460 36642 40516 36652
rect 40516 36372 40572 36382
rect 40516 36278 40572 36316
rect 40684 35700 40740 36652
rect 41020 36484 41076 36494
rect 40796 36426 40852 36438
rect 40796 36374 40798 36426
rect 40850 36374 40852 36426
rect 41020 36402 41022 36428
rect 41074 36402 41076 36428
rect 41020 36390 41076 36402
rect 41244 36454 41300 36876
rect 41244 36402 41246 36454
rect 41298 36402 41300 36454
rect 41244 36390 41300 36402
rect 41356 36426 41412 36438
rect 40796 35924 40852 36374
rect 41356 36374 41358 36426
rect 41410 36374 41412 36426
rect 40796 35868 40964 35924
rect 40796 35700 40852 35710
rect 40684 35698 40852 35700
rect 40684 35646 40798 35698
rect 40850 35646 40852 35698
rect 40684 35644 40852 35646
rect 40796 35634 40852 35644
rect 40908 35700 40964 35868
rect 40908 35634 40964 35644
rect 40236 35474 40292 35486
rect 40236 35422 40238 35474
rect 40290 35422 40292 35474
rect 40236 35028 40292 35422
rect 41356 35252 41412 36374
rect 42028 36036 42084 36876
rect 42028 35970 42084 35980
rect 41580 35588 41636 35598
rect 41580 35494 41636 35532
rect 41356 35186 41412 35196
rect 40236 34962 40292 34972
rect 40684 35028 40740 35038
rect 40684 34934 40740 34972
rect 39508 32610 39564 32620
rect 39788 32618 39844 33068
rect 37996 32510 37998 32562
rect 38050 32510 38052 32562
rect 37996 32498 38052 32510
rect 38668 32564 38724 32574
rect 39788 32566 39790 32618
rect 39842 32566 39844 32618
rect 40124 32609 40180 34188
rect 40348 34804 40404 34814
rect 40236 33346 40292 33358
rect 40236 33294 40238 33346
rect 40290 33294 40292 33346
rect 40236 32788 40292 33294
rect 40236 32722 40292 32732
rect 40348 32618 40404 34748
rect 42588 34804 42644 34814
rect 42588 34710 42644 34748
rect 41580 34244 41636 34254
rect 40796 34132 40852 34142
rect 40796 34038 40852 34076
rect 41580 34130 41636 34188
rect 41580 34078 41582 34130
rect 41634 34078 41636 34130
rect 41580 34066 41636 34078
rect 42812 33570 42868 40572
rect 43036 39844 43092 41945
rect 43036 39778 43092 39788
rect 43372 40962 43428 40974
rect 43372 40910 43374 40962
rect 43426 40910 43428 40962
rect 43372 39732 43428 40910
rect 43484 40402 43540 40414
rect 43484 40350 43486 40402
rect 43538 40350 43540 40402
rect 43484 40180 43540 40350
rect 43484 40114 43540 40124
rect 43932 39844 43988 39854
rect 43932 39750 43988 39788
rect 43372 39666 43428 39676
rect 43596 39620 43652 39630
rect 43484 39618 43652 39620
rect 43484 39566 43598 39618
rect 43650 39566 43652 39618
rect 43484 39564 43652 39566
rect 43260 39508 43316 39518
rect 43260 39414 43316 39452
rect 42924 38722 42980 38734
rect 42924 38670 42926 38722
rect 42978 38670 42980 38722
rect 42924 38276 42980 38670
rect 42924 38210 42980 38220
rect 43372 38612 43428 38622
rect 43372 38050 43428 38556
rect 43372 37998 43374 38050
rect 43426 37998 43428 38050
rect 43372 37986 43428 37998
rect 43036 37826 43092 37838
rect 43036 37774 43038 37826
rect 43090 37774 43092 37826
rect 43036 37268 43092 37774
rect 43036 37202 43092 37212
rect 43148 36594 43204 36606
rect 43148 36542 43150 36594
rect 43202 36542 43204 36594
rect 43148 36372 43204 36542
rect 43148 36306 43204 36316
rect 43148 35924 43204 35934
rect 43148 35138 43204 35868
rect 43484 35812 43540 39564
rect 43596 39554 43652 39564
rect 43708 38836 43764 38846
rect 43708 38742 43764 38780
rect 43708 38276 43764 38286
rect 43708 38182 43764 38220
rect 43596 37154 43652 37166
rect 43596 37102 43598 37154
rect 43650 37102 43652 37154
rect 43596 36932 43652 37102
rect 43596 36866 43652 36876
rect 43820 36454 43876 36466
rect 43820 36402 43822 36454
rect 43874 36402 43876 36454
rect 43820 35924 43876 36402
rect 43820 35858 43876 35868
rect 43148 35086 43150 35138
rect 43202 35086 43204 35138
rect 43148 35074 43204 35086
rect 43260 35756 43540 35812
rect 42812 33518 42814 33570
rect 42866 33518 42868 33570
rect 42812 33506 42868 33518
rect 42476 33346 42532 33358
rect 42476 33294 42478 33346
rect 42530 33294 42532 33346
rect 42140 33236 42196 33246
rect 42140 33234 42420 33236
rect 42140 33182 42142 33234
rect 42194 33182 42420 33234
rect 42140 33180 42420 33182
rect 42140 33170 42196 33180
rect 39788 32554 39844 32566
rect 40012 32590 40068 32602
rect 38668 32470 38724 32508
rect 40012 32538 40014 32590
rect 40066 32538 40068 32590
rect 37660 31106 37940 31108
rect 37660 31054 37662 31106
rect 37714 31054 37940 31106
rect 37660 31052 37940 31054
rect 38108 31780 38164 31790
rect 37660 31042 37716 31052
rect 34300 30604 34580 30660
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 36540 30604 36932 30660
rect 33460 30210 34132 30212
rect 33460 30158 33462 30210
rect 33514 30158 34132 30210
rect 33460 30156 34132 30158
rect 33460 30146 33516 30156
rect 32396 29596 33348 29652
rect 32396 29538 32452 29596
rect 32396 29486 32398 29538
rect 32450 29486 32452 29538
rect 32396 29474 32452 29486
rect 32152 29426 32340 29428
rect 32152 29374 32154 29426
rect 32206 29374 32340 29426
rect 32152 29372 32340 29374
rect 36316 29426 36372 29438
rect 36316 29374 36318 29426
rect 36370 29374 36372 29426
rect 32152 29316 32208 29372
rect 31052 28758 31054 28810
rect 31106 28758 31108 28810
rect 31892 28866 32004 28878
rect 31892 28814 31894 28866
rect 31946 28814 32004 28866
rect 31892 28812 32004 28814
rect 32060 29260 32208 29316
rect 36316 29316 36372 29374
rect 31892 28802 31948 28812
rect 31052 28746 31108 28758
rect 30828 28642 30884 28654
rect 30828 28590 30830 28642
rect 30882 28590 30884 28642
rect 30828 28420 30884 28590
rect 31052 28642 31108 28654
rect 31052 28590 31054 28642
rect 31106 28590 31108 28642
rect 31052 28532 31108 28590
rect 31052 28466 31108 28476
rect 31388 28642 31444 28654
rect 31388 28590 31390 28642
rect 31442 28590 31444 28642
rect 30828 28354 30884 28364
rect 31388 28420 31444 28590
rect 31388 28354 31444 28364
rect 31612 28642 31668 28654
rect 32060 28644 32116 29260
rect 36316 29250 36372 29260
rect 36148 29204 36204 29214
rect 35980 29202 36204 29204
rect 35980 29150 36150 29202
rect 36202 29150 36204 29202
rect 35980 29148 36204 29150
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35868 28754 35924 28766
rect 35868 28702 35870 28754
rect 35922 28702 35924 28754
rect 31612 28590 31614 28642
rect 31666 28590 31668 28642
rect 31612 28532 31668 28590
rect 31164 28084 31220 28094
rect 31164 27990 31220 28028
rect 31612 27188 31668 28476
rect 31612 27122 31668 27132
rect 31948 28588 32116 28644
rect 34524 28644 34580 28654
rect 35420 28644 35476 28654
rect 30940 26290 30996 26302
rect 30940 26238 30942 26290
rect 30994 26238 30996 26290
rect 30940 26180 30996 26238
rect 30940 26114 30996 26124
rect 30604 26068 30660 26078
rect 30604 25974 30660 26012
rect 30716 25620 30772 25630
rect 30716 25526 30772 25564
rect 31948 24836 32004 28588
rect 33740 28418 33796 28430
rect 33740 28366 33742 28418
rect 33794 28366 33796 28418
rect 32060 28084 32116 28094
rect 32060 26908 32116 28028
rect 33740 27972 33796 28366
rect 33292 27916 33796 27972
rect 33964 28028 34468 28084
rect 33964 28026 34020 28028
rect 33964 27974 33966 28026
rect 34018 27974 34020 28026
rect 33964 27962 34020 27974
rect 32508 27885 32564 27897
rect 32508 27833 32510 27885
rect 32562 27833 32564 27885
rect 32508 27300 32564 27833
rect 32508 27234 32564 27244
rect 32172 27188 32228 27198
rect 32172 27094 32228 27132
rect 32956 27074 33012 27086
rect 32956 27022 32958 27074
rect 33010 27022 33012 27074
rect 32956 26908 33012 27022
rect 32060 26852 32228 26908
rect 32172 26334 32228 26852
rect 32172 26282 32174 26334
rect 32226 26282 32228 26334
rect 32172 26270 32228 26282
rect 32396 26852 33012 26908
rect 33180 27076 33236 27086
rect 32060 26178 32116 26190
rect 32060 26126 32062 26178
rect 32114 26126 32116 26178
rect 32060 25620 32116 26126
rect 32060 25554 32116 25564
rect 31948 24770 32004 24780
rect 31500 24498 31556 24510
rect 31500 24446 31502 24498
rect 31554 24446 31556 24498
rect 30492 24220 31220 24276
rect 30156 24052 30212 24062
rect 30156 23958 30212 23996
rect 31052 24052 31108 24062
rect 29932 23268 29988 23278
rect 29932 23154 29988 23212
rect 31052 23266 31108 23996
rect 31052 23214 31054 23266
rect 31106 23214 31108 23266
rect 31052 23202 31108 23214
rect 29932 23102 29934 23154
rect 29986 23102 29988 23154
rect 29932 23090 29988 23102
rect 30808 23156 30864 23166
rect 30808 23062 30864 23100
rect 30808 22596 30864 22606
rect 29932 22372 29988 22382
rect 29932 22278 29988 22316
rect 30604 22372 30660 22382
rect 29708 22092 29988 22148
rect 29596 21970 29652 21980
rect 29204 21698 29428 21700
rect 29204 21646 29206 21698
rect 29258 21646 29428 21698
rect 29204 21644 29428 21646
rect 29764 21812 29820 21822
rect 29204 21634 29260 21644
rect 29764 21642 29820 21756
rect 29484 21586 29540 21598
rect 29484 21534 29486 21586
rect 29538 21534 29540 21586
rect 29372 21476 29428 21486
rect 29372 21026 29428 21420
rect 29372 20974 29374 21026
rect 29426 20974 29428 21026
rect 29372 20962 29428 20974
rect 29036 19964 29428 20020
rect 28812 19394 28868 19404
rect 29148 19236 29204 19246
rect 28700 19234 29204 19236
rect 28700 19182 29150 19234
rect 29202 19182 29204 19234
rect 28700 19180 29204 19182
rect 28476 18788 28532 19180
rect 28644 19010 28700 19022
rect 28644 18958 28646 19010
rect 28698 18958 28700 19010
rect 28644 18910 28700 18958
rect 28644 18900 28756 18910
rect 28644 18844 28700 18900
rect 28756 18844 29092 18900
rect 28700 18806 28756 18844
rect 28476 18732 28644 18788
rect 28252 18498 28308 18508
rect 28476 18450 28532 18462
rect 28476 18398 28478 18450
rect 28530 18398 28532 18450
rect 28252 18340 28308 18350
rect 28252 18246 28308 18284
rect 28140 17892 28196 18172
rect 28364 17892 28420 17902
rect 28140 17890 28420 17892
rect 28140 17838 28366 17890
rect 28418 17838 28420 17890
rect 28140 17836 28420 17838
rect 28364 17826 28420 17836
rect 28028 16930 28084 16940
rect 28476 17108 28532 18398
rect 28588 17444 28644 18732
rect 28812 18452 28868 18462
rect 28812 18358 28868 18396
rect 28700 18340 28756 18350
rect 28700 17666 28756 18284
rect 28700 17614 28702 17666
rect 28754 17614 28756 17666
rect 28700 17602 28756 17614
rect 28588 17388 28980 17444
rect 28476 16882 28532 17052
rect 28476 16830 28478 16882
rect 28530 16830 28532 16882
rect 28476 16818 28532 16830
rect 28588 17220 28644 17230
rect 27468 16716 27636 16772
rect 27692 16772 27748 16782
rect 27468 16660 27524 16716
rect 27468 16594 27524 16604
rect 27580 16548 27636 16558
rect 27468 16212 27524 16222
rect 27244 16156 27468 16212
rect 27132 16046 27134 16098
rect 27186 16046 27188 16098
rect 27132 16034 27188 16046
rect 27468 16098 27524 16156
rect 27468 16046 27470 16098
rect 27522 16046 27524 16098
rect 27468 16034 27524 16046
rect 26124 15876 26180 15886
rect 27580 15876 27636 16492
rect 27692 16098 27748 16716
rect 27804 16770 27860 16782
rect 27804 16718 27806 16770
rect 27858 16718 27860 16770
rect 27804 16548 27860 16718
rect 27804 16482 27860 16492
rect 28588 16334 28644 17164
rect 28532 16322 28644 16334
rect 28532 16270 28534 16322
rect 28586 16270 28644 16322
rect 28532 16268 28644 16270
rect 28532 16258 28588 16268
rect 27692 16046 27694 16098
rect 27746 16046 27748 16098
rect 27692 16034 27748 16046
rect 27804 16100 27860 16110
rect 26124 15316 26180 15820
rect 27468 15820 27636 15876
rect 27468 15428 27524 15820
rect 26124 15222 26180 15260
rect 26796 15314 26852 15326
rect 26796 15262 26798 15314
rect 26850 15262 26852 15314
rect 26012 15138 26068 15148
rect 26460 15202 26516 15214
rect 26460 15150 26462 15202
rect 26514 15150 26516 15202
rect 26460 14532 26516 15150
rect 26460 14466 26516 14476
rect 26516 14308 26572 14318
rect 26796 14308 26852 15262
rect 27244 14532 27300 14542
rect 27244 14438 27300 14476
rect 27468 14530 27524 15372
rect 27580 15204 27636 15242
rect 27580 15138 27636 15148
rect 27804 14868 27860 16044
rect 28364 16100 28420 16110
rect 28364 16006 28420 16044
rect 28028 15876 28084 15886
rect 28028 15782 28084 15820
rect 28700 15316 28756 15326
rect 27468 14478 27470 14530
rect 27522 14478 27524 14530
rect 27636 14812 27860 14868
rect 28140 14980 28196 14990
rect 28700 14980 28756 15260
rect 27636 14586 27692 14812
rect 27636 14534 27638 14586
rect 27690 14534 27692 14586
rect 27636 14522 27692 14534
rect 28140 14530 28196 14924
rect 28382 14924 28756 14980
rect 28382 14754 28438 14924
rect 28382 14702 28384 14754
rect 28436 14702 28438 14754
rect 28382 14690 28438 14702
rect 28924 14644 28980 17388
rect 29036 15540 29092 18844
rect 29148 18465 29204 19180
rect 29148 18413 29150 18465
rect 29202 18413 29204 18465
rect 29148 18116 29204 18413
rect 29260 18676 29316 18686
rect 29260 18338 29316 18620
rect 29260 18286 29262 18338
rect 29314 18286 29316 18338
rect 29260 18274 29316 18286
rect 29372 18116 29428 19964
rect 29484 19460 29540 21534
rect 29596 21586 29652 21598
rect 29596 21534 29598 21586
rect 29650 21534 29652 21586
rect 29764 21590 29766 21642
rect 29818 21590 29820 21642
rect 29764 21578 29820 21590
rect 29932 21586 29988 22092
rect 29596 20020 29652 21534
rect 29932 21534 29934 21586
rect 29986 21534 29988 21586
rect 29932 21522 29988 21534
rect 30044 22036 30100 22046
rect 30044 21028 30100 21980
rect 30380 21588 30436 21598
rect 30380 21494 30436 21532
rect 30604 21418 30660 22316
rect 30808 22370 30864 22540
rect 30808 22318 30810 22370
rect 30862 22318 30864 22370
rect 30808 22306 30864 22318
rect 31052 22260 31108 22270
rect 30604 21366 30606 21418
rect 30658 21366 30660 21418
rect 30940 22258 31108 22260
rect 30940 22206 31054 22258
rect 31106 22206 31108 22258
rect 30940 22204 31108 22206
rect 30604 21354 30660 21366
rect 30716 21364 30772 21374
rect 29820 20972 30100 21028
rect 29708 20804 29764 20814
rect 29708 20710 29764 20748
rect 29596 19954 29652 19964
rect 29820 19796 29876 20972
rect 30716 20970 30772 21308
rect 30716 20918 30718 20970
rect 30770 20918 30772 20970
rect 30716 20906 30772 20918
rect 29932 20802 29988 20814
rect 29932 20750 29934 20802
rect 29986 20750 29988 20802
rect 29932 20356 29988 20750
rect 30380 20804 30436 20814
rect 29932 20300 30212 20356
rect 29932 20132 29988 20142
rect 29932 20038 29988 20076
rect 29820 19730 29876 19740
rect 30156 19908 30212 20300
rect 29484 19404 30100 19460
rect 29484 19402 29540 19404
rect 29484 19350 29486 19402
rect 29538 19350 29540 19402
rect 29484 19338 29540 19350
rect 29484 19234 29540 19246
rect 29484 19182 29486 19234
rect 29538 19182 29540 19234
rect 29484 18340 29540 19182
rect 30044 18450 30100 19404
rect 30156 19236 30212 19852
rect 30156 19170 30212 19180
rect 30268 20018 30324 20030
rect 30268 19966 30270 20018
rect 30322 19966 30324 20018
rect 30268 18452 30324 19966
rect 30044 18398 30046 18450
rect 30098 18398 30100 18450
rect 30044 18386 30100 18398
rect 30156 18450 30324 18452
rect 30156 18398 30270 18450
rect 30322 18398 30324 18450
rect 30156 18396 30324 18398
rect 29484 18274 29540 18284
rect 30156 18228 30212 18396
rect 30268 18386 30324 18396
rect 29876 18172 30212 18228
rect 29372 18060 29764 18116
rect 29148 18050 29204 18060
rect 29372 17666 29428 17678
rect 29372 17614 29374 17666
rect 29426 17614 29428 17666
rect 29372 17220 29428 17614
rect 29372 17154 29428 17164
rect 29596 17668 29652 17678
rect 29484 16884 29540 16894
rect 29372 16882 29540 16884
rect 29372 16830 29486 16882
rect 29538 16830 29540 16882
rect 29372 16828 29540 16830
rect 29148 16100 29204 16110
rect 29372 16100 29428 16828
rect 29484 16818 29540 16828
rect 29596 16660 29652 17612
rect 29708 16772 29764 18060
rect 29876 17890 29932 18172
rect 30380 17892 30436 20748
rect 30492 20802 30548 20814
rect 30492 20750 30494 20802
rect 30546 20750 30548 20802
rect 30492 20132 30548 20750
rect 30492 20066 30548 20076
rect 30716 20020 30772 20030
rect 30716 18564 30772 19964
rect 29876 17838 29878 17890
rect 29930 17838 29932 17890
rect 29876 17826 29932 17838
rect 30268 17836 30436 17892
rect 30548 18226 30604 18238
rect 30548 18174 30550 18226
rect 30602 18174 30604 18226
rect 30156 17668 30212 17678
rect 30044 17666 30212 17668
rect 30044 17614 30158 17666
rect 30210 17614 30212 17666
rect 30044 17612 30212 17614
rect 30044 17108 30100 17612
rect 30156 17602 30212 17612
rect 30268 17444 30324 17836
rect 30380 17668 30436 17678
rect 30380 17574 30436 17612
rect 30548 17668 30604 18174
rect 30716 17902 30772 18508
rect 30660 17890 30772 17902
rect 30660 17838 30662 17890
rect 30714 17838 30772 17890
rect 30660 17836 30772 17838
rect 30828 18676 30884 18686
rect 30660 17826 30716 17836
rect 30548 17602 30604 17612
rect 30268 17388 30436 17444
rect 29932 17052 30100 17108
rect 30156 17108 30212 17118
rect 29820 16996 29876 17006
rect 29820 16938 29876 16940
rect 29820 16886 29822 16938
rect 29874 16886 29876 16938
rect 29820 16874 29876 16886
rect 29708 16706 29764 16716
rect 29932 16770 29988 17052
rect 30156 16882 30212 17052
rect 30156 16830 30158 16882
rect 30210 16830 30212 16882
rect 30156 16818 30212 16830
rect 29932 16718 29934 16770
rect 29986 16718 29988 16770
rect 29204 16044 29428 16100
rect 29148 16006 29204 16044
rect 29036 15474 29092 15484
rect 29372 15428 29428 16044
rect 29484 16604 29652 16660
rect 29932 16660 29988 16718
rect 29932 16604 30100 16660
rect 29484 16054 29540 16604
rect 29932 16324 29988 16334
rect 29596 16212 29652 16222
rect 29596 16118 29652 16156
rect 29932 16210 29988 16268
rect 29932 16158 29934 16210
rect 29986 16158 29988 16210
rect 29932 16146 29988 16158
rect 29484 16002 29486 16054
rect 29538 16002 29540 16054
rect 30044 16083 30100 16604
rect 30044 16031 30046 16083
rect 30098 16031 30100 16083
rect 30044 16019 30100 16031
rect 30268 16098 30324 16110
rect 30268 16046 30270 16098
rect 30322 16046 30324 16098
rect 29484 15988 29540 16002
rect 29484 15922 29540 15932
rect 29484 15428 29540 15438
rect 29372 15426 29540 15428
rect 29372 15374 29486 15426
rect 29538 15374 29540 15426
rect 29372 15372 29540 15374
rect 29484 15362 29540 15372
rect 29820 15428 29876 15438
rect 28924 14578 28980 14588
rect 29484 14644 29540 14654
rect 27468 14466 27524 14478
rect 28140 14478 28142 14530
rect 28194 14478 28196 14530
rect 26908 14308 26964 14318
rect 26796 14306 26964 14308
rect 26796 14254 26910 14306
rect 26962 14254 26964 14306
rect 26796 14252 26964 14254
rect 26516 14214 26572 14252
rect 26908 13748 26964 14252
rect 28140 14308 28196 14478
rect 28140 14242 28196 14252
rect 28588 14532 28644 14542
rect 26908 13682 26964 13692
rect 27692 13748 27748 13758
rect 27692 13654 27748 13692
rect 28476 13634 28532 13646
rect 28476 13582 28478 13634
rect 28530 13582 28532 13634
rect 28476 13188 28532 13582
rect 28476 13122 28532 13132
rect 27356 12962 27412 12974
rect 26852 12906 26908 12918
rect 26684 12852 26740 12862
rect 26572 12850 26740 12852
rect 26572 12798 26686 12850
rect 26738 12798 26740 12850
rect 26572 12796 26740 12798
rect 25564 9158 25566 9210
rect 25618 9158 25620 9210
rect 25564 9146 25620 9158
rect 25676 12348 25956 12404
rect 26404 12738 26460 12750
rect 26404 12686 26406 12738
rect 26458 12686 26460 12738
rect 25340 9042 25508 9044
rect 25340 8990 25342 9042
rect 25394 8990 25508 9042
rect 25340 8988 25508 8990
rect 25564 9069 25620 9081
rect 25564 9017 25566 9069
rect 25618 9017 25620 9069
rect 25340 8978 25396 8988
rect 25564 8596 25620 9017
rect 25564 8530 25620 8540
rect 25228 8484 25284 8494
rect 25228 8370 25284 8428
rect 25676 8372 25732 12348
rect 25900 12180 25956 12190
rect 26404 12180 26460 12686
rect 26572 12292 26628 12796
rect 26684 12786 26740 12796
rect 26852 12854 26854 12906
rect 26906 12854 26908 12906
rect 26852 12404 26908 12854
rect 27356 12910 27358 12962
rect 27410 12910 27412 12962
rect 27356 12852 27412 12910
rect 27356 12786 27412 12796
rect 27598 12852 27654 12862
rect 27598 12850 27860 12852
rect 27598 12798 27600 12850
rect 27652 12798 27860 12850
rect 27598 12796 27860 12798
rect 27598 12786 27654 12796
rect 26852 12348 26964 12404
rect 26572 12198 26628 12236
rect 25900 12178 26460 12180
rect 25900 12126 25902 12178
rect 25954 12126 26460 12178
rect 25900 12124 26460 12126
rect 25900 10052 25956 12124
rect 26740 12122 26796 12134
rect 26740 12070 26742 12122
rect 26794 12070 26796 12122
rect 26142 11956 26198 11966
rect 26142 11862 26198 11900
rect 26012 11732 26068 11742
rect 26012 11506 26068 11676
rect 26740 11620 26796 12070
rect 26908 11732 26964 12348
rect 27244 12178 27300 12190
rect 27244 12126 27246 12178
rect 27298 12126 27300 12178
rect 27244 12068 27300 12126
rect 27804 12178 27860 12796
rect 27804 12126 27806 12178
rect 27858 12126 27860 12178
rect 27804 12114 27860 12126
rect 28252 12740 28308 12750
rect 27244 12002 27300 12012
rect 27486 11956 27542 11966
rect 28140 11956 28196 11966
rect 27486 11954 27860 11956
rect 27486 11902 27488 11954
rect 27540 11902 27860 11954
rect 27486 11900 27860 11902
rect 27486 11890 27542 11900
rect 27020 11732 27076 11742
rect 26908 11676 27020 11732
rect 27020 11666 27076 11676
rect 26740 11554 26796 11564
rect 26012 11454 26014 11506
rect 26066 11454 26068 11506
rect 26012 10276 26068 11454
rect 27804 11284 27860 11900
rect 27916 11954 28196 11956
rect 27916 11902 28142 11954
rect 28194 11902 28196 11954
rect 27916 11900 28196 11902
rect 27916 11506 27972 11900
rect 28140 11890 28196 11900
rect 27916 11454 27918 11506
rect 27970 11454 27972 11506
rect 27916 11442 27972 11454
rect 27804 11228 28196 11284
rect 28028 10610 28084 10622
rect 28028 10558 28030 10610
rect 28082 10558 28084 10610
rect 27244 10500 27300 10510
rect 27244 10406 27300 10444
rect 28028 10388 28084 10558
rect 28140 10610 28196 11228
rect 28140 10558 28142 10610
rect 28194 10558 28196 10610
rect 28140 10546 28196 10558
rect 28252 10388 28308 12684
rect 28588 11396 28644 14476
rect 29484 14530 29540 14588
rect 29484 14478 29486 14530
rect 29538 14478 29540 14530
rect 29484 14466 29540 14478
rect 29242 14420 29298 14430
rect 28700 14418 29298 14420
rect 28700 14366 29244 14418
rect 29296 14366 29298 14418
rect 28700 14364 29298 14366
rect 28700 13412 28756 14364
rect 29242 14354 29298 14364
rect 29820 14362 29876 15372
rect 30156 15316 30212 15326
rect 30268 15316 30324 16046
rect 30156 15314 30324 15316
rect 30156 15262 30158 15314
rect 30210 15262 30324 15314
rect 30156 15260 30324 15262
rect 30156 15148 30212 15260
rect 29820 14310 29822 14362
rect 29874 14310 29876 14362
rect 29820 14298 29876 14310
rect 29988 15092 30212 15148
rect 30380 15148 30436 17388
rect 30492 16884 30548 16894
rect 30492 16790 30548 16828
rect 30828 16884 30884 18620
rect 30828 16818 30884 16828
rect 30828 16714 30884 16726
rect 30828 16662 30830 16714
rect 30882 16662 30884 16714
rect 30604 15988 30660 15998
rect 30492 15428 30548 15438
rect 30492 15370 30548 15372
rect 30492 15318 30494 15370
rect 30546 15318 30548 15370
rect 30492 15306 30548 15318
rect 30604 15202 30660 15932
rect 30604 15150 30606 15202
rect 30658 15150 30660 15202
rect 30380 15092 30548 15148
rect 30604 15138 30660 15150
rect 30716 15314 30772 15326
rect 30716 15262 30718 15314
rect 30770 15262 30772 15314
rect 29988 14474 30044 15092
rect 29988 14422 29990 14474
rect 30042 14422 30044 14474
rect 29988 13860 30044 14422
rect 30380 13860 30436 13870
rect 29988 13858 30436 13860
rect 29988 13806 30382 13858
rect 30434 13806 30436 13858
rect 29988 13804 30436 13806
rect 30380 13794 30436 13804
rect 30492 13636 30548 15092
rect 30604 14980 30660 14990
rect 30604 14588 30660 14924
rect 30716 14756 30772 15262
rect 30828 15092 30884 16662
rect 30940 15148 30996 22204
rect 31052 22194 31108 22204
rect 31164 22036 31220 24220
rect 31388 23492 31444 23502
rect 31388 23154 31444 23436
rect 31388 23102 31390 23154
rect 31442 23102 31444 23154
rect 31388 23090 31444 23102
rect 31500 23156 31556 24446
rect 32396 24388 32452 26852
rect 33180 26526 33236 27020
rect 33292 27059 33348 27916
rect 33740 27902 33796 27916
rect 33740 27850 33742 27902
rect 33794 27850 33796 27902
rect 33740 27838 33796 27850
rect 34076 27858 34132 27870
rect 34076 27806 34078 27858
rect 34130 27806 34132 27858
rect 33292 27007 33294 27059
rect 33346 27007 33348 27059
rect 33292 26995 33348 27007
rect 33404 27186 33460 27198
rect 33404 27134 33406 27186
rect 33458 27134 33460 27186
rect 33180 26514 33292 26526
rect 33180 26462 33238 26514
rect 33290 26462 33292 26514
rect 33180 26460 33292 26462
rect 33236 26450 33292 26460
rect 32508 26292 32564 26302
rect 33068 26292 33124 26302
rect 32508 26290 33068 26292
rect 32508 26238 32510 26290
rect 32562 26238 33068 26290
rect 32508 26236 33068 26238
rect 32508 26226 32564 26236
rect 32620 25618 32676 26236
rect 33068 26198 33124 26236
rect 33404 25732 33460 27134
rect 34076 27188 34132 27806
rect 34076 27122 34132 27132
rect 34412 27186 34468 28028
rect 34412 27134 34414 27186
rect 34466 27134 34468 27186
rect 34412 27122 34468 27134
rect 34524 27970 34580 28588
rect 34524 27918 34526 27970
rect 34578 27918 34580 27970
rect 33628 27076 33684 27086
rect 33628 26982 33684 27020
rect 34524 26908 34580 27918
rect 34748 28614 34804 28626
rect 34748 28562 34750 28614
rect 34802 28562 34804 28614
rect 34748 27636 34804 28562
rect 35420 28550 35476 28588
rect 35756 28598 35812 28610
rect 35756 28546 35758 28598
rect 35810 28546 35812 28598
rect 35756 28084 35812 28546
rect 35868 28196 35924 28702
rect 35980 28532 36036 29148
rect 36148 29138 36204 29148
rect 35980 28466 36036 28476
rect 36428 28642 36484 28654
rect 36428 28590 36430 28642
rect 36482 28590 36484 28642
rect 36260 28420 36316 28430
rect 36260 28326 36316 28364
rect 36428 28308 36484 28590
rect 36428 28242 36484 28252
rect 35868 28140 36260 28196
rect 35756 28018 35812 28028
rect 36204 27860 36260 28140
rect 36428 27860 36484 27870
rect 36204 27858 36484 27860
rect 36204 27806 36430 27858
rect 36482 27806 36484 27858
rect 36204 27804 36484 27806
rect 36428 27794 36484 27804
rect 34300 26852 34580 26908
rect 34636 27580 34804 27636
rect 33628 26292 33684 26302
rect 33628 26198 33684 26236
rect 33404 25676 33684 25732
rect 32620 25566 32622 25618
rect 32674 25566 32676 25618
rect 32620 25554 32676 25566
rect 33292 25478 33348 25490
rect 33292 25426 33294 25478
rect 33346 25426 33348 25478
rect 32508 25396 32564 25406
rect 32508 24749 32564 25340
rect 32508 24697 32510 24749
rect 32562 24697 32564 24749
rect 32956 24724 33012 24734
rect 32508 24685 32564 24697
rect 32732 24722 33012 24724
rect 32732 24670 32958 24722
rect 33010 24670 33012 24722
rect 32732 24668 33012 24670
rect 32396 24332 32564 24388
rect 32396 24164 32452 24174
rect 31500 23090 31556 23100
rect 31836 23938 31892 23950
rect 31836 23886 31838 23938
rect 31890 23886 31892 23938
rect 31120 21980 31220 22036
rect 31500 22932 31556 22942
rect 31120 21624 31176 21980
rect 31120 21572 31122 21624
rect 31174 21572 31176 21624
rect 31120 21140 31176 21572
rect 31500 21486 31556 22876
rect 31724 22930 31780 22942
rect 31724 22878 31726 22930
rect 31778 22878 31780 22930
rect 31612 22146 31668 22158
rect 31612 22094 31614 22146
rect 31666 22094 31668 22146
rect 31612 21812 31668 22094
rect 31612 21746 31668 21756
rect 31500 21476 31612 21486
rect 31500 21474 31668 21476
rect 31500 21422 31558 21474
rect 31610 21422 31668 21474
rect 31500 21420 31668 21422
rect 31556 21410 31668 21420
rect 31120 21084 31220 21140
rect 31164 20580 31220 21084
rect 31332 20580 31388 20590
rect 31164 20524 31332 20580
rect 31332 20486 31388 20524
rect 31388 20018 31444 20030
rect 31388 19966 31390 20018
rect 31442 19966 31444 20018
rect 31388 19908 31444 19966
rect 31388 19842 31444 19852
rect 31388 18564 31444 18574
rect 31388 18450 31444 18508
rect 31388 18398 31390 18450
rect 31442 18398 31444 18450
rect 31388 17666 31444 18398
rect 31388 17614 31390 17666
rect 31442 17614 31444 17666
rect 31388 17602 31444 17614
rect 31612 17332 31668 21410
rect 31724 20804 31780 22878
rect 31836 22372 31892 23886
rect 32172 23714 32228 23726
rect 32172 23662 32174 23714
rect 32226 23662 32228 23714
rect 32172 23268 32228 23662
rect 32396 23378 32452 24108
rect 32396 23326 32398 23378
rect 32450 23326 32452 23378
rect 32396 23314 32452 23326
rect 32172 23202 32228 23212
rect 32060 23156 32116 23166
rect 32060 23062 32116 23100
rect 32508 23156 32564 24332
rect 32732 23380 32788 24668
rect 32956 24658 33012 24668
rect 33292 24052 33348 25426
rect 33628 24724 33684 25676
rect 34300 24948 34356 26852
rect 34504 26292 34560 26302
rect 34504 26290 34580 26292
rect 34504 26238 34506 26290
rect 34558 26238 34580 26290
rect 34504 26226 34580 26238
rect 33852 24892 34356 24948
rect 34524 24948 34580 26226
rect 34636 25732 34692 27580
rect 35868 27524 35924 27534
rect 36540 27524 36596 30604
rect 37772 30210 37828 30222
rect 37772 30158 37774 30210
rect 37826 30158 37828 30210
rect 37604 29988 37660 29998
rect 37772 29988 37828 30158
rect 38108 30210 38164 31724
rect 39564 31780 39620 31790
rect 39564 31686 39620 31724
rect 40012 30772 40068 32538
rect 40124 32597 40236 32609
rect 40124 32545 40182 32597
rect 40234 32545 40236 32597
rect 40348 32566 40350 32618
rect 40402 32566 40404 32618
rect 40348 32554 40404 32566
rect 40124 32535 40236 32545
rect 40180 32533 40236 32535
rect 42252 31892 42308 31902
rect 42252 31798 42308 31836
rect 40012 30706 40068 30716
rect 40348 31778 40404 31790
rect 40348 31726 40350 31778
rect 40402 31726 40404 31778
rect 40348 30324 40404 31726
rect 41468 30996 41524 31006
rect 41468 30994 41748 30996
rect 41468 30942 41470 30994
rect 41522 30942 41748 30994
rect 41468 30940 41748 30942
rect 41468 30930 41524 30940
rect 41300 30772 41356 30782
rect 41300 30770 41636 30772
rect 41300 30718 41302 30770
rect 41354 30718 41636 30770
rect 41300 30716 41636 30718
rect 41300 30706 41356 30716
rect 40460 30324 40516 30334
rect 40348 30268 40460 30324
rect 40460 30230 40516 30268
rect 38108 30158 38110 30210
rect 38162 30158 38164 30210
rect 38108 30146 38164 30158
rect 38556 30210 38612 30222
rect 38556 30158 38558 30210
rect 38610 30158 38612 30210
rect 37604 29986 37828 29988
rect 37604 29934 37606 29986
rect 37658 29934 37828 29986
rect 37604 29932 37828 29934
rect 37604 29922 37660 29932
rect 37772 29876 37828 29932
rect 37772 29820 38164 29876
rect 37436 29441 37492 29453
rect 36876 29428 36932 29438
rect 36876 29334 36932 29372
rect 37212 29426 37268 29438
rect 37212 29374 37214 29426
rect 37266 29374 37268 29426
rect 37212 29316 37268 29374
rect 37212 29250 37268 29260
rect 37324 29428 37380 29438
rect 36708 29202 36764 29214
rect 36708 29150 36710 29202
rect 36762 29150 36764 29202
rect 36708 28644 36764 29150
rect 36708 28578 36764 28588
rect 36988 28754 37044 28766
rect 36988 28702 36990 28754
rect 37042 28702 37044 28754
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35084 26852 35140 26862
rect 35084 26290 35140 26796
rect 35084 26238 35086 26290
rect 35138 26238 35140 26290
rect 35084 26226 35140 26238
rect 35868 26290 35924 27468
rect 35868 26238 35870 26290
rect 35922 26238 35924 26290
rect 35868 26226 35924 26238
rect 35980 27468 36596 27524
rect 36652 28420 36708 28430
rect 34748 26068 34804 26078
rect 34748 25974 34804 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34636 25666 34692 25676
rect 34972 25396 35028 25406
rect 34972 25302 35028 25340
rect 34524 24892 34916 24948
rect 33740 24724 33796 24734
rect 33628 24722 33796 24724
rect 33628 24670 33742 24722
rect 33794 24670 33796 24722
rect 33628 24668 33796 24670
rect 33740 24658 33796 24668
rect 33292 23986 33348 23996
rect 33628 24052 33684 24062
rect 33628 23958 33684 23996
rect 32844 23940 32900 23950
rect 32844 23938 33180 23940
rect 32844 23886 32846 23938
rect 32898 23886 33180 23938
rect 32844 23884 33180 23886
rect 32844 23874 32900 23884
rect 32732 23314 32788 23324
rect 33124 23378 33180 23884
rect 33124 23326 33126 23378
rect 33178 23326 33180 23378
rect 33124 23314 33180 23326
rect 33572 23380 33628 23390
rect 33572 23286 33628 23324
rect 32508 23090 32564 23100
rect 33292 23156 33348 23166
rect 33292 23062 33348 23100
rect 33740 23156 33796 23166
rect 33852 23156 33908 24892
rect 34860 23380 34916 24892
rect 35644 24610 35700 24622
rect 35644 24558 35646 24610
rect 35698 24558 35700 24610
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35532 23940 35588 23950
rect 35532 23846 35588 23884
rect 35644 23716 35700 24558
rect 35980 24276 36036 27468
rect 36316 27188 36372 27198
rect 36316 27094 36372 27132
rect 36652 27076 36708 28364
rect 36652 27010 36708 27020
rect 36876 28308 36932 28318
rect 36876 27188 36932 28252
rect 36988 27524 37044 28702
rect 37324 28642 37380 29372
rect 36988 27458 37044 27468
rect 37100 28598 37156 28610
rect 37100 28546 37102 28598
rect 37154 28546 37156 28598
rect 36092 26964 36148 26974
rect 36092 25732 36148 26908
rect 36876 26740 36932 27132
rect 36988 27046 37044 27058
rect 36988 26994 36990 27046
rect 37042 26994 37044 27046
rect 36988 26964 37044 26994
rect 36988 26898 37044 26908
rect 36876 26684 37044 26740
rect 36204 25732 36260 25742
rect 36092 25730 36260 25732
rect 36092 25678 36206 25730
rect 36258 25678 36260 25730
rect 36092 25676 36260 25678
rect 36204 25666 36260 25676
rect 36988 25620 37044 26684
rect 36876 25564 37044 25620
rect 37100 25620 37156 28546
rect 37324 28590 37326 28642
rect 37378 28590 37380 28642
rect 37212 28532 37268 28542
rect 37212 27858 37268 28476
rect 37212 27806 37214 27858
rect 37266 27806 37268 27858
rect 37212 27794 37268 27806
rect 37324 26404 37380 28590
rect 37436 29389 37438 29441
rect 37490 29389 37492 29441
rect 37436 28532 37492 29389
rect 37436 28466 37492 28476
rect 37548 29314 37604 29326
rect 37548 29262 37550 29314
rect 37602 29262 37604 29314
rect 37548 27860 37604 29262
rect 37548 27794 37604 27804
rect 37772 29316 37828 29326
rect 37772 27746 37828 29260
rect 37884 28644 37940 28654
rect 37884 28550 37940 28588
rect 37772 27694 37774 27746
rect 37826 27694 37828 27746
rect 37772 26908 37828 27694
rect 37996 27300 38052 27310
rect 37996 27206 38052 27244
rect 37324 26338 37380 26348
rect 37548 26852 37828 26908
rect 38108 26908 38164 29820
rect 38556 28532 38612 30158
rect 39676 30210 39732 30222
rect 39676 30158 39678 30210
rect 39730 30158 39732 30210
rect 38892 29986 38948 29998
rect 38892 29934 38894 29986
rect 38946 29934 38948 29986
rect 38668 28756 38724 28766
rect 38668 28662 38724 28700
rect 38556 27076 38612 28476
rect 38892 28084 38948 29934
rect 39508 29988 39564 29998
rect 39676 29988 39732 30158
rect 39508 29986 39732 29988
rect 39508 29934 39510 29986
rect 39562 29934 39732 29986
rect 39508 29932 39732 29934
rect 39508 29922 39564 29932
rect 39676 29876 39732 29932
rect 39676 29820 39956 29876
rect 39340 29316 39396 29326
rect 39340 29222 39396 29260
rect 38892 28018 38948 28028
rect 39676 27860 39732 27870
rect 39676 27766 39732 27804
rect 38556 27010 38612 27020
rect 39676 27076 39732 27086
rect 39676 26982 39732 27020
rect 38108 26852 38276 26908
rect 36540 25508 36596 25518
rect 36540 25414 36596 25452
rect 36316 25284 36372 25294
rect 36204 25228 36316 25284
rect 33740 23154 33908 23156
rect 33740 23102 33742 23154
rect 33794 23102 33908 23154
rect 33740 23100 33908 23102
rect 33740 23090 33796 23100
rect 31836 22306 31892 22316
rect 31948 22370 32004 22382
rect 31948 22318 31950 22370
rect 32002 22318 32004 22370
rect 31948 22148 32004 22318
rect 33852 22372 33908 23100
rect 34524 23324 34916 23380
rect 35532 23660 35700 23716
rect 35868 24220 36036 24276
rect 36092 24749 36148 24761
rect 36092 24697 36094 24749
rect 36146 24697 36148 24749
rect 34188 22372 34244 22382
rect 33852 22306 33908 22316
rect 33964 22370 34244 22372
rect 33964 22318 34190 22370
rect 34242 22318 34244 22370
rect 33964 22316 34244 22318
rect 31948 22092 32228 22148
rect 32004 21812 32060 21822
rect 32004 21810 32116 21812
rect 32004 21758 32006 21810
rect 32058 21758 32116 21810
rect 32004 21746 32116 21758
rect 32060 21700 32116 21746
rect 32060 21364 32116 21644
rect 32172 21588 32228 22092
rect 32340 22146 32396 22158
rect 32340 22094 32342 22146
rect 32394 22094 32396 22146
rect 32340 22036 32396 22094
rect 32340 21970 32396 21980
rect 33292 22148 33348 22158
rect 32172 21522 32228 21532
rect 32956 21812 33012 21822
rect 32956 21586 33012 21756
rect 32956 21534 32958 21586
rect 33010 21534 33012 21586
rect 32060 21308 32228 21364
rect 32060 21140 32116 21150
rect 32060 21026 32116 21084
rect 32060 20974 32062 21026
rect 32114 20974 32116 21026
rect 32060 20962 32116 20974
rect 31724 20738 31780 20748
rect 31724 19794 31780 19806
rect 31724 19742 31726 19794
rect 31778 19742 31780 19794
rect 31724 18564 31780 19742
rect 32172 19796 32228 21308
rect 32396 20802 32452 20814
rect 32396 20750 32398 20802
rect 32450 20750 32452 20802
rect 32396 20244 32452 20750
rect 32508 20804 32564 20814
rect 32508 20710 32564 20748
rect 32956 20804 33012 21534
rect 33292 20914 33348 22092
rect 33852 22148 33908 22158
rect 33852 22054 33908 22092
rect 33740 21474 33796 21486
rect 33740 21422 33742 21474
rect 33794 21422 33796 21474
rect 33740 21140 33796 21422
rect 33964 21140 34020 22316
rect 34188 22306 34244 22316
rect 34524 21812 34580 23324
rect 34860 23156 34916 23194
rect 34860 23090 34916 23100
rect 35532 23156 35588 23660
rect 35532 23090 35588 23100
rect 35736 23156 35792 23166
rect 35868 23156 35924 24220
rect 36092 24164 36148 24697
rect 36092 24098 36148 24108
rect 35980 24052 36036 24062
rect 35980 23958 36036 23996
rect 36204 23940 36260 25228
rect 36316 25218 36372 25228
rect 36876 25172 36932 25564
rect 36988 25478 37044 25490
rect 36988 25426 36990 25478
rect 37042 25426 37044 25478
rect 36988 25396 37044 25426
rect 36988 25330 37044 25340
rect 37100 25284 37156 25564
rect 37100 25218 37156 25228
rect 37436 25732 37492 25742
rect 37436 25284 37492 25676
rect 36876 25116 37044 25172
rect 36988 25060 37044 25116
rect 36988 25004 37156 25060
rect 36148 23908 36260 23940
rect 36148 23856 36150 23908
rect 36202 23884 36260 23908
rect 36316 23940 36372 23950
rect 36372 23884 36484 23940
rect 36202 23856 36204 23884
rect 36148 23844 36204 23856
rect 36316 23846 36372 23884
rect 35736 23154 35812 23156
rect 35736 23102 35738 23154
rect 35790 23102 35812 23154
rect 35736 23090 35812 23102
rect 35868 23100 36148 23156
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35084 22372 35140 22382
rect 35084 22278 35140 22316
rect 35644 21812 35700 21822
rect 34524 21756 35028 21812
rect 34860 21588 34916 21598
rect 33964 21084 34468 21140
rect 33740 21074 33796 21084
rect 33292 20862 33294 20914
rect 33346 20862 33348 20914
rect 33292 20850 33348 20862
rect 32956 20738 33012 20748
rect 33516 20804 33572 20814
rect 32396 20188 33218 20244
rect 33162 20130 33218 20188
rect 33162 20078 33164 20130
rect 33216 20078 33218 20130
rect 33162 20066 33218 20078
rect 32172 19730 32228 19740
rect 33404 20018 33460 20030
rect 33404 19966 33406 20018
rect 33458 19966 33460 20018
rect 33404 19012 33460 19966
rect 33404 18946 33460 18956
rect 31724 18498 31780 18508
rect 32060 18676 32116 18686
rect 32060 18450 32116 18620
rect 32060 18398 32062 18450
rect 32114 18398 32116 18450
rect 32060 18386 32116 18398
rect 33516 18450 33572 20748
rect 34412 20692 34468 21084
rect 34412 20636 34562 20692
rect 33908 20580 33964 20590
rect 33908 20074 33964 20524
rect 33908 20022 33910 20074
rect 33962 20022 33964 20074
rect 34506 20130 34562 20636
rect 34506 20078 34508 20130
rect 34560 20078 34562 20130
rect 34506 20066 34562 20078
rect 34748 20356 34804 20366
rect 33908 20010 33964 20022
rect 34076 20020 34132 20030
rect 34748 20020 34804 20300
rect 34076 19236 34132 19964
rect 34636 20018 34804 20020
rect 34636 19966 34750 20018
rect 34802 19966 34804 20018
rect 34636 19964 34804 19966
rect 33852 19180 34132 19236
rect 34188 19234 34244 19246
rect 34188 19182 34190 19234
rect 34242 19182 34244 19234
rect 33516 18398 33518 18450
rect 33570 18398 33572 18450
rect 33516 18386 33572 18398
rect 33740 19012 33796 19022
rect 32396 18228 32452 18238
rect 32396 18134 32452 18172
rect 31724 18004 31780 18014
rect 31724 17666 31780 17948
rect 31836 17834 31892 17846
rect 31836 17782 31838 17834
rect 31890 17782 31892 17834
rect 31836 17780 31892 17782
rect 31836 17714 31892 17724
rect 32060 17836 32340 17892
rect 31724 17614 31726 17666
rect 31778 17614 31780 17666
rect 31724 17556 31780 17614
rect 31724 17490 31780 17500
rect 31612 17276 31780 17332
rect 31164 17108 31220 17118
rect 31052 16324 31108 16334
rect 31052 16098 31108 16268
rect 31052 16046 31054 16098
rect 31106 16046 31108 16098
rect 31052 16034 31108 16046
rect 31052 15316 31108 15326
rect 31052 15222 31108 15260
rect 30940 15092 31108 15148
rect 30828 15026 30884 15036
rect 30716 14700 30996 14756
rect 30604 14532 30772 14588
rect 30604 14420 30660 14430
rect 30604 14326 30660 14364
rect 30380 13580 30548 13636
rect 28700 13356 29092 13412
rect 29036 12962 29092 13356
rect 29372 13188 29428 13198
rect 29372 13094 29428 13132
rect 29036 12910 29038 12962
rect 29090 12910 29092 12962
rect 29036 12898 29092 12910
rect 30268 12964 30324 12974
rect 30380 12964 30436 13580
rect 30604 13524 30660 13534
rect 30268 12962 30436 12964
rect 30268 12910 30270 12962
rect 30322 12910 30436 12962
rect 30268 12908 30436 12910
rect 30492 13468 30604 13524
rect 30268 12898 30324 12908
rect 29708 12740 29764 12750
rect 28868 12404 28924 12414
rect 28924 12348 29092 12404
rect 28868 12310 28924 12348
rect 28700 11396 28756 11406
rect 28588 11394 28756 11396
rect 28588 11342 28702 11394
rect 28754 11342 28756 11394
rect 28588 11340 28756 11342
rect 28700 11330 28756 11340
rect 29036 11394 29092 12348
rect 29036 11342 29038 11394
rect 29090 11342 29092 11394
rect 29036 11330 29092 11342
rect 29708 12178 29764 12684
rect 29708 12126 29710 12178
rect 29762 12126 29764 12178
rect 28476 10500 28532 10510
rect 28476 10406 28532 10444
rect 27804 10332 28308 10388
rect 26012 10210 26068 10220
rect 27112 10276 27168 10286
rect 25900 9996 26068 10052
rect 25228 8318 25230 8370
rect 25282 8318 25284 8370
rect 25228 8306 25284 8318
rect 25564 8316 25676 8372
rect 25564 7586 25620 8316
rect 25676 8278 25732 8316
rect 25900 9042 25956 9054
rect 25900 8990 25902 9042
rect 25954 8990 25956 9042
rect 25770 8148 25826 8158
rect 25770 8054 25826 8092
rect 25900 7924 25956 8990
rect 26012 8258 26068 9996
rect 26236 9826 26292 9838
rect 26236 9774 26238 9826
rect 26290 9774 26292 9826
rect 26236 9604 26292 9774
rect 27112 9826 27168 10220
rect 27112 9774 27114 9826
rect 27166 9774 27168 9826
rect 27112 9762 27168 9774
rect 26236 9538 26292 9548
rect 27356 9714 27412 9726
rect 27356 9662 27358 9714
rect 27410 9662 27412 9714
rect 26012 8206 26014 8258
rect 26066 8206 26068 8258
rect 26684 8372 26740 8382
rect 26684 8258 26740 8316
rect 26012 8148 26068 8206
rect 26012 8082 26068 8092
rect 26516 8202 26572 8214
rect 26516 8150 26518 8202
rect 26570 8150 26572 8202
rect 25900 7858 25956 7868
rect 26516 7812 26572 8150
rect 26684 8206 26686 8258
rect 26738 8206 26740 8258
rect 26684 8036 26740 8206
rect 26684 7970 26740 7980
rect 27188 8148 27244 8158
rect 27188 8034 27244 8092
rect 27188 7982 27190 8034
rect 27242 7982 27244 8034
rect 25564 7534 25566 7586
rect 25618 7534 25620 7586
rect 25564 7522 25620 7534
rect 26124 7756 26572 7812
rect 27020 7924 27076 7934
rect 25732 7418 25788 7430
rect 25732 7366 25734 7418
rect 25786 7366 25788 7418
rect 25732 6916 25788 7366
rect 26124 7252 26180 7756
rect 26236 7588 26292 7598
rect 26236 7474 26292 7532
rect 26236 7422 26238 7474
rect 26290 7422 26292 7474
rect 26236 7410 26292 7422
rect 26908 7474 26964 7486
rect 26908 7422 26910 7474
rect 26962 7422 26964 7474
rect 26478 7252 26534 7262
rect 26031 7196 26180 7252
rect 26236 7250 26534 7252
rect 26236 7198 26480 7250
rect 26532 7198 26534 7250
rect 26236 7196 26534 7198
rect 25116 6638 25118 6690
rect 25170 6638 25172 6690
rect 25116 6626 25172 6638
rect 25452 6860 25788 6916
rect 25900 7028 25956 7038
rect 24556 5966 24558 6018
rect 24610 5966 24612 6018
rect 24556 5954 24612 5966
rect 25340 6020 25396 6030
rect 24444 5182 24446 5234
rect 24498 5182 24500 5234
rect 24444 5170 24500 5182
rect 25004 5908 25060 5918
rect 25004 5234 25060 5852
rect 25340 5906 25396 5964
rect 25340 5854 25342 5906
rect 25394 5854 25396 5906
rect 25340 5842 25396 5854
rect 25452 5908 25508 6860
rect 25788 6580 25844 6590
rect 25788 6486 25844 6524
rect 25900 6244 25956 6972
rect 26031 6634 26087 7196
rect 26031 6582 26033 6634
rect 26085 6582 26087 6634
rect 26031 6468 26087 6582
rect 26031 6402 26087 6412
rect 26236 6356 26292 7196
rect 26478 7186 26534 7196
rect 26908 7028 26964 7422
rect 27020 7362 27076 7868
rect 27188 7924 27244 7982
rect 27188 7858 27244 7868
rect 27020 7310 27022 7362
rect 27074 7310 27076 7362
rect 27020 7298 27076 7310
rect 27244 7501 27300 7513
rect 27244 7449 27246 7501
rect 27298 7449 27300 7501
rect 26908 6962 26964 6972
rect 27244 7028 27300 7449
rect 27356 7476 27412 9662
rect 27636 8036 27692 8046
rect 27636 7942 27692 7980
rect 27580 7476 27636 7486
rect 27356 7474 27636 7476
rect 27356 7422 27582 7474
rect 27634 7422 27636 7474
rect 27356 7420 27636 7422
rect 27580 7410 27636 7420
rect 27804 7252 27860 10332
rect 29148 9042 29204 9054
rect 29484 9044 29540 9054
rect 29148 8990 29150 9042
rect 29202 8990 29204 9042
rect 29148 8932 29204 8990
rect 29148 8866 29204 8876
rect 29372 9042 29540 9044
rect 29372 8990 29486 9042
rect 29538 8990 29540 9042
rect 29372 8988 29540 8990
rect 28812 8818 28868 8830
rect 28812 8766 28814 8818
rect 28866 8766 28868 8818
rect 28812 8148 28868 8766
rect 29260 8260 29316 8270
rect 29260 8166 29316 8204
rect 28812 8082 28868 8092
rect 28644 8036 28700 8046
rect 28644 7698 28700 7980
rect 29372 7924 29428 8988
rect 29484 8978 29540 8988
rect 29708 8932 29764 12126
rect 30492 12178 30548 13468
rect 30604 13458 30660 13468
rect 30604 13188 30660 13198
rect 30604 13094 30660 13132
rect 30492 12126 30494 12178
rect 30546 12126 30548 12178
rect 30492 12114 30548 12126
rect 30716 11732 30772 14532
rect 30940 14530 30996 14700
rect 30940 14478 30942 14530
rect 30994 14478 30996 14530
rect 30940 13300 30996 14478
rect 31052 13412 31108 15092
rect 31164 14420 31220 17052
rect 31388 16884 31444 16894
rect 31388 16098 31444 16828
rect 31612 16884 31668 16894
rect 31612 16790 31668 16828
rect 31388 16046 31390 16098
rect 31442 16046 31444 16098
rect 31388 16034 31444 16046
rect 31500 16660 31556 16670
rect 31500 16266 31556 16604
rect 31500 16214 31502 16266
rect 31554 16214 31556 16266
rect 31500 15316 31556 16214
rect 31500 15250 31556 15260
rect 31388 15204 31444 15242
rect 31724 15148 31780 17276
rect 31836 16921 31892 16933
rect 31836 16869 31838 16921
rect 31890 16869 31892 16921
rect 31836 16660 31892 16869
rect 32060 16884 32116 17836
rect 32284 17834 32340 17836
rect 32284 17782 32286 17834
rect 32338 17782 32340 17834
rect 32284 17770 32340 17782
rect 32172 17666 32228 17678
rect 32172 17614 32174 17666
rect 32226 17614 32228 17666
rect 32172 17556 32228 17614
rect 32172 17490 32228 17500
rect 32508 17666 32564 17678
rect 32508 17614 32510 17666
rect 32562 17614 32564 17666
rect 32284 17444 32340 17454
rect 32284 16884 32340 17388
rect 32060 16818 32116 16828
rect 32172 16882 32340 16884
rect 32172 16830 32286 16882
rect 32338 16830 32340 16882
rect 32172 16828 32340 16830
rect 31948 16772 32004 16782
rect 31948 16678 32004 16716
rect 31836 16594 31892 16604
rect 31948 16548 32004 16558
rect 31948 16322 32004 16492
rect 31948 16270 31950 16322
rect 32002 16270 32004 16322
rect 31948 16258 32004 16270
rect 32004 15428 32060 15438
rect 32004 15334 32060 15372
rect 31388 15138 31444 15148
rect 31612 15092 31780 15148
rect 31332 14644 31388 14654
rect 31332 14550 31388 14588
rect 31164 14354 31220 14364
rect 31052 13346 31108 13356
rect 30940 13234 30996 13244
rect 31500 13076 31556 13086
rect 31500 12962 31556 13020
rect 31500 12910 31502 12962
rect 31554 12910 31556 12962
rect 31500 12898 31556 12910
rect 31164 12740 31220 12750
rect 31164 12646 31220 12684
rect 30716 11676 31108 11732
rect 29820 11394 29876 11406
rect 29820 11342 29822 11394
rect 29874 11342 29876 11394
rect 29820 11060 29876 11342
rect 29820 10994 29876 11004
rect 30940 10386 30996 10398
rect 30940 10334 30942 10386
rect 30994 10334 30996 10386
rect 30268 10164 30324 10174
rect 30268 10050 30324 10108
rect 30268 9998 30270 10050
rect 30322 9998 30324 10050
rect 30268 9986 30324 9998
rect 30604 9826 30660 9838
rect 30604 9774 30606 9826
rect 30658 9774 30660 9826
rect 30604 9716 30660 9774
rect 30604 9650 30660 9660
rect 30940 9044 30996 10334
rect 30940 8978 30996 8988
rect 29708 8866 29764 8876
rect 29820 8818 29876 8830
rect 29820 8766 29822 8818
rect 29874 8766 29876 8818
rect 29820 8372 29876 8766
rect 29820 8306 29876 8316
rect 28644 7646 28646 7698
rect 28698 7646 28700 7698
rect 27916 7476 27972 7486
rect 27916 7474 28532 7476
rect 27916 7422 27918 7474
rect 27970 7422 28532 7474
rect 27916 7420 28532 7422
rect 27916 7410 27972 7420
rect 27804 7196 27972 7252
rect 27244 6962 27300 6972
rect 26908 6692 26964 6702
rect 26908 6690 27188 6692
rect 26908 6638 26910 6690
rect 26962 6638 27188 6690
rect 26908 6636 27188 6638
rect 26908 6626 26964 6636
rect 26236 6300 26852 6356
rect 25900 6188 26516 6244
rect 26460 6018 26516 6188
rect 26460 5966 26462 6018
rect 26514 5966 26516 6018
rect 26460 5954 26516 5966
rect 25452 5842 25508 5852
rect 26216 5908 26272 5918
rect 26216 5814 26272 5852
rect 26796 5906 26852 6300
rect 26796 5854 26798 5906
rect 26850 5854 26852 5906
rect 26796 5842 26852 5854
rect 27132 5908 27188 6636
rect 27244 6690 27300 6702
rect 27244 6638 27246 6690
rect 27298 6638 27300 6690
rect 27244 6356 27300 6638
rect 27916 6356 27972 7196
rect 28364 7028 28420 7038
rect 28364 6914 28420 6972
rect 28364 6862 28366 6914
rect 28418 6862 28420 6914
rect 28364 6850 28420 6862
rect 28252 6804 28308 6814
rect 28120 6692 28176 6702
rect 28120 6598 28176 6636
rect 27244 6290 27300 6300
rect 27468 6300 27972 6356
rect 27132 5852 27300 5908
rect 27132 5682 27188 5694
rect 27132 5630 27134 5682
rect 27186 5630 27188 5682
rect 25004 5182 25006 5234
rect 25058 5182 25060 5234
rect 25004 5170 25060 5182
rect 26908 5236 26964 5246
rect 27132 5236 27188 5630
rect 26908 5234 27188 5236
rect 26908 5182 26910 5234
rect 26962 5182 27188 5234
rect 26908 5180 27188 5182
rect 26908 5170 26964 5180
rect 25788 5124 25844 5134
rect 25788 4900 25844 5068
rect 26796 5124 26852 5134
rect 25788 4844 26068 4900
rect 24332 4386 24388 4396
rect 26012 4338 26068 4844
rect 26012 4286 26014 4338
rect 26066 4286 26068 4338
rect 26012 4274 26068 4286
rect 26796 4338 26852 5068
rect 27244 4564 27300 5852
rect 27468 5236 27524 6300
rect 28252 6244 28308 6748
rect 28476 6580 28532 7420
rect 28644 6804 28700 7646
rect 29130 7868 29428 7924
rect 29932 8260 29988 8270
rect 29130 7586 29186 7868
rect 29130 7534 29132 7586
rect 29184 7534 29186 7586
rect 29130 7522 29186 7534
rect 29484 7588 29540 7598
rect 29932 7542 29988 8204
rect 30156 7924 30212 7934
rect 29372 7476 29428 7486
rect 29372 7382 29428 7420
rect 28644 6738 28700 6748
rect 29372 6692 29428 6702
rect 28476 6524 28868 6580
rect 28252 6188 28420 6244
rect 27692 6132 27748 6142
rect 27692 5906 27748 6076
rect 27692 5854 27694 5906
rect 27746 5854 27748 5906
rect 27692 5842 27748 5854
rect 28364 5348 28420 6188
rect 28812 6018 28868 6524
rect 28812 5966 28814 6018
rect 28866 5966 28868 6018
rect 28812 5954 28868 5966
rect 29372 6018 29428 6636
rect 29372 5966 29374 6018
rect 29426 5966 29428 6018
rect 29372 5954 29428 5966
rect 29484 6690 29540 7532
rect 29876 7530 29988 7542
rect 29876 7478 29878 7530
rect 29930 7478 29988 7530
rect 30044 7588 30100 7598
rect 30044 7494 30100 7532
rect 29876 7476 29988 7478
rect 29876 7466 29932 7476
rect 29484 6638 29486 6690
rect 29538 6638 29540 6690
rect 28568 5908 28624 5918
rect 28568 5814 28624 5852
rect 28252 5292 28420 5348
rect 27524 5180 27748 5236
rect 27468 5170 27524 5180
rect 27692 5122 27748 5180
rect 27692 5070 27694 5122
rect 27746 5070 27748 5122
rect 27692 5058 27748 5070
rect 28028 5124 28084 5134
rect 28028 5030 28084 5068
rect 27244 4498 27300 4508
rect 26796 4286 26798 4338
rect 26850 4286 26852 4338
rect 26796 4274 26852 4286
rect 25564 3780 25620 3790
rect 25564 3686 25620 3724
rect 27860 3668 27916 3678
rect 28252 3668 28308 5292
rect 28364 5122 28420 5134
rect 28364 5070 28366 5122
rect 28418 5070 28420 5122
rect 28364 3780 28420 5070
rect 28700 4452 28756 4462
rect 28588 4396 28700 4452
rect 29484 4452 29540 6638
rect 29652 6692 29708 6702
rect 29652 6598 29708 6636
rect 30156 6690 30212 7868
rect 31052 7588 31108 11676
rect 31612 10164 31668 15092
rect 32060 13748 32116 13758
rect 32042 13746 32116 13748
rect 32042 13694 32062 13746
rect 32114 13694 32116 13746
rect 32042 13682 32116 13694
rect 31724 13524 31780 13534
rect 31724 13430 31780 13468
rect 31724 13300 31780 13310
rect 31724 11620 31780 13244
rect 32042 13186 32098 13682
rect 32042 13134 32044 13186
rect 32096 13134 32098 13186
rect 32042 13122 32098 13134
rect 31724 11554 31780 11564
rect 31836 12180 31892 12190
rect 31724 11396 31780 11406
rect 31724 11282 31780 11340
rect 31724 11230 31726 11282
rect 31778 11230 31780 11282
rect 31724 10500 31780 11230
rect 31836 10637 31892 12124
rect 32172 11732 32228 16828
rect 32284 16818 32340 16828
rect 32508 16324 32564 17614
rect 32844 17668 32900 17678
rect 32844 17574 32900 17612
rect 33180 17444 33236 17454
rect 33180 17350 33236 17388
rect 32508 16258 32564 16268
rect 33740 16322 33796 18956
rect 33852 17780 33908 19180
rect 34020 19012 34076 19022
rect 34020 18918 34076 18956
rect 34058 17892 34114 17902
rect 34188 17892 34244 19182
rect 34524 19012 34580 19022
rect 34300 19010 34580 19012
rect 34300 18958 34526 19010
rect 34578 18958 34580 19010
rect 34300 18956 34580 18958
rect 34300 18450 34356 18956
rect 34524 18946 34580 18956
rect 34636 18676 34692 19964
rect 34748 19954 34804 19964
rect 34860 19234 34916 21532
rect 34860 19182 34862 19234
rect 34914 19182 34916 19234
rect 34860 19170 34916 19182
rect 34972 18788 35028 21756
rect 35644 21474 35700 21756
rect 35644 21422 35646 21474
rect 35698 21422 35700 21474
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 20916 35252 20926
rect 35196 20636 35252 20860
rect 35196 20580 35308 20636
rect 35084 20186 35140 20198
rect 35084 20134 35086 20186
rect 35138 20134 35140 20186
rect 35084 20020 35140 20134
rect 35252 20074 35308 20580
rect 35644 20580 35700 21422
rect 35756 20916 35812 23090
rect 35980 22932 36036 22942
rect 35980 22838 36036 22876
rect 35960 22314 36016 22326
rect 35960 22262 35962 22314
rect 36014 22262 36016 22314
rect 35960 21812 36016 22262
rect 35960 21746 36016 21756
rect 35756 20850 35812 20860
rect 35644 20514 35700 20524
rect 35812 20578 35868 20590
rect 35812 20526 35814 20578
rect 35866 20526 35868 20578
rect 35812 20356 35868 20526
rect 35812 20290 35868 20300
rect 35252 20022 35254 20074
rect 35306 20022 35308 20074
rect 35252 20010 35308 20022
rect 35868 20020 35924 20030
rect 35084 19954 35140 19964
rect 35532 19908 35588 19918
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 19348 35252 19358
rect 35532 19348 35588 19852
rect 35868 19458 35924 19964
rect 35868 19406 35870 19458
rect 35922 19406 35924 19458
rect 35868 19394 35924 19406
rect 35980 19906 36036 19918
rect 35980 19854 35982 19906
rect 36034 19854 36036 19906
rect 35196 19346 35588 19348
rect 35196 19294 35198 19346
rect 35250 19294 35588 19346
rect 35196 19292 35588 19294
rect 35196 19282 35252 19292
rect 35532 19234 35588 19292
rect 35980 19348 36036 19854
rect 35980 19282 36036 19292
rect 35532 19182 35534 19234
rect 35586 19182 35588 19234
rect 35532 19170 35588 19182
rect 34972 18732 35252 18788
rect 34300 18398 34302 18450
rect 34354 18398 34356 18450
rect 34300 18386 34356 18398
rect 34524 18620 34692 18676
rect 35196 18676 35252 18732
rect 35196 18620 35476 18676
rect 34058 17890 34244 17892
rect 34058 17838 34060 17890
rect 34112 17838 34244 17890
rect 34058 17836 34244 17838
rect 34300 17892 34356 17902
rect 34058 17826 34114 17836
rect 33852 17714 33908 17724
rect 34300 17666 34356 17836
rect 34300 17614 34302 17666
rect 34354 17614 34356 17666
rect 33740 16270 33742 16322
rect 33794 16270 33796 16322
rect 32284 16098 32340 16110
rect 32284 16046 32286 16098
rect 32338 16046 32340 16098
rect 32284 15876 32340 16046
rect 32676 15876 32732 15886
rect 32284 15874 32732 15876
rect 32284 15822 32678 15874
rect 32730 15822 32732 15874
rect 32284 15820 32732 15822
rect 32284 15428 32340 15820
rect 32676 15810 32732 15820
rect 32396 15428 32452 15438
rect 32284 15372 32396 15428
rect 32284 12964 32340 12974
rect 32284 12870 32340 12908
rect 32396 12404 32452 15372
rect 32956 15316 33012 15326
rect 32956 15222 33012 15260
rect 33292 15202 33348 15214
rect 33292 15150 33294 15202
rect 33346 15150 33348 15202
rect 33068 13746 33124 13758
rect 33068 13694 33070 13746
rect 33122 13694 33124 13746
rect 32956 13524 33012 13534
rect 32956 12962 33012 13468
rect 32788 12906 32844 12918
rect 32788 12854 32790 12906
rect 32842 12854 32844 12906
rect 32956 12910 32958 12962
rect 33010 12910 33012 12962
rect 32956 12898 33012 12910
rect 32788 12404 32844 12854
rect 33068 12740 33124 13694
rect 33292 13524 33348 15150
rect 33740 15148 33796 16270
rect 33628 15092 33796 15148
rect 34076 17556 34132 17566
rect 34076 16098 34132 17500
rect 34300 17108 34356 17614
rect 34524 17444 34580 18620
rect 35420 18228 35476 18620
rect 35868 18564 35924 18574
rect 35756 18340 35812 18350
rect 35420 18172 35644 18228
rect 35588 18116 35644 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 34804 17892 34860 17902
rect 34804 17722 34860 17836
rect 34804 17670 34806 17722
rect 34858 17670 34860 17722
rect 34804 17658 34860 17670
rect 34972 17780 35028 17790
rect 34972 17666 35028 17724
rect 35588 17722 35644 18060
rect 34972 17614 34974 17666
rect 35026 17614 35028 17666
rect 34972 17602 35028 17614
rect 35420 17668 35476 17678
rect 35588 17670 35590 17722
rect 35642 17670 35644 17722
rect 35588 17658 35644 17670
rect 35420 17574 35476 17612
rect 35756 17444 35812 18284
rect 35868 17668 35924 18508
rect 36092 18116 36148 23100
rect 36428 23154 36484 23884
rect 36428 23102 36430 23154
rect 36482 23102 36484 23154
rect 36428 23090 36484 23102
rect 37100 23044 37156 25004
rect 37436 24946 37492 25228
rect 37436 24894 37438 24946
rect 37490 24894 37492 24946
rect 37436 24882 37492 24894
rect 37548 24724 37604 26852
rect 37772 26404 37828 26414
rect 37772 26310 37828 26348
rect 37548 24658 37604 24668
rect 37660 26180 37716 26190
rect 37548 23938 37604 23950
rect 37548 23886 37550 23938
rect 37602 23886 37604 23938
rect 37548 23492 37604 23886
rect 37660 23770 37716 26124
rect 37996 25618 38052 25630
rect 37996 25566 37998 25618
rect 38050 25566 38052 25618
rect 37996 25508 38052 25566
rect 37996 25442 38052 25452
rect 38220 24276 38276 26852
rect 38556 26404 38612 26414
rect 38556 26290 38612 26348
rect 39432 26292 39488 26302
rect 38556 26238 38558 26290
rect 38610 26238 38612 26290
rect 38556 26226 38612 26238
rect 39228 26290 39488 26292
rect 39228 26238 39434 26290
rect 39486 26238 39488 26290
rect 39228 26236 39488 26238
rect 39228 24948 39284 26236
rect 39432 26226 39488 26236
rect 39676 26066 39732 26078
rect 39676 26014 39678 26066
rect 39730 26014 39732 26066
rect 39676 25060 39732 26014
rect 39900 25620 39956 29820
rect 41580 29652 41636 30716
rect 41132 29596 41636 29652
rect 40012 29453 40068 29465
rect 40012 29401 40014 29453
rect 40066 29401 40068 29453
rect 40908 29428 40964 29438
rect 40012 25732 40068 29401
rect 40796 29426 40964 29428
rect 40796 29374 40910 29426
rect 40962 29374 40964 29426
rect 40796 29372 40964 29374
rect 40572 28532 40628 28542
rect 40796 28532 40852 29372
rect 40908 29362 40964 29372
rect 40572 28530 40852 28532
rect 40572 28478 40574 28530
rect 40626 28478 40852 28530
rect 40572 28476 40852 28478
rect 40908 28642 40964 28654
rect 40908 28590 40910 28642
rect 40962 28590 40964 28642
rect 40572 28466 40628 28476
rect 40460 27860 40516 27870
rect 40236 27858 40516 27860
rect 40236 27806 40462 27858
rect 40514 27806 40516 27858
rect 40236 27804 40516 27806
rect 40236 26526 40292 27804
rect 40460 27794 40516 27804
rect 40180 26514 40292 26526
rect 40180 26462 40182 26514
rect 40234 26462 40292 26514
rect 40180 26460 40292 26462
rect 40684 27074 40740 28476
rect 40908 27310 40964 28590
rect 40852 27298 40964 27310
rect 40852 27246 40854 27298
rect 40906 27246 40964 27298
rect 40852 27244 40964 27246
rect 41020 28084 41076 28094
rect 40852 27234 40908 27244
rect 40684 27022 40686 27074
rect 40738 27022 40740 27074
rect 40180 26450 40236 26460
rect 40348 26292 40404 26302
rect 40348 26290 40516 26292
rect 40348 26238 40350 26290
rect 40402 26238 40516 26290
rect 40348 26236 40516 26238
rect 40348 26226 40404 26236
rect 40348 25732 40404 25742
rect 40012 25676 40292 25732
rect 39900 25564 40180 25620
rect 39788 25478 39844 25490
rect 39788 25426 39790 25478
rect 39842 25426 39844 25478
rect 39788 25284 39844 25426
rect 39788 25218 39844 25228
rect 39900 25396 39956 25406
rect 39900 25060 39956 25340
rect 39676 24994 39732 25004
rect 39788 25004 39956 25060
rect 38892 24892 39284 24948
rect 38220 24220 38500 24276
rect 38220 24052 38276 24062
rect 38220 23938 38276 23996
rect 37940 23882 37996 23894
rect 37940 23830 37942 23882
rect 37994 23830 37996 23882
rect 38220 23886 38222 23938
rect 38274 23886 38276 23938
rect 38220 23874 38276 23886
rect 37940 23828 37996 23830
rect 37940 23772 38164 23828
rect 37660 23718 37662 23770
rect 37714 23718 37716 23770
rect 37660 23706 37716 23718
rect 38108 23716 38164 23772
rect 38108 23660 38276 23716
rect 37548 23426 37604 23436
rect 38108 23492 38164 23502
rect 37304 23156 37360 23166
rect 37548 23156 37604 23166
rect 37996 23156 38052 23166
rect 37304 23154 37492 23156
rect 37304 23102 37306 23154
rect 37358 23102 37492 23154
rect 37304 23100 37492 23102
rect 37304 23090 37360 23100
rect 37100 22978 37156 22988
rect 37436 22820 37492 23100
rect 37548 23154 38052 23156
rect 37548 23102 37550 23154
rect 37602 23102 37998 23154
rect 38050 23102 38052 23154
rect 37548 23100 38052 23102
rect 37548 23090 37604 23100
rect 37996 23090 38052 23100
rect 38108 23042 38164 23436
rect 38108 22990 38110 23042
rect 38162 22990 38164 23042
rect 38108 22978 38164 22990
rect 37436 22764 37716 22820
rect 36204 22596 36260 22606
rect 36204 22502 36260 22540
rect 36988 22372 37044 22382
rect 36988 22278 37044 22316
rect 37660 19460 37716 22764
rect 38108 22708 38164 22718
rect 38108 22594 38164 22652
rect 38108 22542 38110 22594
rect 38162 22542 38164 22594
rect 38108 22530 38164 22542
rect 38220 22484 38276 23660
rect 38332 23181 38388 23193
rect 38332 23129 38334 23181
rect 38386 23129 38388 23181
rect 38332 22596 38388 23129
rect 38332 22530 38388 22540
rect 38220 22418 38276 22428
rect 37864 22316 37920 22326
rect 37864 22314 37940 22316
rect 37864 22262 37866 22314
rect 37918 22262 37940 22314
rect 37864 22250 37940 22262
rect 37772 21812 37828 21822
rect 37772 21698 37828 21756
rect 37772 21646 37774 21698
rect 37826 21646 37828 21698
rect 37772 21634 37828 21646
rect 37884 20132 37940 22250
rect 37548 19404 37716 19460
rect 37772 20076 37940 20132
rect 38444 20132 38500 24220
rect 38892 24164 38948 24892
rect 39116 24724 39172 24762
rect 39116 24658 39172 24668
rect 39788 24388 39844 25004
rect 39992 24724 40048 24734
rect 39992 24630 40048 24668
rect 39788 24332 40068 24388
rect 38892 24108 39172 24164
rect 38911 23882 38967 23894
rect 38668 23828 38724 23838
rect 38911 23830 38913 23882
rect 38965 23830 38967 23882
rect 38668 23826 38836 23828
rect 38668 23774 38670 23826
rect 38722 23774 38836 23826
rect 38668 23772 38836 23774
rect 38668 23762 38724 23772
rect 38668 23154 38724 23166
rect 38668 23102 38670 23154
rect 38722 23102 38724 23154
rect 38556 22932 38612 22942
rect 38556 22370 38612 22876
rect 38668 22708 38724 23102
rect 38668 22642 38724 22652
rect 38668 22484 38724 22494
rect 38668 22390 38724 22428
rect 38556 22318 38558 22370
rect 38610 22318 38612 22370
rect 38556 22306 38612 22318
rect 38780 22372 38836 23772
rect 38911 23380 38967 23830
rect 38892 23324 38967 23380
rect 38892 22708 38948 23324
rect 38892 22642 38948 22652
rect 39004 23154 39060 23166
rect 39004 23102 39006 23154
rect 39058 23102 39060 23154
rect 39004 22596 39060 23102
rect 39004 22530 39060 22540
rect 38780 22316 38892 22372
rect 38836 22314 38892 22316
rect 38836 22262 38838 22314
rect 38890 22262 38892 22314
rect 38836 22250 38892 22262
rect 38556 21812 38612 21822
rect 38556 21252 38612 21756
rect 39116 21812 39172 24108
rect 39676 23940 39732 23950
rect 39676 23380 39732 23884
rect 39788 23940 39844 23950
rect 40012 23940 40068 24332
rect 39788 23938 40068 23940
rect 39788 23886 39790 23938
rect 39842 23886 40068 23938
rect 39788 23884 40068 23886
rect 39788 23874 39844 23884
rect 39228 23324 39732 23380
rect 39228 22370 39284 23324
rect 39228 22318 39230 22370
rect 39282 22318 39284 22370
rect 39228 22306 39284 22318
rect 39452 23154 39508 23166
rect 39452 23102 39454 23154
rect 39506 23102 39508 23154
rect 39116 21746 39172 21756
rect 39452 21252 39508 23102
rect 39788 22930 39844 22942
rect 39788 22878 39790 22930
rect 39842 22878 39844 22930
rect 39676 22372 39732 22382
rect 38556 21196 38724 21252
rect 38668 21140 38724 21196
rect 38612 21084 38724 21140
rect 39340 21196 39508 21252
rect 39564 22370 39732 22372
rect 39564 22318 39678 22370
rect 39730 22318 39732 22370
rect 39564 22316 39732 22318
rect 39564 21588 39620 22316
rect 39676 22306 39732 22316
rect 38612 20858 38668 21084
rect 39340 20926 39396 21196
rect 39340 20914 39414 20926
rect 39340 20862 39360 20914
rect 39412 20862 39414 20914
rect 39340 20860 39414 20862
rect 38612 20806 38614 20858
rect 38666 20806 38668 20858
rect 39358 20850 39414 20860
rect 38612 20794 38668 20806
rect 39116 20802 39172 20814
rect 39116 20750 39118 20802
rect 39170 20750 39172 20802
rect 37156 19348 37212 19358
rect 37156 19290 37212 19292
rect 36988 19236 37044 19246
rect 37156 19238 37158 19290
rect 37210 19238 37212 19290
rect 37156 19226 37212 19238
rect 36988 19122 37044 19180
rect 36988 19070 36990 19122
rect 37042 19070 37044 19122
rect 36988 18564 37044 19070
rect 36988 18498 37044 18508
rect 36204 18452 36260 18462
rect 37548 18452 37604 19404
rect 37772 19348 37828 20076
rect 38444 20066 38500 20076
rect 38780 20692 38836 20702
rect 38780 20634 38836 20636
rect 38780 20582 38782 20634
rect 38834 20582 38836 20634
rect 38668 20020 38724 20030
rect 37884 19908 37940 19918
rect 37884 19906 38612 19908
rect 37884 19854 37886 19906
rect 37938 19854 38612 19906
rect 37884 19852 38612 19854
rect 37884 19842 37940 19852
rect 38556 19458 38612 19852
rect 38556 19406 38558 19458
rect 38610 19406 38612 19458
rect 38556 19394 38612 19406
rect 37772 19282 37828 19292
rect 38668 19348 38724 19964
rect 38668 19282 38724 19292
rect 37660 19234 37716 19246
rect 37660 19182 37662 19234
rect 37714 19182 37716 19234
rect 37660 18676 37716 19182
rect 37902 19236 37958 19246
rect 38220 19236 38276 19246
rect 37902 19234 38276 19236
rect 37902 19182 37904 19234
rect 37956 19182 38222 19234
rect 38274 19182 38276 19234
rect 37902 19180 38276 19182
rect 37902 19170 37958 19180
rect 38220 19170 38276 19180
rect 38780 19236 38836 20582
rect 38780 19170 38836 19180
rect 37660 18610 37716 18620
rect 36260 18396 36372 18452
rect 36204 18358 36260 18396
rect 36092 18060 36260 18116
rect 35868 17602 35924 17612
rect 36092 17668 36148 17678
rect 36092 17574 36148 17612
rect 34524 17388 35252 17444
rect 34300 17042 34356 17052
rect 34076 16046 34078 16098
rect 34130 16046 34132 16098
rect 34076 15148 34132 16046
rect 34188 16884 34244 16894
rect 34188 16098 34244 16828
rect 34188 16046 34190 16098
rect 34242 16046 34244 16098
rect 34188 16034 34244 16046
rect 34524 15988 34580 15998
rect 34524 15894 34580 15932
rect 34076 15092 34244 15148
rect 33628 13636 33684 15092
rect 34188 14530 34244 15092
rect 34188 14478 34190 14530
rect 34242 14478 34244 14530
rect 34188 14466 34244 14478
rect 34524 15090 34580 15102
rect 34524 15038 34526 15090
rect 34578 15038 34580 15090
rect 33852 14308 33908 14318
rect 33292 13458 33348 13468
rect 33516 13580 33684 13636
rect 33740 14306 33908 14308
rect 33740 14254 33854 14306
rect 33906 14254 33908 14306
rect 33740 14252 33908 14254
rect 33516 13086 33572 13580
rect 33460 13074 33572 13086
rect 33460 13022 33462 13074
rect 33514 13022 33572 13074
rect 33460 13020 33572 13022
rect 33628 13412 33684 13422
rect 33460 12964 33516 13020
rect 33460 12898 33516 12908
rect 33068 12674 33124 12684
rect 31836 10585 31838 10637
rect 31890 10585 31892 10637
rect 31836 10573 31892 10585
rect 32060 11676 32228 11732
rect 32284 12348 32452 12404
rect 32732 12348 32844 12404
rect 31724 10444 31892 10500
rect 31612 10098 31668 10108
rect 31444 9994 31500 10006
rect 31444 9942 31446 9994
rect 31498 9942 31500 9994
rect 31444 9940 31500 9942
rect 31444 9884 31780 9940
rect 31724 9826 31780 9884
rect 31612 9770 31668 9782
rect 31612 9718 31614 9770
rect 31666 9718 31668 9770
rect 31724 9774 31726 9826
rect 31778 9774 31780 9826
rect 31724 9762 31780 9774
rect 31612 9604 31668 9718
rect 31836 9604 31892 10444
rect 31612 9548 31892 9604
rect 31948 9044 32004 9054
rect 31948 8950 32004 8988
rect 31164 8372 31220 8382
rect 31164 8278 31220 8316
rect 31948 8258 32004 8270
rect 31948 8206 31950 8258
rect 32002 8206 32004 8258
rect 31948 8148 32004 8206
rect 32060 8260 32116 11676
rect 32284 11508 32340 12348
rect 32172 11452 32340 11508
rect 32396 12068 32452 12078
rect 32732 12068 32788 12348
rect 33628 12205 33684 13356
rect 33628 12153 33630 12205
rect 33682 12153 33684 12205
rect 33628 12141 33684 12153
rect 33740 12852 33796 14252
rect 33852 14242 33908 14252
rect 34524 13972 34580 15038
rect 33964 13916 34580 13972
rect 34636 13972 34692 17388
rect 34804 17108 34860 17118
rect 34804 17014 34860 17052
rect 35196 17106 35252 17388
rect 35196 17054 35198 17106
rect 35250 17054 35252 17106
rect 35196 17042 35252 17054
rect 35532 17388 35812 17444
rect 34972 16884 35028 16894
rect 34860 15316 34916 15326
rect 34972 15316 35028 16828
rect 35532 16882 35588 17388
rect 35980 17108 36036 17118
rect 35532 16830 35534 16882
rect 35586 16830 35588 16882
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35532 16100 35588 16830
rect 35644 16884 35700 16894
rect 35644 16790 35700 16828
rect 35644 16100 35700 16110
rect 35532 16098 35700 16100
rect 35532 16046 35646 16098
rect 35698 16046 35700 16098
rect 35532 16044 35700 16046
rect 35644 16034 35700 16044
rect 35308 15876 35364 15886
rect 35308 15782 35364 15820
rect 34860 15314 35028 15316
rect 34860 15262 34862 15314
rect 34914 15262 35028 15314
rect 34860 15260 35028 15262
rect 35196 15314 35252 15326
rect 35196 15262 35198 15314
rect 35250 15262 35252 15314
rect 34860 15250 34916 15260
rect 35196 15148 35252 15262
rect 34954 15092 35252 15148
rect 35532 15092 35588 15102
rect 34954 14754 35010 15092
rect 35532 14998 35588 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34954 14702 34956 14754
rect 35008 14702 35010 14754
rect 34954 14690 35010 14702
rect 35196 14532 35252 14542
rect 35980 14532 36036 17052
rect 35196 14438 35252 14476
rect 35700 14474 35756 14486
rect 35700 14422 35702 14474
rect 35754 14422 35756 14474
rect 35980 14466 36036 14476
rect 35700 14308 35756 14422
rect 35700 14242 35756 14252
rect 35868 14420 35924 14430
rect 34636 13916 35028 13972
rect 32396 12066 32788 12068
rect 32396 12014 32398 12066
rect 32450 12014 32788 12066
rect 32396 12012 32788 12014
rect 32172 9380 32228 11452
rect 32284 11350 32340 11362
rect 32284 11298 32286 11350
rect 32338 11298 32340 11350
rect 32284 11284 32340 11298
rect 32284 11218 32340 11228
rect 32396 11172 32452 12012
rect 32508 11396 32564 11406
rect 32508 11302 32564 11340
rect 33068 11396 33124 11406
rect 32396 11106 32452 11116
rect 32508 11226 32564 11238
rect 32508 11174 32510 11226
rect 32562 11174 32564 11226
rect 32508 11060 32564 11174
rect 32508 10994 32564 11004
rect 32620 10724 32676 10734
rect 32620 10610 32676 10668
rect 32620 10558 32622 10610
rect 32674 10558 32676 10610
rect 32620 10546 32676 10558
rect 33068 10610 33124 11340
rect 33068 10558 33070 10610
rect 33122 10558 33124 10610
rect 33068 10546 33124 10558
rect 32452 10388 32508 10398
rect 32396 10386 32508 10388
rect 32396 10334 32454 10386
rect 32506 10334 32508 10386
rect 32396 10322 32508 10334
rect 32620 10388 32676 10398
rect 32396 9604 32452 10322
rect 32508 9940 32564 9950
rect 32620 9940 32676 10332
rect 32508 9938 32676 9940
rect 32508 9886 32510 9938
rect 32562 9886 32676 9938
rect 32508 9884 32676 9886
rect 32508 9874 32564 9884
rect 32396 9548 33572 9604
rect 32172 9314 32228 9324
rect 33516 9042 33572 9548
rect 33516 8990 33518 9042
rect 33570 8990 33572 9042
rect 33516 8978 33572 8990
rect 32956 8932 33012 8942
rect 32284 8818 32340 8830
rect 32284 8766 32286 8818
rect 32338 8766 32340 8818
rect 32284 8260 32340 8766
rect 32060 8204 32228 8260
rect 32004 8092 32116 8148
rect 31948 8082 32004 8092
rect 31052 7522 31108 7532
rect 30156 6638 30158 6690
rect 30210 6638 30212 6690
rect 30156 6468 30212 6638
rect 30156 6402 30212 6412
rect 30268 7474 30324 7486
rect 30268 7422 30270 7474
rect 30322 7422 30324 7474
rect 30268 6132 30324 7422
rect 30604 7252 30660 7262
rect 30604 7250 31556 7252
rect 30604 7198 30606 7250
rect 30658 7198 31556 7250
rect 30604 7196 31556 7198
rect 30604 7186 30660 7196
rect 30398 6692 30454 6702
rect 30716 6692 30772 6702
rect 30398 6690 30772 6692
rect 30398 6638 30400 6690
rect 30452 6638 30718 6690
rect 30770 6638 30772 6690
rect 30398 6636 30772 6638
rect 30398 6626 30454 6636
rect 30716 6626 30772 6636
rect 31052 6468 31108 6478
rect 31052 6466 31332 6468
rect 31052 6414 31054 6466
rect 31106 6414 31332 6466
rect 31052 6412 31332 6414
rect 31052 6402 31108 6412
rect 30156 6076 30324 6132
rect 29596 5908 29652 5918
rect 29596 5236 29652 5852
rect 30156 5572 30212 6076
rect 31276 5906 31332 6412
rect 31276 5854 31278 5906
rect 31330 5854 31332 5906
rect 31276 5842 31332 5854
rect 30156 5516 30436 5572
rect 29596 5234 29764 5236
rect 29596 5182 29598 5234
rect 29650 5182 29764 5234
rect 29596 5180 29764 5182
rect 29596 5170 29652 5180
rect 29708 4900 29764 5180
rect 30380 4900 30436 5516
rect 31500 5234 31556 7196
rect 31668 6468 31724 6478
rect 31668 6374 31724 6412
rect 32060 5908 32116 8092
rect 32172 6132 32228 8204
rect 32284 8194 32340 8204
rect 32172 6066 32228 6076
rect 32060 5906 32340 5908
rect 32060 5854 32062 5906
rect 32114 5854 32340 5906
rect 32060 5852 32340 5854
rect 32060 5842 32116 5852
rect 31500 5182 31502 5234
rect 31554 5182 31556 5234
rect 31500 5170 31556 5182
rect 32284 5122 32340 5852
rect 32284 5070 32286 5122
rect 32338 5070 32340 5122
rect 29708 4844 29820 4900
rect 30380 4844 30566 4900
rect 29596 4452 29652 4462
rect 29484 4450 29652 4452
rect 29484 4398 29598 4450
rect 29650 4398 29652 4450
rect 29484 4396 29652 4398
rect 28588 4116 28644 4396
rect 28700 4358 28756 4396
rect 29596 4386 29652 4396
rect 29764 4394 29820 4844
rect 28364 3714 28420 3724
rect 28532 4060 28644 4116
rect 29036 4340 29092 4350
rect 29764 4342 29766 4394
rect 29818 4342 29820 4394
rect 30510 4450 30566 4844
rect 30510 4398 30512 4450
rect 30564 4398 30566 4450
rect 30510 4386 30566 4398
rect 29764 4330 29820 4342
rect 30268 4340 30324 4350
rect 27860 3666 28308 3668
rect 27860 3614 27862 3666
rect 27914 3614 28308 3666
rect 27860 3612 28308 3614
rect 27860 3602 27916 3612
rect 24108 3490 24164 3500
rect 24556 3556 24612 3566
rect 28252 3556 28308 3612
rect 28532 3610 28588 4060
rect 28364 3556 28420 3566
rect 28252 3554 28420 3556
rect 28252 3502 28366 3554
rect 28418 3502 28420 3554
rect 28532 3558 28534 3610
rect 28586 3558 28588 3610
rect 28532 3546 28588 3558
rect 29036 3554 29092 4284
rect 30268 4246 30324 4284
rect 29278 3780 29334 3790
rect 29278 3686 29334 3724
rect 32284 3778 32340 5070
rect 32956 5122 33012 8876
rect 33740 8372 33796 12796
rect 33852 13634 33908 13646
rect 33852 13582 33854 13634
rect 33906 13582 33908 13634
rect 33852 12404 33908 13582
rect 33852 12338 33908 12348
rect 33964 12068 34020 13916
rect 34076 13524 34132 13534
rect 34076 12964 34132 13468
rect 34188 12964 34244 12974
rect 34076 12962 34244 12964
rect 34076 12910 34190 12962
rect 34242 12910 34244 12962
rect 34076 12908 34244 12910
rect 34188 12898 34244 12908
rect 34356 12964 34412 12974
rect 34356 12870 34412 12908
rect 34860 12964 34916 12974
rect 34972 12964 35028 13916
rect 35756 13634 35812 13646
rect 35756 13582 35758 13634
rect 35810 13582 35812 13634
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35756 13188 35812 13582
rect 35868 13524 35924 14364
rect 35868 13458 35924 13468
rect 35980 14308 36036 14318
rect 35980 13636 36036 14252
rect 35980 13300 36036 13580
rect 34860 12962 35028 12964
rect 34860 12910 34862 12962
rect 34914 12910 35028 12962
rect 34860 12908 35028 12910
rect 34860 12898 34916 12908
rect 34972 12740 35028 12908
rect 35420 13132 35812 13188
rect 35868 13244 36036 13300
rect 36092 13972 36148 13982
rect 36092 13746 36148 13916
rect 36092 13694 36094 13746
rect 36146 13694 36148 13746
rect 35420 12964 35476 13132
rect 34972 12674 35028 12684
rect 35102 12850 35158 12862
rect 35102 12798 35104 12850
rect 35156 12798 35158 12850
rect 35102 12516 35158 12798
rect 35102 12450 35158 12460
rect 35420 12292 35476 12908
rect 35756 12964 35812 12974
rect 35756 12870 35812 12908
rect 35588 12740 35644 12750
rect 35868 12740 35924 13244
rect 36092 13076 36148 13694
rect 36092 13010 36148 13020
rect 35420 12226 35476 12236
rect 35532 12738 35644 12740
rect 35532 12686 35590 12738
rect 35642 12686 35644 12738
rect 35532 12674 35644 12686
rect 35756 12684 35924 12740
rect 35980 12964 36036 12974
rect 36204 12964 36260 18060
rect 36316 17892 36372 18396
rect 37548 18386 37604 18396
rect 36764 18338 36820 18350
rect 36764 18286 36766 18338
rect 36818 18286 36820 18338
rect 36764 18116 36820 18286
rect 36764 18050 36820 18060
rect 38668 18338 38724 18350
rect 38668 18286 38670 18338
rect 38722 18286 38724 18338
rect 36316 17826 36372 17836
rect 37212 17892 37268 17902
rect 37212 17798 37268 17836
rect 38668 17892 38724 18286
rect 38668 17826 38724 17836
rect 36334 17668 36390 17678
rect 36876 17668 36932 17678
rect 36334 17666 36932 17668
rect 36334 17614 36336 17666
rect 36388 17614 36878 17666
rect 36930 17614 36932 17666
rect 36334 17612 36932 17614
rect 36334 17602 36390 17612
rect 36876 17602 36932 17612
rect 39116 16884 39172 20750
rect 39564 19908 39620 21532
rect 39676 21588 39732 21598
rect 39788 21588 39844 22878
rect 39676 21586 39844 21588
rect 39676 21534 39678 21586
rect 39730 21534 39844 21586
rect 39676 21532 39844 21534
rect 40012 22036 40068 22046
rect 39676 21522 39732 21532
rect 39882 20692 39938 20702
rect 39882 20690 39956 20692
rect 39882 20638 39884 20690
rect 39936 20638 39956 20690
rect 39882 20626 39956 20638
rect 39900 20018 39956 20626
rect 39900 19966 39902 20018
rect 39954 19966 39956 20018
rect 39900 19954 39956 19966
rect 39564 19842 39620 19852
rect 39770 19460 39826 19470
rect 40012 19460 40068 21980
rect 40124 21364 40180 25564
rect 40236 24948 40292 25676
rect 40236 24882 40292 24892
rect 40236 24498 40292 24510
rect 40236 24446 40238 24498
rect 40290 24446 40292 24498
rect 40236 23940 40292 24446
rect 40236 23874 40292 23884
rect 40348 23938 40404 25676
rect 40348 23886 40350 23938
rect 40402 23886 40404 23938
rect 40348 23874 40404 23886
rect 40460 25508 40516 26236
rect 40460 23604 40516 25452
rect 40684 25396 40740 27022
rect 40796 25620 40852 25630
rect 40796 25526 40852 25564
rect 40684 25330 40740 25340
rect 40908 25396 40964 25406
rect 40684 25060 40740 25070
rect 40684 23938 40740 25004
rect 40684 23886 40686 23938
rect 40738 23886 40740 23938
rect 40684 23874 40740 23886
rect 40908 23899 40964 25340
rect 41020 24749 41076 28028
rect 41132 27858 41188 29596
rect 41244 29441 41300 29453
rect 41244 29389 41246 29441
rect 41298 29389 41300 29441
rect 41244 29316 41300 29389
rect 41244 28644 41300 29260
rect 41356 29314 41412 29326
rect 41356 29262 41358 29314
rect 41410 29262 41412 29314
rect 41356 28756 41412 29262
rect 41692 28868 41748 30940
rect 42364 30994 42420 33180
rect 42364 30942 42366 30994
rect 42418 30942 42420 30994
rect 42364 30930 42420 30942
rect 41916 30772 41972 30782
rect 41916 29453 41972 30716
rect 42364 30212 42420 30222
rect 42476 30212 42532 33294
rect 43148 33012 43204 33022
rect 43148 32450 43204 32956
rect 43148 32398 43150 32450
rect 43202 32398 43204 32450
rect 43148 32386 43204 32398
rect 43260 31892 43316 35756
rect 43484 35588 43540 35598
rect 43484 34914 43540 35532
rect 43484 34862 43486 34914
rect 43538 34862 43540 34914
rect 43484 34850 43540 34862
rect 43484 34018 43540 34030
rect 43484 33966 43486 34018
rect 43538 33966 43540 34018
rect 43484 33348 43540 33966
rect 43708 33348 43764 33358
rect 43484 33346 43764 33348
rect 43484 33294 43710 33346
rect 43762 33294 43764 33346
rect 43484 33292 43764 33294
rect 43708 33282 43764 33292
rect 43372 33124 43428 33134
rect 43372 33122 43876 33124
rect 43372 33070 43374 33122
rect 43426 33070 43876 33122
rect 43372 33068 43876 33070
rect 43372 33058 43428 33068
rect 43820 32589 43876 33068
rect 43820 32537 43822 32589
rect 43874 32537 43876 32589
rect 43820 32525 43876 32537
rect 43260 31826 43316 31836
rect 42868 31556 42924 31566
rect 42868 31554 42980 31556
rect 42868 31502 42870 31554
rect 42922 31502 42980 31554
rect 42868 31490 42980 31502
rect 42700 30772 42756 30782
rect 42700 30678 42756 30716
rect 42364 30210 42532 30212
rect 42364 30158 42366 30210
rect 42418 30158 42532 30210
rect 42364 30156 42532 30158
rect 42924 30324 42980 31490
rect 42364 30146 42420 30156
rect 42924 29998 42980 30268
rect 42924 29988 43036 29998
rect 42924 29986 43092 29988
rect 42924 29934 42982 29986
rect 43034 29934 43092 29986
rect 42924 29932 43092 29934
rect 42980 29922 43092 29932
rect 41916 29401 41918 29453
rect 41970 29401 41972 29453
rect 41916 29389 41972 29401
rect 41692 28802 41748 28812
rect 41356 28690 41412 28700
rect 41244 28578 41300 28588
rect 41692 28642 41748 28654
rect 41692 28590 41694 28642
rect 41746 28590 41748 28642
rect 41132 27806 41134 27858
rect 41186 27806 41188 27858
rect 41132 27794 41188 27806
rect 41244 27300 41300 27310
rect 41020 24697 41022 24749
rect 41074 24697 41076 24749
rect 41020 24685 41076 24697
rect 41132 27074 41188 27086
rect 41132 27022 41134 27074
rect 41186 27022 41188 27074
rect 41020 24052 41076 24062
rect 41020 23958 41076 23996
rect 40908 23847 40910 23899
rect 40962 23847 40964 23899
rect 40908 23835 40964 23847
rect 40460 23548 41076 23604
rect 40460 23268 40516 23278
rect 40460 23154 40516 23212
rect 40460 23102 40462 23154
rect 40514 23102 40516 23154
rect 40460 23090 40516 23102
rect 41020 23154 41076 23548
rect 41020 23102 41022 23154
rect 41074 23102 41076 23154
rect 41020 23090 41076 23102
rect 40292 22932 40348 22942
rect 41132 22932 41188 27022
rect 41244 26317 41300 27244
rect 41692 27300 41748 28590
rect 41916 27746 41972 27758
rect 41916 27694 41918 27746
rect 41970 27694 41972 27746
rect 41916 27300 41972 27694
rect 41916 27244 42084 27300
rect 41692 27234 41748 27244
rect 41916 27076 41972 27086
rect 41244 26265 41246 26317
rect 41298 26265 41300 26317
rect 41244 26253 41300 26265
rect 41468 27074 41972 27076
rect 41468 27022 41918 27074
rect 41970 27022 41972 27074
rect 41468 27020 41972 27022
rect 40292 22930 41188 22932
rect 40292 22878 40294 22930
rect 40346 22878 41188 22930
rect 40292 22876 41188 22878
rect 41244 23938 41300 23950
rect 41244 23886 41246 23938
rect 41298 23886 41300 23938
rect 40292 22866 40348 22876
rect 41244 22820 41300 23886
rect 41356 23169 41412 23194
rect 41356 23156 41358 23169
rect 41410 23156 41412 23169
rect 41356 23090 41412 23100
rect 41468 23042 41524 27020
rect 41916 27010 41972 27020
rect 42028 26908 42084 27244
rect 41916 26852 42084 26908
rect 42140 27076 42196 27086
rect 42140 26908 42196 27020
rect 43036 26908 43092 29922
rect 43372 29652 43428 29662
rect 43372 29558 43428 29596
rect 43596 28868 43652 28878
rect 43596 28756 43652 28812
rect 43596 28754 43764 28756
rect 43596 28702 43598 28754
rect 43650 28702 43764 28754
rect 43596 28700 43764 28702
rect 43596 28690 43652 28700
rect 43484 28644 43540 28654
rect 43484 27188 43540 28588
rect 43708 27524 43764 28700
rect 44212 28420 44268 28430
rect 44212 28418 44436 28420
rect 44212 28366 44214 28418
rect 44266 28366 44436 28418
rect 44212 28364 44436 28366
rect 44212 28354 44268 28364
rect 43820 27748 43876 27758
rect 43820 27746 44212 27748
rect 43820 27694 43822 27746
rect 43874 27694 44212 27746
rect 43820 27692 44212 27694
rect 43820 27682 43876 27692
rect 43708 27468 44100 27524
rect 43484 27132 43988 27188
rect 43708 26964 43764 26974
rect 42140 26852 42308 26908
rect 43036 26852 43204 26908
rect 41692 24948 41748 24958
rect 41692 23910 41748 24892
rect 41692 23858 41694 23910
rect 41746 23858 41748 23910
rect 41692 23846 41748 23858
rect 41916 23492 41972 26852
rect 42252 26514 42308 26852
rect 42252 26462 42254 26514
rect 42306 26462 42308 26514
rect 42252 26450 42308 26462
rect 42943 25450 42999 25462
rect 42700 25396 42756 25406
rect 42700 25302 42756 25340
rect 42943 25398 42945 25450
rect 42997 25398 42999 25450
rect 42364 24948 42420 24958
rect 42364 24854 42420 24892
rect 42943 24836 42999 25398
rect 43148 24948 43204 26852
rect 43708 26178 43764 26908
rect 43820 26962 43876 26974
rect 43820 26910 43822 26962
rect 43874 26910 43876 26962
rect 43820 26628 43876 26910
rect 43820 26562 43876 26572
rect 43932 26404 43988 27132
rect 43876 26348 43988 26404
rect 44044 26404 44100 27468
rect 43876 26346 43932 26348
rect 43876 26294 43878 26346
rect 43930 26294 43932 26346
rect 43876 26282 43932 26294
rect 44044 26346 44100 26348
rect 44044 26294 44046 26346
rect 44098 26294 44100 26346
rect 44044 26282 44100 26294
rect 44156 26180 44212 27692
rect 44380 26908 44436 28364
rect 43708 26126 43710 26178
rect 43762 26126 43764 26178
rect 43708 26114 43764 26126
rect 44044 26124 44212 26180
rect 44268 26852 44436 26908
rect 44268 26292 44324 26852
rect 43820 25508 43876 25518
rect 43820 25414 43876 25452
rect 43148 24892 43652 24948
rect 42943 24780 43316 24836
rect 41916 23426 41972 23436
rect 43036 23268 43092 23278
rect 42159 23156 42215 23166
rect 41468 22990 41470 23042
rect 41522 22990 41524 23042
rect 41468 22978 41524 22990
rect 42140 23154 42215 23156
rect 42140 23102 42161 23154
rect 42213 23102 42215 23154
rect 42140 23090 42215 23102
rect 43036 23154 43092 23212
rect 43036 23102 43038 23154
rect 43090 23102 43092 23154
rect 43036 23090 43092 23102
rect 41916 22930 41972 22942
rect 41916 22878 41918 22930
rect 41970 22878 41972 22930
rect 41916 22820 41972 22878
rect 41244 22764 41972 22820
rect 40572 22708 40628 22718
rect 40460 22372 40516 22382
rect 40124 21298 40180 21308
rect 40348 22370 40516 22372
rect 40348 22318 40462 22370
rect 40514 22318 40516 22370
rect 40348 22316 40516 22318
rect 40124 20804 40180 20814
rect 40124 20468 40180 20748
rect 40124 20402 40180 20412
rect 40348 20244 40404 22316
rect 40460 22306 40516 22316
rect 40236 20188 40404 20244
rect 40460 21586 40516 21598
rect 40460 21534 40462 21586
rect 40514 21534 40516 21586
rect 40460 20244 40516 21534
rect 40572 21476 40628 22652
rect 42140 21700 42196 23090
rect 43036 22820 43092 22830
rect 42252 22708 42308 22718
rect 42252 22260 42308 22652
rect 42924 22596 42980 22606
rect 42924 22502 42980 22540
rect 42364 22260 42420 22270
rect 42252 22258 42420 22260
rect 42252 22206 42366 22258
rect 42418 22206 42420 22258
rect 42252 22204 42420 22206
rect 42364 22194 42420 22204
rect 42140 21634 42196 21644
rect 41132 21588 41188 21598
rect 41132 21494 41188 21532
rect 41916 21476 41972 21486
rect 40572 21420 40684 21476
rect 40628 20858 40684 21420
rect 41916 21474 42196 21476
rect 41916 21422 41918 21474
rect 41970 21422 42196 21474
rect 41916 21420 42196 21422
rect 41916 21410 41972 21420
rect 42140 21028 42196 21420
rect 42252 21028 42308 21038
rect 42140 21026 42308 21028
rect 42140 20974 42254 21026
rect 42306 20974 42308 21026
rect 42140 20972 42308 20974
rect 42252 20962 42308 20972
rect 40628 20806 40630 20858
rect 40682 20806 40684 20858
rect 40628 20794 40684 20806
rect 41300 20804 41356 20814
rect 41300 20710 41356 20748
rect 42588 20804 42644 20814
rect 42906 20804 42962 20814
rect 42588 20802 42962 20804
rect 42588 20750 42590 20802
rect 42642 20750 42908 20802
rect 42960 20750 42962 20802
rect 42588 20748 42962 20750
rect 42588 20738 42644 20748
rect 42906 20738 42962 20748
rect 40796 20692 40852 20702
rect 40796 20598 40852 20636
rect 41860 20578 41916 20590
rect 41860 20526 41862 20578
rect 41914 20526 41916 20578
rect 40460 20188 40964 20244
rect 40236 20130 40292 20188
rect 40236 20078 40238 20130
rect 40290 20078 40292 20130
rect 40236 20066 40292 20078
rect 40796 20018 40852 20030
rect 40796 19966 40798 20018
rect 40850 19966 40852 20018
rect 39770 19366 39826 19404
rect 39900 19404 40068 19460
rect 40124 19908 40180 19918
rect 39452 19236 39508 19246
rect 39340 18452 39396 18462
rect 39340 17666 39396 18396
rect 39452 18450 39508 19180
rect 39452 18398 39454 18450
rect 39506 18398 39508 18450
rect 39452 18386 39508 18398
rect 39788 18452 39844 18462
rect 39788 18358 39844 18396
rect 39340 17614 39342 17666
rect 39394 17614 39396 17666
rect 39340 17602 39396 17614
rect 39788 17220 39844 17230
rect 39116 16818 39172 16828
rect 39676 16884 39732 16894
rect 39788 16884 39844 17164
rect 39676 16882 39844 16884
rect 39676 16830 39678 16882
rect 39730 16830 39790 16882
rect 39842 16830 39844 16882
rect 39676 16828 39844 16830
rect 39676 16818 39732 16828
rect 39340 16658 39396 16670
rect 39340 16606 39342 16658
rect 39394 16606 39396 16658
rect 37660 16324 37716 16334
rect 37100 16322 37716 16324
rect 37100 16270 37662 16322
rect 37714 16270 37716 16322
rect 37100 16268 37716 16270
rect 36540 15876 36596 15886
rect 36372 15540 36428 15550
rect 36372 15204 36428 15484
rect 36372 15138 36428 15148
rect 36540 15148 36596 15820
rect 36764 15316 36820 15326
rect 36764 15222 36820 15260
rect 37100 15314 37156 16268
rect 37660 16258 37716 16268
rect 38444 16212 38500 16222
rect 37324 16098 37380 16110
rect 37324 16046 37326 16098
rect 37378 16046 37380 16098
rect 37100 15262 37102 15314
rect 37154 15262 37156 15314
rect 36540 15092 36708 15148
rect 36372 14532 36428 14542
rect 36372 14438 36428 14476
rect 36204 12908 36372 12964
rect 35084 12180 35140 12190
rect 35084 12086 35140 12124
rect 33964 11396 34020 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35532 11620 35588 12674
rect 35420 11564 35588 11620
rect 35644 12292 35700 12302
rect 34300 11508 34356 11518
rect 33964 11340 34132 11396
rect 33944 11172 34000 11182
rect 33944 10666 34000 11116
rect 33944 10614 33946 10666
rect 33998 10614 34000 10666
rect 33944 10602 34000 10614
rect 34076 9044 34132 11340
rect 34188 10612 34244 10622
rect 34188 10518 34244 10556
rect 34076 8988 34244 9044
rect 34076 8820 34132 8830
rect 33740 8316 34020 8372
rect 33964 6804 34020 8316
rect 34076 8370 34132 8764
rect 34076 8318 34078 8370
rect 34130 8318 34132 8370
rect 34076 8306 34132 8318
rect 32956 5070 32958 5122
rect 33010 5070 33012 5122
rect 32956 5058 33012 5070
rect 33628 6748 34020 6804
rect 32284 3726 32286 3778
rect 32338 3726 32340 3778
rect 32284 3714 32340 3726
rect 33404 4338 33460 4350
rect 33404 4286 33406 4338
rect 33458 4286 33460 4338
rect 33404 3778 33460 4286
rect 33628 4340 33684 6748
rect 33964 6692 34020 6748
rect 34188 7476 34244 8988
rect 34300 9042 34356 11452
rect 34524 11508 34580 11518
rect 34524 11506 34916 11508
rect 34524 11454 34526 11506
rect 34578 11454 34916 11506
rect 34524 11452 34916 11454
rect 34524 11442 34580 11452
rect 34860 11396 34916 11452
rect 34300 8990 34302 9042
rect 34354 8990 34356 9042
rect 34300 8978 34356 8990
rect 34412 10724 34468 10734
rect 34412 9938 34468 10668
rect 34636 10724 34692 10734
rect 34860 10724 34916 11340
rect 34860 10668 34972 10724
rect 34636 10610 34692 10668
rect 34636 10558 34638 10610
rect 34690 10558 34692 10610
rect 34916 10666 34972 10668
rect 34916 10614 34918 10666
rect 34970 10614 34972 10666
rect 34916 10602 34972 10614
rect 35420 10610 35476 11564
rect 34636 10546 34692 10558
rect 35420 10558 35422 10610
rect 35474 10558 35476 10610
rect 35420 10546 35476 10558
rect 35532 11366 35588 11378
rect 35532 11314 35534 11366
rect 35586 11314 35588 11366
rect 35084 10498 35140 10510
rect 35084 10446 35086 10498
rect 35138 10446 35140 10498
rect 35084 10388 35140 10446
rect 35084 10322 35140 10332
rect 35532 10276 35588 11314
rect 35644 10500 35700 12236
rect 35756 10836 35812 12684
rect 35980 11788 36036 12908
rect 36148 12740 36204 12778
rect 36148 12674 36204 12684
rect 36092 12516 36148 12526
rect 36092 12178 36148 12460
rect 36092 12126 36094 12178
rect 36146 12126 36148 12178
rect 36092 12114 36148 12126
rect 36316 12180 36372 12908
rect 36428 12404 36484 12414
rect 36428 12310 36484 12348
rect 36316 12124 36484 12180
rect 35980 11732 36260 11788
rect 35868 11508 35924 11518
rect 35868 11414 35924 11452
rect 35980 11396 36036 11406
rect 35980 11327 35982 11340
rect 36034 11327 36036 11340
rect 35980 11302 36036 11327
rect 36204 11396 36260 11732
rect 36204 11302 36260 11340
rect 35756 10780 36148 10836
rect 35644 10434 35700 10444
rect 35196 10220 35460 10230
rect 35532 10220 35924 10276
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34412 9886 34414 9938
rect 34466 9886 34468 9938
rect 34412 8484 34468 9886
rect 35196 9828 35252 9838
rect 35196 9734 35252 9772
rect 35532 9492 35588 9502
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34300 8428 34468 8484
rect 34300 7924 34356 8428
rect 35532 8270 35588 9436
rect 35868 9268 35924 10220
rect 36092 9782 36148 10780
rect 36072 9770 36148 9782
rect 36072 9718 36074 9770
rect 36126 9718 36148 9770
rect 36072 9660 36148 9718
rect 36204 10498 36260 10510
rect 36204 10446 36206 10498
rect 36258 10446 36260 10498
rect 35868 9202 35924 9212
rect 36204 9156 36260 10446
rect 36428 10276 36484 12124
rect 36652 10836 36708 15092
rect 36876 15092 36932 15102
rect 36876 13746 36932 15036
rect 37100 14756 37156 15262
rect 37212 15316 37268 15326
rect 37212 15222 37268 15260
rect 37100 14690 37156 14700
rect 37156 14474 37212 14486
rect 36988 14420 37044 14430
rect 36988 14326 37044 14364
rect 37156 14422 37158 14474
rect 37210 14422 37212 14474
rect 37156 13860 37212 14422
rect 37324 13972 37380 16046
rect 38444 16098 38500 16156
rect 39340 16212 39396 16606
rect 39340 16146 39396 16156
rect 38444 16046 38446 16098
rect 38498 16046 38500 16098
rect 38444 16034 38500 16046
rect 38948 16042 39004 16054
rect 38202 15988 38258 15998
rect 38948 15990 38950 16042
rect 39002 15990 39004 16042
rect 39788 15998 39844 16828
rect 39900 16212 39956 19404
rect 40012 19234 40068 19246
rect 40012 19182 40014 19234
rect 40066 19182 40068 19234
rect 40012 17668 40068 19182
rect 40124 18450 40180 19852
rect 40124 18398 40126 18450
rect 40178 18398 40180 18450
rect 40124 18386 40180 18398
rect 40236 19796 40292 19806
rect 40124 17780 40180 17790
rect 40236 17780 40292 19740
rect 40796 19460 40852 19966
rect 40796 19394 40852 19404
rect 40516 19348 40572 19358
rect 40516 19290 40572 19292
rect 40516 19238 40518 19290
rect 40570 19238 40572 19290
rect 40516 19226 40572 19238
rect 40908 19236 40964 20188
rect 41692 20020 41748 20030
rect 41468 20018 41748 20020
rect 41468 19966 41694 20018
rect 41746 19966 41748 20018
rect 41468 19964 41748 19966
rect 41132 19796 41188 19806
rect 41132 19702 41188 19740
rect 40908 19142 40964 19180
rect 40684 19124 40740 19134
rect 40684 18116 40740 19068
rect 40796 18452 40852 18462
rect 40796 18358 40852 18396
rect 40684 18050 40740 18060
rect 40124 17778 40292 17780
rect 40124 17726 40126 17778
rect 40178 17726 40292 17778
rect 40124 17724 40292 17726
rect 40124 17714 40180 17724
rect 40012 17108 40068 17612
rect 41076 17220 41132 17230
rect 40124 17108 40180 17118
rect 40012 17106 40180 17108
rect 40012 17054 40126 17106
rect 40178 17054 40180 17106
rect 40012 17052 40180 17054
rect 40124 17042 40180 17052
rect 41076 17106 41132 17164
rect 41076 17054 41078 17106
rect 41130 17054 41132 17106
rect 41076 17042 41132 17054
rect 41468 17006 41524 19964
rect 41692 19954 41748 19964
rect 41860 20020 41916 20526
rect 41860 19954 41916 19964
rect 42924 20020 42980 20030
rect 43036 20020 43092 22764
rect 43260 22484 43316 24780
rect 43372 23716 43428 23726
rect 43372 23714 43540 23716
rect 43372 23662 43374 23714
rect 43426 23662 43540 23714
rect 43372 23660 43540 23662
rect 43372 23650 43428 23660
rect 43372 23492 43428 23502
rect 43372 23042 43428 23436
rect 43484 23198 43540 23660
rect 43484 23156 43486 23198
rect 43538 23156 43540 23198
rect 43484 23068 43540 23100
rect 43372 22990 43374 23042
rect 43426 22990 43428 23042
rect 43372 22978 43428 22990
rect 43596 22820 43652 24892
rect 43932 24500 43988 24510
rect 43932 24406 43988 24444
rect 44044 24052 44100 26124
rect 44156 25956 44212 25966
rect 44156 24500 44212 25900
rect 44268 24722 44324 26236
rect 44380 26628 44436 26638
rect 44380 25508 44436 26572
rect 44380 25442 44436 25452
rect 44268 24670 44270 24722
rect 44322 24670 44324 24722
rect 44268 24658 44324 24670
rect 44380 24724 44436 24734
rect 44156 24444 44324 24500
rect 43820 23996 44100 24052
rect 43820 23268 43876 23996
rect 43820 23154 43876 23212
rect 43820 23102 43822 23154
rect 43874 23102 43876 23154
rect 43820 23090 43876 23102
rect 43596 22754 43652 22764
rect 43260 22428 43428 22484
rect 43167 22314 43223 22326
rect 43167 22262 43169 22314
rect 43221 22262 43223 22314
rect 43167 22260 43223 22262
rect 43167 22204 43316 22260
rect 43148 20804 43204 20814
rect 43148 20710 43204 20748
rect 43260 20132 43316 22204
rect 42924 20018 43092 20020
rect 42924 19966 42926 20018
rect 42978 19966 43038 20018
rect 43090 19966 43092 20018
rect 42924 19964 43092 19966
rect 42924 19954 42980 19964
rect 42028 19796 42084 19806
rect 41580 19794 42084 19796
rect 41580 19742 42030 19794
rect 42082 19742 42084 19794
rect 41580 19740 42084 19742
rect 41580 18450 41636 19740
rect 42028 19730 42084 19740
rect 42588 19794 42644 19806
rect 42588 19742 42590 19794
rect 42642 19742 42644 19794
rect 42588 19572 42644 19742
rect 42588 19516 42980 19572
rect 41804 19348 41860 19358
rect 41580 18398 41582 18450
rect 41634 18398 41636 18450
rect 41580 18386 41636 18398
rect 41692 19234 41748 19246
rect 41692 19182 41694 19234
rect 41746 19182 41748 19234
rect 41692 17108 41748 19182
rect 41804 18116 41860 19292
rect 42700 18676 42756 18686
rect 41804 18060 42084 18116
rect 42028 17778 42084 18060
rect 42700 17780 42756 18620
rect 42028 17726 42030 17778
rect 42082 17726 42084 17778
rect 42028 17714 42084 17726
rect 42252 17724 42756 17780
rect 42812 18340 42868 18350
rect 42812 17780 42868 18284
rect 42252 17556 42308 17724
rect 42812 17666 42868 17724
rect 42812 17614 42814 17666
rect 42866 17614 42868 17666
rect 42812 17602 42868 17614
rect 41692 17042 41748 17052
rect 42196 17500 42308 17556
rect 42570 17556 42626 17566
rect 42570 17554 42644 17556
rect 42570 17502 42572 17554
rect 42624 17502 42644 17554
rect 41450 16994 41524 17006
rect 41450 16942 41452 16994
rect 41504 16942 41524 16994
rect 41450 16940 41524 16942
rect 41450 16930 41506 16940
rect 42196 16938 42252 17500
rect 42570 17490 42644 17502
rect 41692 16884 41748 16894
rect 42196 16886 42198 16938
rect 42250 16886 42252 16938
rect 42364 16996 42420 17006
rect 42364 16902 42420 16940
rect 42196 16874 42252 16886
rect 42588 16882 42644 17490
rect 42924 17444 42980 19516
rect 43036 18452 43092 19964
rect 43148 20076 43316 20132
rect 43148 19348 43204 20076
rect 43372 20020 43428 22428
rect 44044 22372 44100 22382
rect 44268 22372 44324 24444
rect 44044 22370 44324 22372
rect 44044 22318 44046 22370
rect 44098 22318 44324 22370
rect 44044 22316 44324 22318
rect 44044 22306 44100 22316
rect 44380 22036 44436 24668
rect 43820 21980 44436 22036
rect 44492 24500 44548 24510
rect 43148 19282 43204 19292
rect 43260 19964 43428 20020
rect 43484 21700 43540 21710
rect 43820 21700 43876 21980
rect 43036 18386 43092 18396
rect 43148 19124 43204 19134
rect 41692 16790 41748 16828
rect 42588 16830 42590 16882
rect 42642 16830 42644 16882
rect 42588 16818 42644 16830
rect 42812 17388 42980 17444
rect 43148 17498 43204 19068
rect 43260 18676 43316 19964
rect 43372 19796 43428 19806
rect 43372 19702 43428 19740
rect 43484 19348 43540 21644
rect 43708 21698 43876 21700
rect 43708 21646 43822 21698
rect 43874 21646 43876 21698
rect 43708 21644 43876 21646
rect 43708 21476 43764 21644
rect 43820 21634 43876 21644
rect 43652 21420 43764 21476
rect 43652 20858 43708 21420
rect 43652 20806 43654 20858
rect 43706 20806 43708 20858
rect 43652 20794 43708 20806
rect 44268 20804 44324 20814
rect 43596 20634 43652 20646
rect 43596 20582 43598 20634
rect 43650 20582 43652 20634
rect 43596 19684 43652 20582
rect 43596 19618 43652 19628
rect 43708 20020 43764 20030
rect 43708 19572 43764 19964
rect 43708 19506 43764 19516
rect 44044 19908 44100 19918
rect 43596 19348 43652 19358
rect 43260 18610 43316 18620
rect 43372 19346 43652 19348
rect 43372 19294 43598 19346
rect 43650 19294 43652 19346
rect 43372 19292 43652 19294
rect 43372 18228 43428 19292
rect 43596 19282 43652 19292
rect 43484 18676 43540 18686
rect 43484 18450 43540 18620
rect 43484 18398 43486 18450
rect 43538 18398 43540 18450
rect 43484 18386 43540 18398
rect 43596 18452 43652 18462
rect 43316 18172 43428 18228
rect 43316 17722 43372 18172
rect 43316 17670 43318 17722
rect 43370 17670 43372 17722
rect 43316 17658 43372 17670
rect 43148 17446 43150 17498
rect 43202 17446 43204 17498
rect 42812 16884 42868 17388
rect 42924 17108 42980 17118
rect 42924 17014 42980 17052
rect 43148 16996 43204 17446
rect 43596 17118 43652 18396
rect 43540 17106 43652 17118
rect 43540 17054 43542 17106
rect 43594 17054 43652 17106
rect 43540 17052 43652 17054
rect 43820 18340 43876 18350
rect 43820 17220 43876 18284
rect 43932 17780 43988 17790
rect 43932 17686 43988 17724
rect 43820 17108 43876 17164
rect 43932 17108 43988 17118
rect 43820 17106 43988 17108
rect 43820 17054 43934 17106
rect 43986 17054 43988 17106
rect 43820 17052 43988 17054
rect 43540 17042 43596 17052
rect 43932 17042 43988 17052
rect 43148 16930 43204 16940
rect 42812 16818 42868 16828
rect 43540 16324 43596 16334
rect 39900 16146 39956 16156
rect 40292 16212 40348 16222
rect 40292 16118 40348 16156
rect 43540 16210 43596 16268
rect 43540 16158 43542 16210
rect 43594 16158 43596 16210
rect 43540 16146 43596 16158
rect 38202 15986 38276 15988
rect 38202 15934 38204 15986
rect 38256 15934 38276 15986
rect 38202 15922 38276 15934
rect 37324 13906 37380 13916
rect 37660 15204 37716 15214
rect 37660 14530 37716 15148
rect 37996 15202 38052 15214
rect 37996 15150 37998 15202
rect 38050 15150 38052 15202
rect 37660 14478 37662 14530
rect 37714 14478 37716 14530
rect 37660 13972 37716 14478
rect 37772 14756 37828 14766
rect 37772 14196 37828 14700
rect 37996 14756 38052 15150
rect 37996 14690 38052 14700
rect 38220 14532 38276 15922
rect 38948 15540 39004 15990
rect 39116 15988 39172 15998
rect 39788 15986 39900 15998
rect 39788 15934 39846 15986
rect 39898 15934 39900 15986
rect 39788 15932 39900 15934
rect 39116 15894 39172 15932
rect 39844 15922 39900 15932
rect 41468 15988 41524 15998
rect 38948 15484 39956 15540
rect 39900 15426 39956 15484
rect 39900 15374 39902 15426
rect 39954 15374 39956 15426
rect 39900 15148 39956 15374
rect 41468 15426 41524 15932
rect 41468 15374 41470 15426
rect 41522 15374 41524 15426
rect 40796 15316 40852 15326
rect 39900 15092 40068 15148
rect 38780 14756 38836 14766
rect 38780 14662 38836 14700
rect 38444 14532 38500 14542
rect 38220 14530 38500 14532
rect 38220 14478 38446 14530
rect 38498 14478 38500 14530
rect 38220 14476 38500 14478
rect 38444 14466 38500 14476
rect 37902 14420 37958 14430
rect 37902 14326 37958 14364
rect 39116 14420 39172 14430
rect 37772 14140 38052 14196
rect 37660 13906 37716 13916
rect 36876 13694 36878 13746
rect 36930 13694 36932 13746
rect 36876 13682 36932 13694
rect 37100 13804 37212 13860
rect 37100 12852 37156 13804
rect 37996 13412 38052 14140
rect 39116 13746 39172 14364
rect 39116 13694 39118 13746
rect 39170 13694 39172 13746
rect 39116 13682 39172 13694
rect 38780 13636 38836 13646
rect 38780 13542 38836 13580
rect 39452 13524 39508 13534
rect 37100 12758 37156 12796
rect 37884 13356 38052 13412
rect 39004 13522 39508 13524
rect 39004 13470 39454 13522
rect 39506 13470 39508 13522
rect 39004 13468 39508 13470
rect 37324 12205 37380 12217
rect 37324 12180 37326 12205
rect 37378 12180 37380 12205
rect 37324 12113 37380 12124
rect 37772 12180 37828 12190
rect 37884 12180 37940 13356
rect 39004 13074 39060 13468
rect 39452 13458 39508 13468
rect 39004 13022 39006 13074
rect 39058 13022 39060 13074
rect 39004 13010 39060 13022
rect 39788 12964 39844 12974
rect 39788 12870 39844 12908
rect 37828 12124 37940 12180
rect 38892 12852 38948 12862
rect 37212 11394 37268 11406
rect 37212 11342 37214 11394
rect 37266 11342 37268 11394
rect 37212 11284 37268 11342
rect 37212 11218 37268 11228
rect 36652 10770 36708 10780
rect 36428 10220 36820 10276
rect 36316 10052 36372 10062
rect 36316 9958 36372 9996
rect 36540 10052 36596 10062
rect 34636 8258 34692 8270
rect 34412 8202 34468 8214
rect 34412 8150 34414 8202
rect 34466 8150 34468 8202
rect 34412 8148 34468 8150
rect 34412 8082 34468 8092
rect 34636 8206 34638 8258
rect 34690 8206 34692 8258
rect 34636 7924 34692 8206
rect 35512 8258 35588 8270
rect 35512 8206 35514 8258
rect 35566 8206 35588 8258
rect 35512 8204 35588 8206
rect 35980 9100 36260 9156
rect 35512 8194 35568 8204
rect 35756 8148 35812 8158
rect 34300 7868 34692 7924
rect 35644 8146 35812 8148
rect 35644 8094 35758 8146
rect 35810 8094 35812 8146
rect 35644 8092 35812 8094
rect 34076 6692 34132 6702
rect 33964 6690 34132 6692
rect 33964 6638 34078 6690
rect 34130 6638 34132 6690
rect 33964 6636 34132 6638
rect 34076 6626 34132 6636
rect 33834 6580 33890 6590
rect 33834 6578 34020 6580
rect 33834 6526 33836 6578
rect 33888 6526 34020 6578
rect 33834 6524 34020 6526
rect 33834 6514 33890 6524
rect 33740 6132 33796 6142
rect 33964 6132 34020 6524
rect 33964 6076 34132 6132
rect 33740 6018 33796 6076
rect 33740 5966 33742 6018
rect 33794 5966 33796 6018
rect 33740 5954 33796 5966
rect 33908 5908 33964 5918
rect 33908 5814 33964 5852
rect 34076 5460 34132 6076
rect 34188 5908 34244 7420
rect 35420 7252 35476 7262
rect 35420 7250 35588 7252
rect 35420 7198 35422 7250
rect 35474 7198 35588 7250
rect 35420 7196 35588 7198
rect 35420 7186 35476 7196
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35420 6692 35476 6702
rect 34580 6634 34636 6646
rect 34580 6582 34582 6634
rect 34634 6582 34636 6634
rect 35252 6634 35308 6646
rect 34580 6132 34636 6582
rect 34748 6580 34804 6590
rect 35084 6580 35140 6590
rect 34748 6578 35140 6580
rect 34748 6526 34750 6578
rect 34802 6526 35086 6578
rect 35138 6526 35140 6578
rect 34748 6524 35140 6526
rect 34748 6356 34804 6524
rect 35084 6514 35140 6524
rect 35252 6582 35254 6634
rect 35306 6582 35308 6634
rect 34748 6290 34804 6300
rect 35252 6244 35308 6582
rect 35252 6178 35308 6188
rect 34580 6076 34916 6132
rect 34412 5908 34468 5918
rect 34188 5906 34468 5908
rect 34188 5854 34414 5906
rect 34466 5854 34468 5906
rect 34188 5852 34468 5854
rect 34412 5842 34468 5852
rect 34654 5684 34710 5694
rect 34654 5590 34710 5628
rect 33964 5404 34132 5460
rect 33740 5124 33796 5134
rect 33740 5030 33796 5068
rect 33628 4274 33684 4284
rect 33964 4004 34020 5404
rect 34860 4564 34916 6076
rect 35420 6018 35476 6636
rect 35420 5966 35422 6018
rect 35474 5966 35476 6018
rect 35420 5954 35476 5966
rect 35532 6020 35588 7196
rect 35644 6580 35700 8092
rect 35756 8082 35812 8092
rect 35756 7476 35812 7486
rect 35756 7382 35812 7420
rect 35980 7362 36036 9100
rect 36204 8932 36260 8942
rect 36204 8838 36260 8876
rect 36540 8596 36596 9996
rect 36652 9069 36708 9081
rect 36652 9017 36654 9069
rect 36706 9017 36708 9069
rect 36652 8820 36708 9017
rect 36652 8754 36708 8764
rect 36372 8540 36596 8596
rect 36372 8372 36428 8540
rect 36204 8370 36428 8372
rect 36204 8318 36374 8370
rect 36426 8318 36428 8370
rect 36204 8316 36428 8318
rect 36092 8036 36148 8046
rect 36092 7518 36148 7980
rect 36092 7466 36094 7518
rect 36146 7466 36148 7518
rect 36092 7454 36148 7466
rect 35980 7310 35982 7362
rect 36034 7310 36036 7362
rect 35980 7298 36036 7310
rect 36204 7140 36260 8316
rect 36372 8306 36428 8316
rect 36540 8372 36596 8382
rect 36428 7476 36484 7486
rect 36540 7476 36596 8316
rect 36428 7474 36596 7476
rect 36428 7422 36430 7474
rect 36482 7422 36596 7474
rect 36428 7420 36596 7422
rect 36428 7410 36484 7420
rect 35644 6514 35700 6524
rect 35756 7084 36260 7140
rect 35756 6690 35812 7084
rect 35756 6638 35758 6690
rect 35810 6638 35812 6690
rect 35756 6468 35812 6638
rect 35998 6580 36054 6590
rect 35756 6402 35812 6412
rect 35868 6578 36054 6580
rect 35868 6526 36000 6578
rect 36052 6526 36054 6578
rect 35868 6524 36054 6526
rect 35532 5954 35588 5964
rect 35663 5908 35719 5946
rect 35644 5852 35663 5908
rect 35644 5842 35719 5852
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35644 5234 35700 5842
rect 35868 5796 35924 6524
rect 35998 6514 36054 6524
rect 36540 6132 36596 6142
rect 36540 5906 36596 6076
rect 36540 5854 36542 5906
rect 36594 5854 36596 5906
rect 36540 5842 36596 5854
rect 35644 5182 35646 5234
rect 35698 5182 35700 5234
rect 35644 5170 35700 5182
rect 35756 5740 35924 5796
rect 35756 4900 35812 5740
rect 35868 5572 35924 5582
rect 35868 5124 35924 5516
rect 35980 5124 36036 5134
rect 35868 5122 36036 5124
rect 35868 5070 35982 5122
rect 36034 5070 36036 5122
rect 35868 5068 36036 5070
rect 35980 5058 36036 5068
rect 36316 5124 36372 5134
rect 36316 5030 36372 5068
rect 36652 5124 36708 5134
rect 35756 4844 36484 4900
rect 34860 4498 34916 4508
rect 36092 4564 36148 4574
rect 36092 4450 36148 4508
rect 36092 4398 36094 4450
rect 36146 4398 36148 4450
rect 36092 4386 36148 4398
rect 34188 4228 34244 4238
rect 34188 4226 34468 4228
rect 34188 4174 34190 4226
rect 34242 4174 34468 4226
rect 34188 4172 34468 4174
rect 34188 4162 34244 4172
rect 33964 3948 34356 4004
rect 33404 3726 33406 3778
rect 33458 3726 33460 3778
rect 33404 3714 33460 3726
rect 28252 3500 28420 3502
rect 24556 3474 24558 3500
rect 24610 3474 24612 3500
rect 28364 3490 28420 3500
rect 29036 3502 29038 3554
rect 29090 3502 29092 3554
rect 29036 3490 29092 3502
rect 34300 3554 34356 3948
rect 34412 3780 34468 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34636 3780 34692 3790
rect 34412 3778 34692 3780
rect 34412 3726 34638 3778
rect 34690 3726 34692 3778
rect 34412 3724 34692 3726
rect 34636 3714 34692 3724
rect 34300 3502 34302 3554
rect 34354 3502 34356 3554
rect 34300 3490 34356 3502
rect 36428 3554 36484 4844
rect 36652 3780 36708 5068
rect 36764 4900 36820 10220
rect 36876 9826 36932 9838
rect 37660 9828 37716 9838
rect 36876 9774 36878 9826
rect 36930 9774 36932 9826
rect 36876 8036 36932 9774
rect 37436 9826 37716 9828
rect 37436 9774 37662 9826
rect 37714 9774 37716 9826
rect 37436 9772 37716 9774
rect 37324 9044 37380 9054
rect 37212 8372 37268 8382
rect 37212 8258 37268 8316
rect 37212 8206 37214 8258
rect 37266 8206 37268 8258
rect 37212 8194 37268 8206
rect 37044 8036 37100 8046
rect 36876 8034 37100 8036
rect 36876 7982 37046 8034
rect 37098 7982 37100 8034
rect 36876 7980 37100 7982
rect 37044 7970 37100 7980
rect 37212 8036 37268 8046
rect 36988 7812 37044 7822
rect 36876 7588 36932 7598
rect 36876 5122 36932 7532
rect 36988 7474 37044 7756
rect 36988 7422 36990 7474
rect 37042 7422 37044 7474
rect 36988 7410 37044 7422
rect 37100 7700 37156 7710
rect 37100 6802 37156 7644
rect 37100 6750 37102 6802
rect 37154 6750 37156 6802
rect 37100 6738 37156 6750
rect 36988 6692 37044 6702
rect 36988 6598 37044 6636
rect 37212 6580 37268 7980
rect 37324 7700 37380 8988
rect 37324 7634 37380 7644
rect 37324 7474 37380 7486
rect 37324 7422 37326 7474
rect 37378 7422 37380 7474
rect 37324 6804 37380 7422
rect 37324 6738 37380 6748
rect 37100 6524 37268 6580
rect 37324 6634 37380 6646
rect 37324 6582 37326 6634
rect 37378 6582 37380 6634
rect 37100 5950 37156 6524
rect 37324 6468 37380 6582
rect 37100 5898 37102 5950
rect 37154 5898 37156 5950
rect 37100 5886 37156 5898
rect 37212 6412 37380 6468
rect 37212 5460 37268 6412
rect 37436 6356 37492 9772
rect 37660 9762 37716 9772
rect 37548 8260 37604 8270
rect 37548 8178 37550 8204
rect 37602 8178 37604 8204
rect 37548 8166 37604 8178
rect 37772 7700 37828 12124
rect 38780 10612 38836 10622
rect 38780 10518 38836 10556
rect 38108 10500 38164 10510
rect 37884 10498 38164 10500
rect 37884 10446 38110 10498
rect 38162 10446 38164 10498
rect 37884 10444 38164 10446
rect 37884 8372 37940 10444
rect 38108 10434 38164 10444
rect 37996 9268 38052 9278
rect 37996 9174 38052 9212
rect 37884 7924 37940 8316
rect 38892 8148 38948 12796
rect 38687 8092 38948 8148
rect 39004 11954 39060 11966
rect 39004 11902 39006 11954
rect 39058 11902 39060 11954
rect 39004 8148 39060 11902
rect 39900 11508 39956 11518
rect 39116 11506 39956 11508
rect 39116 11454 39902 11506
rect 39954 11454 39956 11506
rect 39116 11452 39956 11454
rect 39116 10610 39172 11452
rect 39900 11442 39956 11452
rect 40012 11396 40068 15092
rect 40796 14532 40852 15260
rect 40572 14530 40852 14532
rect 40572 14478 40798 14530
rect 40850 14478 40852 14530
rect 40572 14476 40852 14478
rect 40460 13748 40516 13758
rect 40460 13654 40516 13692
rect 40124 13522 40180 13534
rect 40124 13470 40126 13522
rect 40178 13470 40180 13522
rect 40124 13076 40180 13470
rect 40124 13010 40180 13020
rect 40572 12964 40628 14476
rect 40796 14466 40852 14476
rect 41188 13972 41244 13982
rect 41188 13878 41244 13916
rect 41468 13860 41524 15374
rect 43652 15540 43708 15550
rect 41636 15316 41692 15326
rect 41636 15314 41860 15316
rect 41636 15262 41638 15314
rect 41690 15262 41860 15314
rect 41636 15260 41860 15262
rect 41636 15250 41692 15260
rect 41580 15092 41636 15102
rect 41580 14642 41636 15036
rect 41580 14590 41582 14642
rect 41634 14590 41636 14642
rect 41580 14578 41636 14590
rect 41468 13766 41524 13804
rect 41636 14196 41692 14206
rect 41636 13690 41692 14140
rect 41636 13638 41638 13690
rect 41690 13638 41692 13690
rect 41636 13300 41692 13638
rect 41804 13524 41860 15260
rect 42140 15314 42196 15326
rect 42140 15262 42142 15314
rect 42194 15262 42196 15314
rect 42140 14868 42196 15262
rect 42700 15314 42756 15326
rect 42700 15262 42702 15314
rect 42754 15262 42756 15314
rect 42382 15092 42438 15102
rect 42382 14998 42438 15036
rect 42140 14802 42196 14812
rect 42140 14308 42196 14318
rect 42700 14308 42756 15262
rect 43036 15204 43092 15242
rect 43652 15148 43708 15484
rect 43036 15138 43092 15148
rect 42140 13746 42196 14252
rect 42382 14252 42756 14308
rect 43372 15092 43428 15102
rect 42382 13858 42438 14252
rect 42382 13806 42384 13858
rect 42436 13806 42438 13858
rect 42382 13794 42438 13806
rect 43148 13972 43204 13982
rect 42140 13694 42142 13746
rect 42194 13694 42196 13746
rect 42140 13682 42196 13694
rect 42906 13748 42962 13758
rect 42906 13654 42962 13692
rect 43148 13746 43204 13916
rect 43148 13694 43150 13746
rect 43202 13694 43204 13746
rect 43148 13682 43204 13694
rect 41804 13458 41860 13468
rect 41580 13244 41692 13300
rect 43260 13412 43316 13422
rect 41356 13076 41412 13086
rect 41356 12982 41412 13020
rect 40572 12870 40628 12908
rect 40908 12180 40964 12190
rect 40908 12086 40964 12124
rect 40143 11396 40199 11406
rect 40012 11394 40199 11396
rect 39116 10558 39118 10610
rect 39170 10558 39172 10610
rect 39116 10546 39172 10558
rect 39228 11366 39284 11378
rect 39228 11314 39230 11366
rect 39282 11314 39284 11366
rect 40012 11342 40145 11394
rect 40197 11342 40199 11394
rect 40012 11340 40199 11342
rect 40143 11330 40199 11340
rect 41020 11394 41076 11406
rect 41020 11342 41022 11394
rect 41074 11342 41076 11394
rect 39228 8260 39284 11314
rect 39788 11284 39844 11294
rect 39452 10724 39508 10734
rect 39340 10649 39396 10661
rect 39340 10597 39342 10649
rect 39394 10597 39396 10649
rect 39340 10276 39396 10597
rect 39340 10210 39396 10220
rect 39452 9940 39508 10668
rect 39676 10612 39732 10622
rect 39676 10518 39732 10556
rect 39564 10498 39620 10510
rect 39564 10446 39566 10498
rect 39618 10446 39620 10498
rect 39564 10052 39620 10446
rect 39788 10388 39844 11228
rect 40012 10724 40068 10734
rect 40012 10610 40068 10668
rect 41020 10724 41076 11342
rect 41468 11284 41524 11294
rect 41468 11190 41524 11228
rect 41580 11172 41636 13244
rect 43260 12850 43316 13356
rect 43372 12964 43428 15036
rect 43596 15092 43708 15148
rect 44044 15148 44100 19852
rect 44268 19358 44324 20748
rect 44492 20804 44548 24444
rect 44492 20738 44548 20748
rect 44212 19346 44324 19358
rect 44212 19294 44214 19346
rect 44266 19294 44324 19346
rect 44212 19292 44324 19294
rect 44380 19572 44436 19582
rect 44212 19282 44268 19292
rect 44212 18452 44268 18462
rect 44212 18358 44268 18396
rect 44268 17668 44324 17678
rect 44380 17668 44436 19516
rect 44268 17666 44436 17668
rect 44268 17614 44270 17666
rect 44322 17614 44436 17666
rect 44268 17612 44436 17614
rect 44268 17602 44324 17612
rect 44268 16882 44324 16894
rect 44268 16830 44270 16882
rect 44322 16830 44324 16882
rect 44268 16222 44324 16830
rect 44380 16324 44436 17612
rect 44380 16258 44436 16268
rect 44212 16212 44324 16222
rect 44268 16156 44324 16212
rect 44212 16118 44268 16156
rect 44044 15092 44156 15148
rect 43596 14868 43652 15092
rect 43596 14802 43652 14812
rect 43484 14418 43540 14430
rect 43484 14366 43486 14418
rect 43538 14366 43540 14418
rect 43484 14196 43540 14366
rect 44100 14308 44156 15092
rect 44100 14214 44156 14252
rect 43484 14130 43540 14140
rect 43484 13914 43540 13926
rect 43484 13862 43486 13914
rect 43538 13862 43540 13914
rect 43484 13860 43540 13862
rect 43484 13794 43540 13804
rect 43652 13690 43708 13702
rect 43652 13638 43654 13690
rect 43706 13638 43708 13690
rect 43484 13524 43540 13534
rect 43484 13188 43540 13468
rect 43652 13412 43708 13638
rect 43652 13346 43708 13356
rect 43484 13132 43764 13188
rect 43596 12964 43652 12974
rect 43372 12962 43652 12964
rect 43372 12910 43598 12962
rect 43650 12910 43652 12962
rect 43372 12908 43652 12910
rect 43596 12898 43652 12908
rect 43260 12798 43262 12850
rect 43314 12798 43316 12850
rect 41692 12180 41748 12190
rect 41692 12086 41748 12124
rect 41711 11844 41767 11854
rect 41711 11394 41767 11788
rect 43260 11844 43316 12798
rect 43708 12740 43764 13132
rect 44380 12852 44436 12862
rect 43596 12684 43764 12740
rect 43932 12738 43988 12750
rect 43932 12686 43934 12738
rect 43986 12686 43988 12738
rect 43596 12292 43652 12684
rect 43260 11778 43316 11788
rect 43372 12290 43652 12292
rect 43372 12238 43598 12290
rect 43650 12238 43652 12290
rect 43372 12236 43652 12238
rect 41711 11342 41713 11394
rect 41765 11342 41767 11394
rect 41711 11330 41767 11342
rect 42588 11396 42644 11406
rect 42812 11396 42868 11406
rect 43372 11396 43428 12236
rect 43596 12226 43652 12236
rect 43932 12180 43988 12686
rect 43932 12114 43988 12124
rect 44212 12068 44268 12078
rect 44156 12066 44268 12068
rect 44156 12014 44214 12066
rect 44266 12014 44268 12066
rect 44156 12002 44268 12014
rect 43932 11620 43988 11630
rect 43932 11526 43988 11564
rect 42588 11394 42868 11396
rect 42588 11342 42590 11394
rect 42642 11342 42814 11394
rect 42866 11342 42868 11394
rect 42588 11340 42868 11342
rect 42588 11330 42644 11340
rect 41580 11116 41692 11172
rect 41636 11060 41692 11116
rect 41020 10658 41076 10668
rect 41487 11004 41692 11060
rect 41487 10666 41543 11004
rect 40012 10558 40014 10610
rect 40066 10558 40068 10610
rect 40012 10546 40068 10558
rect 41244 10612 41300 10622
rect 41487 10614 41489 10666
rect 41541 10614 41543 10666
rect 41487 10602 41543 10614
rect 42364 10612 42420 10622
rect 42364 10610 42644 10612
rect 41244 10518 41300 10556
rect 42364 10558 42366 10610
rect 42418 10558 42644 10610
rect 42364 10556 42644 10558
rect 42364 10546 42420 10556
rect 39788 10332 40068 10388
rect 39564 9996 39732 10052
rect 39228 8194 39284 8204
rect 39340 9884 39620 9940
rect 37996 7924 38052 7934
rect 37884 7868 37996 7924
rect 37996 7858 38052 7868
rect 37772 7634 37828 7644
rect 37996 7588 38052 7598
rect 37716 7532 37772 7542
rect 37716 7530 37940 7532
rect 37716 7478 37718 7530
rect 37770 7478 37940 7530
rect 37716 7476 37940 7478
rect 37716 7466 37772 7476
rect 37660 7362 37716 7374
rect 37660 7310 37662 7362
rect 37714 7310 37716 7362
rect 37660 7252 37716 7310
rect 37884 7364 37940 7476
rect 37996 7474 38052 7532
rect 37996 7422 37998 7474
rect 38050 7422 38052 7474
rect 38687 7530 38743 8092
rect 39004 8082 39060 8092
rect 39340 7924 39396 9884
rect 39564 9826 39620 9884
rect 39564 9774 39566 9826
rect 39618 9774 39620 9826
rect 39564 9762 39620 9774
rect 39452 9716 39508 9726
rect 39452 9492 39508 9660
rect 39452 9436 39620 9492
rect 39564 9210 39620 9436
rect 39564 9158 39566 9210
rect 39618 9158 39620 9210
rect 39564 9146 39620 9158
rect 39676 9156 39732 9996
rect 39900 9828 39956 9838
rect 39900 9734 39956 9772
rect 39676 9100 39788 9156
rect 39732 9098 39788 9100
rect 39452 9044 39508 9054
rect 39732 9046 39734 9098
rect 39786 9046 39788 9098
rect 39732 9034 39788 9046
rect 39452 8950 39508 8988
rect 39900 8484 39956 8494
rect 39788 8260 39844 8270
rect 39788 8166 39844 8204
rect 38687 7478 38689 7530
rect 38741 7478 38743 7530
rect 38687 7466 38743 7478
rect 38892 7868 39396 7924
rect 39564 7924 39620 7934
rect 37996 7410 38052 7422
rect 37884 7298 37940 7308
rect 38444 7364 38500 7374
rect 38444 7270 38500 7308
rect 37660 7186 37716 7196
rect 37324 6300 37492 6356
rect 37548 6916 37604 6926
rect 37324 6074 37380 6300
rect 37324 6022 37326 6074
rect 37378 6022 37380 6074
rect 37324 6010 37380 6022
rect 37436 5908 37492 5918
rect 37548 5908 37604 6860
rect 38892 6916 38948 7868
rect 39564 7474 39620 7868
rect 39564 7422 39566 7474
rect 39618 7422 39620 7474
rect 39564 7410 39620 7422
rect 39900 7362 39956 8428
rect 40012 7518 40068 10332
rect 40180 10386 40236 10398
rect 40180 10334 40182 10386
rect 40234 10334 40236 10386
rect 40180 9828 40236 10334
rect 40180 9762 40236 9772
rect 40684 9826 40740 9838
rect 40684 9774 40686 9826
rect 40738 9774 40740 9826
rect 40460 9716 40516 9726
rect 40348 9268 40404 9278
rect 40012 7466 40014 7518
rect 40066 7466 40068 7518
rect 40012 7454 40068 7466
rect 40124 9042 40180 9054
rect 40124 8990 40126 9042
rect 40178 8990 40180 9042
rect 39900 7310 39902 7362
rect 39954 7310 39956 7362
rect 39900 7298 39956 7310
rect 40124 7252 40180 8990
rect 40348 8230 40404 9212
rect 40348 8178 40350 8230
rect 40402 8178 40404 8230
rect 40348 8166 40404 8178
rect 40348 7476 40404 7486
rect 40460 7476 40516 9660
rect 40684 8484 40740 9774
rect 42588 9716 42644 10556
rect 42588 9622 42644 9660
rect 41020 8932 41076 8942
rect 41020 8838 41076 8876
rect 40684 8418 40740 8428
rect 40348 7474 40516 7476
rect 40348 7422 40350 7474
rect 40402 7422 40516 7474
rect 40908 8260 40964 8270
rect 40908 7501 40964 8204
rect 41692 8036 41748 8046
rect 41692 7942 41748 7980
rect 40908 7449 40910 7501
rect 40962 7449 40964 7501
rect 40908 7437 40964 7449
rect 42252 7476 42308 7486
rect 40348 7420 40516 7422
rect 40348 7410 40404 7420
rect 42252 7382 42308 7420
rect 40124 7186 40180 7196
rect 42700 7140 42756 11340
rect 42812 11330 42868 11340
rect 43148 11340 43428 11396
rect 43540 11396 43596 11406
rect 42980 11172 43036 11182
rect 42980 11078 43036 11116
rect 43148 10948 43204 11340
rect 43540 11302 43596 11340
rect 43055 10892 43204 10948
rect 43055 10666 43111 10892
rect 43055 10614 43057 10666
rect 43109 10614 43111 10666
rect 43055 10602 43111 10614
rect 43932 10612 43988 10650
rect 43932 10546 43988 10556
rect 42812 10386 42868 10398
rect 42812 10334 42814 10386
rect 42866 10334 42868 10386
rect 42812 7588 42868 10334
rect 43820 10164 43876 10174
rect 42924 9826 42980 9838
rect 42924 9774 42926 9826
rect 42978 9774 42980 9826
rect 42924 9716 42980 9774
rect 42924 9650 42980 9660
rect 43092 9602 43148 9614
rect 43092 9550 43094 9602
rect 43146 9550 43148 9602
rect 43092 9044 43148 9550
rect 43820 9062 43876 10108
rect 44156 9828 44212 12002
rect 44268 11396 44324 11406
rect 44380 11396 44436 12796
rect 44324 11340 44436 11396
rect 44268 11302 44324 11340
rect 44380 11172 44436 11182
rect 44268 9828 44324 9838
rect 44156 9826 44324 9828
rect 44156 9774 44270 9826
rect 44322 9774 44324 9826
rect 44156 9772 44324 9774
rect 43932 9604 43988 9614
rect 43932 9510 43988 9548
rect 44268 9492 44324 9772
rect 44268 9426 44324 9436
rect 43092 8978 43148 8988
rect 43708 9044 43764 9054
rect 43708 8950 43764 8988
rect 43820 9010 43822 9062
rect 43874 9010 43876 9062
rect 42812 7522 42868 7532
rect 42924 8930 42980 8942
rect 42924 8878 42926 8930
rect 42978 8878 42980 8930
rect 42924 7364 42980 8878
rect 43820 8932 43876 9010
rect 43820 8596 43876 8876
rect 43988 8820 44044 8830
rect 43988 8818 44212 8820
rect 43988 8766 43990 8818
rect 44042 8766 44212 8818
rect 43988 8764 44212 8766
rect 43988 8754 44044 8764
rect 43820 8540 44100 8596
rect 43932 8260 43988 8270
rect 43820 8258 43988 8260
rect 43820 8206 43934 8258
rect 43986 8206 43988 8258
rect 43820 8204 43988 8206
rect 43820 7489 43876 8204
rect 43932 8194 43988 8204
rect 43820 7476 43822 7489
rect 43874 7476 43876 7489
rect 43820 7410 43876 7420
rect 44044 7474 44100 8540
rect 44044 7422 44046 7474
rect 44098 7422 44100 7474
rect 44044 7410 44100 7422
rect 42924 7298 42980 7308
rect 43708 7364 43764 7374
rect 43708 7270 43764 7308
rect 42700 7084 43092 7140
rect 38892 6850 38948 6860
rect 37660 6690 37716 6702
rect 37660 6638 37662 6690
rect 37714 6638 37716 6690
rect 39228 6692 39284 6702
rect 37660 6580 37716 6638
rect 37660 6514 37716 6524
rect 38780 6662 38836 6674
rect 38780 6610 38782 6662
rect 38834 6610 38836 6662
rect 37436 5906 37604 5908
rect 37436 5854 37438 5906
rect 37490 5854 37604 5906
rect 37436 5852 37604 5854
rect 37436 5842 37492 5852
rect 38780 5796 38836 6610
rect 38780 5730 38836 5740
rect 38892 5908 38948 5918
rect 36876 5070 36878 5122
rect 36930 5070 36932 5122
rect 36876 5058 36932 5070
rect 36988 5404 37268 5460
rect 36764 4844 36932 4900
rect 36764 3780 36820 3790
rect 36652 3778 36820 3780
rect 36652 3726 36766 3778
rect 36818 3726 36820 3778
rect 36652 3724 36820 3726
rect 36764 3714 36820 3724
rect 36428 3502 36430 3554
rect 36482 3502 36484 3554
rect 36428 3490 36484 3502
rect 24556 3462 24612 3474
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 36876 2772 36932 4844
rect 36988 4450 37044 5404
rect 37660 5124 37716 5134
rect 37660 5030 37716 5068
rect 38780 5124 38836 5134
rect 38500 4900 38556 4910
rect 36988 4398 36990 4450
rect 37042 4398 37044 4450
rect 36988 4386 37044 4398
rect 37231 4564 37287 4574
rect 37231 4394 37287 4508
rect 38500 4562 38556 4844
rect 38500 4510 38502 4562
rect 38554 4510 38556 4562
rect 38500 4498 38556 4510
rect 37231 4342 37233 4394
rect 37285 4342 37287 4394
rect 37231 4330 37287 4342
rect 38108 4340 38164 4350
rect 38332 4340 38388 4350
rect 38108 4338 38388 4340
rect 38108 4286 38110 4338
rect 38162 4286 38334 4338
rect 38386 4286 38388 4338
rect 38108 4284 38388 4286
rect 38108 4274 38164 4284
rect 38332 4228 38388 4284
rect 38332 4162 38388 4172
rect 38556 4340 38612 4350
rect 38556 3678 38612 4284
rect 38500 3666 38612 3678
rect 38500 3614 38502 3666
rect 38554 3614 38612 3666
rect 38500 3612 38612 3614
rect 38780 3666 38836 5068
rect 38780 3614 38782 3666
rect 38834 3614 38836 3666
rect 38500 3602 38556 3612
rect 38780 3602 38836 3614
rect 38892 3539 38948 5852
rect 39228 4450 39284 6636
rect 41356 6580 41412 6590
rect 41356 6486 41412 6524
rect 43036 6580 43092 7084
rect 40124 6468 40180 6478
rect 40124 6374 40180 6412
rect 39564 6244 39620 6254
rect 39340 5908 39396 5918
rect 39340 5794 39396 5852
rect 39340 5742 39342 5794
rect 39394 5742 39396 5794
rect 39340 5730 39396 5742
rect 39564 5234 39620 6188
rect 39564 5182 39566 5234
rect 39618 5182 39620 5234
rect 39564 4900 39620 5182
rect 39228 4398 39230 4450
rect 39282 4398 39284 4450
rect 39228 4386 39284 4398
rect 39471 4844 39620 4900
rect 39676 6132 39732 6142
rect 39471 4394 39527 4844
rect 38892 3487 38894 3539
rect 38946 3487 38948 3539
rect 39116 4340 39172 4350
rect 39471 4342 39473 4394
rect 39525 4342 39527 4394
rect 39471 4330 39527 4342
rect 39116 3554 39172 4284
rect 39676 3780 39732 6076
rect 40908 6132 40964 6142
rect 40236 5933 40292 5945
rect 40236 5881 40238 5933
rect 40290 5881 40292 5933
rect 40236 5796 40292 5881
rect 40908 5906 40964 6076
rect 41692 6020 41748 6030
rect 41692 5933 41748 5964
rect 40908 5854 40910 5906
rect 40962 5854 40964 5906
rect 40908 5842 40964 5854
rect 41244 5921 41300 5933
rect 41244 5908 41246 5921
rect 41298 5908 41300 5921
rect 41692 5881 41694 5933
rect 41746 5881 41748 5933
rect 41692 5869 41748 5881
rect 41244 5829 41300 5852
rect 40236 5730 40292 5740
rect 41356 5796 41412 5806
rect 42700 5796 42756 5806
rect 41356 5794 41860 5796
rect 41356 5742 41358 5794
rect 41410 5742 41860 5794
rect 41356 5740 41860 5742
rect 41356 5730 41412 5740
rect 39900 5236 39956 5246
rect 39900 5122 39956 5180
rect 39900 5070 39902 5122
rect 39954 5070 39956 5122
rect 39900 5058 39956 5070
rect 40684 5124 40740 5134
rect 40684 5030 40740 5068
rect 40348 5012 40404 5022
rect 40348 4340 40404 4956
rect 40348 4246 40404 4284
rect 41356 4228 41412 4238
rect 41356 4134 41412 4172
rect 39676 3724 39956 3780
rect 39900 3666 39956 3724
rect 39900 3614 39902 3666
rect 39954 3614 39956 3666
rect 39900 3602 39956 3614
rect 41804 3666 41860 5740
rect 42700 5702 42756 5740
rect 43036 5122 43092 6524
rect 43260 6802 43316 6814
rect 43260 6750 43262 6802
rect 43314 6750 43316 6802
rect 43036 5070 43038 5122
rect 43090 5070 43092 5122
rect 43036 5058 43092 5070
rect 43148 6468 43204 6478
rect 43148 5124 43204 6412
rect 43260 5236 43316 6750
rect 44044 6692 44100 6702
rect 44156 6692 44212 8764
rect 44044 6690 44212 6692
rect 44044 6638 44046 6690
rect 44098 6638 44212 6690
rect 44044 6636 44212 6638
rect 44044 6626 44100 6636
rect 44380 6468 44436 11116
rect 44044 6412 44436 6468
rect 43932 5348 43988 5358
rect 43932 5254 43988 5292
rect 43484 5236 43540 5246
rect 43260 5234 43540 5236
rect 43260 5182 43486 5234
rect 43538 5182 43540 5234
rect 43260 5180 43540 5182
rect 43484 5170 43540 5180
rect 43148 5092 43428 5124
rect 43148 5068 43318 5092
rect 43316 5040 43318 5068
rect 43370 5040 43428 5092
rect 43316 5028 43428 5040
rect 41804 3614 41806 3666
rect 41858 3614 41860 3666
rect 41804 3602 41860 3614
rect 42140 5012 42196 5022
rect 39116 3502 39118 3554
rect 39170 3502 39172 3554
rect 39116 3490 39172 3502
rect 38892 3475 38948 3487
rect 42140 3444 42196 4956
rect 42588 5012 42644 5022
rect 43372 5012 43428 5028
rect 43372 4956 43764 5012
rect 42588 4918 42644 4956
rect 43260 4226 43316 4238
rect 43260 4174 43262 4226
rect 43314 4174 43316 4226
rect 42868 3722 42924 3734
rect 42868 3670 42870 3722
rect 42922 3670 42924 3722
rect 42868 3668 42924 3670
rect 42588 3612 42924 3668
rect 43260 3668 43316 4174
rect 43596 3668 43652 3678
rect 43260 3666 43652 3668
rect 43260 3614 43598 3666
rect 43650 3614 43652 3666
rect 43260 3612 43652 3614
rect 42588 3554 42644 3612
rect 43596 3602 43652 3612
rect 42588 3502 42590 3554
rect 42642 3502 42644 3554
rect 43708 3539 43764 4956
rect 44044 4338 44100 6412
rect 44268 6132 44324 6142
rect 44268 5460 44324 6076
rect 44268 5122 44324 5404
rect 44268 5070 44270 5122
rect 44322 5070 44324 5122
rect 44268 5058 44324 5070
rect 44044 4286 44046 4338
rect 44098 4286 44100 4338
rect 44044 4274 44100 4286
rect 42588 3490 42644 3502
rect 42700 3498 42756 3510
rect 42140 3378 42196 3388
rect 42700 3446 42702 3498
rect 42754 3446 42756 3498
rect 43708 3487 43710 3539
rect 43762 3487 43764 3539
rect 43932 4228 43988 4238
rect 43932 3554 43988 4172
rect 43932 3502 43934 3554
rect 43986 3502 43988 3554
rect 43932 3490 43988 3502
rect 43708 3475 43764 3487
rect 42700 3444 42756 3446
rect 42700 3378 42756 3388
rect 36876 2706 36932 2716
<< via2 >>
rect 41692 43036 41748 43092
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 20748 39564 20804 39620
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19740 38834 19796 38836
rect 19740 38782 19742 38834
rect 19742 38782 19794 38834
rect 19794 38782 19796 38834
rect 19740 38780 19796 38782
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 21532 39116 21588 39172
rect 20748 38780 20804 38836
rect 20188 38668 20244 38724
rect 21868 38668 21924 38724
rect 20748 38050 20804 38052
rect 20748 37998 20750 38050
rect 20750 37998 20802 38050
rect 20802 37998 20804 38050
rect 20748 37996 20804 37998
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20188 37324 20244 37380
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 6076 33346 6132 33348
rect 6076 33294 6078 33346
rect 6078 33294 6130 33346
rect 6130 33294 6132 33346
rect 6076 33292 6132 33294
rect 10424 35698 10480 35700
rect 10424 35646 10426 35698
rect 10426 35646 10478 35698
rect 10478 35646 10480 35698
rect 10424 35644 10480 35646
rect 11116 35644 11172 35700
rect 10332 35308 10388 35364
rect 9100 35084 9156 35140
rect 8652 33292 8708 33348
rect 9100 33346 9156 33348
rect 9100 33294 9102 33346
rect 9102 33294 9154 33346
rect 9154 33294 9156 33346
rect 9100 33292 9156 33294
rect 11004 35196 11060 35252
rect 11004 34524 11060 34580
rect 11695 35308 11751 35364
rect 11452 35196 11508 35252
rect 12572 35698 12628 35700
rect 12572 35646 12574 35698
rect 12574 35646 12626 35698
rect 12626 35646 12628 35698
rect 12572 35644 12628 35646
rect 12012 35084 12068 35140
rect 10668 34076 10724 34132
rect 11004 34130 11060 34132
rect 11004 34078 11006 34130
rect 11006 34078 11058 34130
rect 11058 34078 11060 34130
rect 11004 34076 11060 34078
rect 9772 33404 9828 33460
rect 9884 33852 9940 33908
rect 11788 34524 11844 34580
rect 11116 33740 11172 33796
rect 11788 33458 11844 33460
rect 11788 33406 11790 33458
rect 11790 33406 11842 33458
rect 11842 33406 11844 33458
rect 11788 33404 11844 33406
rect 12292 33740 12348 33796
rect 13020 34636 13076 34692
rect 13020 34076 13076 34132
rect 13356 35084 13412 35140
rect 13692 34690 13748 34692
rect 13692 34638 13694 34690
rect 13694 34638 13746 34690
rect 13746 34638 13748 34690
rect 13692 34636 13748 34638
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 21532 37324 21588 37380
rect 20636 37100 20692 37156
rect 20524 36988 20580 37044
rect 21644 37100 21700 37156
rect 23100 40124 23156 40180
rect 24668 41132 24724 41188
rect 23212 40348 23268 40404
rect 22648 39452 22704 39508
rect 22988 39116 23044 39172
rect 23940 40348 23996 40404
rect 24444 40290 24500 40292
rect 24444 40238 24446 40290
rect 24446 40238 24498 40290
rect 24498 40238 24500 40290
rect 24444 40236 24500 40238
rect 23436 40124 23492 40180
rect 24332 39676 24388 39732
rect 24108 39618 24164 39620
rect 24108 39566 24110 39618
rect 24110 39566 24162 39618
rect 24162 39566 24164 39618
rect 24108 39564 24164 39566
rect 23436 38892 23492 38948
rect 23548 39452 23604 39508
rect 22988 38050 23044 38052
rect 22988 37998 22990 38050
rect 22990 37998 23042 38050
rect 23042 37998 23044 38050
rect 22988 37996 23044 37998
rect 22316 37772 22372 37828
rect 21980 37548 22036 37604
rect 22652 37324 22708 37380
rect 22316 37266 22372 37268
rect 22316 37214 22318 37266
rect 22318 37214 22370 37266
rect 22370 37214 22372 37266
rect 22316 37212 22372 37214
rect 26012 41186 26068 41188
rect 26012 41134 26014 41186
rect 26014 41134 26066 41186
rect 26066 41134 26068 41186
rect 26012 41132 26068 41134
rect 24780 41020 24836 41076
rect 25732 41074 25788 41076
rect 25732 41022 25734 41074
rect 25734 41022 25786 41074
rect 25786 41022 25788 41074
rect 25732 41020 25788 41022
rect 26236 40908 26292 40964
rect 25116 40402 25172 40404
rect 25116 40350 25118 40402
rect 25118 40350 25170 40402
rect 25170 40350 25172 40402
rect 25116 40348 25172 40350
rect 24332 38892 24388 38948
rect 24108 38108 24164 38164
rect 25900 40290 25956 40292
rect 25900 40238 25902 40290
rect 25902 40238 25954 40290
rect 25954 40238 25956 40290
rect 25900 40236 25956 40238
rect 23660 37996 23716 38052
rect 23436 37884 23492 37940
rect 23100 37212 23156 37268
rect 23436 37266 23492 37268
rect 23436 37214 23438 37266
rect 23438 37214 23490 37266
rect 23490 37214 23492 37266
rect 23436 37212 23492 37214
rect 23828 38050 23884 38052
rect 23828 37998 23830 38050
rect 23830 37998 23882 38050
rect 23882 37998 23884 38050
rect 23828 37996 23884 37998
rect 23940 37548 23996 37604
rect 22876 37100 22932 37156
rect 21868 36988 21924 37044
rect 22652 36988 22708 37044
rect 22148 36594 22204 36596
rect 22148 36542 22150 36594
rect 22150 36542 22202 36594
rect 22202 36542 22204 36594
rect 22148 36540 22204 36542
rect 21756 36428 21812 36484
rect 21980 36428 22036 36484
rect 21868 36316 21924 36372
rect 14028 33740 14084 33796
rect 14812 33740 14868 33796
rect 13132 33628 13188 33684
rect 12908 33404 12964 33460
rect 12460 33180 12516 33236
rect 9660 32508 9716 32564
rect 10332 32562 10388 32564
rect 10332 32510 10334 32562
rect 10334 32510 10386 32562
rect 10386 32510 10388 32562
rect 10332 32508 10388 32510
rect 8316 32284 8372 32340
rect 12460 32284 12516 32340
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 15820 33628 15876 33684
rect 15932 33292 15988 33348
rect 16156 33404 16212 33460
rect 15036 32284 15092 32340
rect 15596 31778 15652 31780
rect 15596 31726 15598 31778
rect 15598 31726 15650 31778
rect 15650 31726 15652 31778
rect 15596 31724 15652 31726
rect 13916 30492 13972 30548
rect 17388 34914 17444 34916
rect 17388 34862 17390 34914
rect 17390 34862 17442 34914
rect 17442 34862 17444 34914
rect 17388 34860 17444 34862
rect 17276 33628 17332 33684
rect 21420 35308 21476 35364
rect 18172 33740 18228 33796
rect 16772 33570 16828 33572
rect 16772 33518 16774 33570
rect 16774 33518 16826 33570
rect 16826 33518 16828 33570
rect 16772 33516 16828 33518
rect 16268 31724 16324 31780
rect 17052 33346 17108 33348
rect 17052 33294 17054 33346
rect 17054 33294 17106 33346
rect 17106 33294 17108 33346
rect 17052 33292 17108 33294
rect 16604 32620 16660 32676
rect 15148 30492 15204 30548
rect 14812 30210 14868 30212
rect 14812 30158 14814 30210
rect 14814 30158 14866 30210
rect 14866 30158 14868 30210
rect 14812 30156 14868 30158
rect 12684 29148 12740 29204
rect 13468 29148 13524 29204
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 15148 29036 15204 29092
rect 16044 30156 16100 30212
rect 17444 32338 17500 32340
rect 17444 32286 17446 32338
rect 17446 32286 17498 32338
rect 17498 32286 17500 32338
rect 17444 32284 17500 32286
rect 17948 33068 18004 33124
rect 17724 32620 17780 32676
rect 18620 34914 18676 34916
rect 18620 34862 18622 34914
rect 18622 34862 18674 34914
rect 18674 34862 18676 34914
rect 18620 34860 18676 34862
rect 24444 38050 24500 38052
rect 24444 37998 24446 38050
rect 24446 37998 24498 38050
rect 24498 37998 24500 38050
rect 24444 37996 24500 37998
rect 25004 37884 25060 37940
rect 24108 36988 24164 37044
rect 22988 36540 23044 36596
rect 22764 36482 22820 36484
rect 22764 36430 22766 36482
rect 22766 36430 22818 36482
rect 22818 36430 22820 36482
rect 22764 36428 22820 36430
rect 23268 36370 23324 36372
rect 23268 36318 23270 36370
rect 23270 36318 23322 36370
rect 23322 36318 23324 36370
rect 23268 36316 23324 36318
rect 22092 35308 22148 35364
rect 23436 35644 23492 35700
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 18284 33516 18340 33572
rect 18396 33292 18452 33348
rect 18172 33234 18228 33236
rect 18172 33182 18174 33234
rect 18174 33182 18226 33234
rect 18226 33182 18228 33234
rect 18172 33180 18228 33182
rect 18172 32508 18228 32564
rect 16716 30492 16772 30548
rect 17612 31724 17668 31780
rect 19964 33068 20020 33124
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19292 32620 19348 32676
rect 17836 30604 17892 30660
rect 17724 30268 17780 30324
rect 18620 29932 18676 29988
rect 17052 29148 17108 29204
rect 10444 27804 10500 27860
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 11788 27858 11844 27860
rect 11788 27806 11790 27858
rect 11790 27806 11842 27858
rect 11842 27806 11844 27858
rect 11788 27804 11844 27806
rect 12796 27804 12852 27860
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 10220 26290 10276 26292
rect 10220 26238 10222 26290
rect 10222 26238 10274 26290
rect 10274 26238 10276 26290
rect 10220 26236 10276 26238
rect 17836 29260 17892 29316
rect 18956 29260 19012 29316
rect 14140 27298 14196 27300
rect 14140 27246 14142 27298
rect 14142 27246 14194 27298
rect 14194 27246 14196 27298
rect 14140 27244 14196 27246
rect 12684 26236 12740 26292
rect 11116 25452 11172 25508
rect 9884 25228 9940 25284
rect 10332 25228 10388 25284
rect 10892 25116 10948 25172
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 10276 24050 10332 24052
rect 10276 23998 10278 24050
rect 10278 23998 10330 24050
rect 10330 23998 10332 24050
rect 10276 23996 10332 23998
rect 11228 25228 11284 25284
rect 10892 23996 10948 24052
rect 9884 23212 9940 23268
rect 10556 23212 10612 23268
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 6300 20690 6356 20692
rect 6300 20638 6302 20690
rect 6302 20638 6354 20690
rect 6354 20638 6356 20690
rect 6300 20636 6356 20638
rect 8260 21532 8316 21588
rect 9436 21586 9492 21588
rect 9436 21534 9438 21586
rect 9438 21534 9490 21586
rect 9490 21534 9492 21586
rect 9436 21532 9492 21534
rect 9772 22876 9828 22932
rect 11452 25228 11508 25284
rect 12236 25228 12292 25284
rect 12348 25340 12404 25396
rect 13020 25506 13076 25508
rect 13020 25454 13022 25506
rect 13022 25454 13074 25506
rect 13074 25454 13076 25506
rect 13020 25452 13076 25454
rect 13356 25340 13412 25396
rect 11676 23212 11732 23268
rect 10892 23154 10948 23156
rect 10892 23102 10894 23154
rect 10894 23102 10946 23154
rect 10946 23102 10948 23154
rect 10892 23100 10948 23102
rect 12796 23100 12852 23156
rect 10780 22988 10836 23044
rect 12572 22988 12628 23044
rect 12684 22930 12740 22932
rect 12684 22878 12686 22930
rect 12686 22878 12738 22930
rect 12738 22878 12740 22930
rect 12684 22876 12740 22878
rect 12796 22316 12852 22372
rect 14588 27132 14644 27188
rect 14476 27074 14532 27076
rect 14476 27022 14478 27074
rect 14478 27022 14530 27074
rect 14530 27022 14532 27074
rect 14476 27020 14532 27022
rect 15596 27186 15652 27188
rect 15596 27134 15598 27186
rect 15598 27134 15650 27186
rect 15650 27134 15652 27186
rect 15596 27132 15652 27134
rect 15148 25004 15204 25060
rect 15708 24220 15764 24276
rect 14812 23996 14868 24052
rect 15596 24050 15652 24052
rect 15596 23998 15598 24050
rect 15598 23998 15650 24050
rect 15650 23998 15652 24050
rect 15596 23996 15652 23998
rect 14252 23884 14308 23940
rect 15708 23923 15764 23940
rect 15708 23884 15710 23923
rect 15710 23884 15762 23923
rect 15762 23884 15764 23923
rect 18844 27244 18900 27300
rect 19068 27132 19124 27188
rect 16604 25004 16660 25060
rect 17836 26290 17892 26292
rect 17836 26238 17838 26290
rect 17838 26238 17890 26290
rect 17890 26238 17892 26290
rect 17836 26236 17892 26238
rect 18732 26290 18788 26292
rect 18732 26238 18734 26290
rect 18734 26238 18786 26290
rect 18786 26238 18788 26290
rect 18732 26236 18788 26238
rect 16828 24668 16884 24724
rect 19628 31724 19684 31780
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20076 30380 20132 30436
rect 19908 30156 19964 30212
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19740 29538 19796 29540
rect 19740 29486 19742 29538
rect 19742 29486 19794 29538
rect 19794 29486 19796 29538
rect 19740 29484 19796 29486
rect 20300 29484 20356 29540
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20748 33068 20804 33124
rect 21644 32562 21700 32564
rect 21644 32510 21646 32562
rect 21646 32510 21698 32562
rect 21698 32510 21700 32562
rect 21644 32508 21700 32510
rect 23268 35308 23324 35364
rect 28644 40908 28700 40964
rect 27020 40236 27076 40292
rect 27356 39730 27412 39732
rect 27356 39678 27358 39730
rect 27358 39678 27410 39730
rect 27410 39678 27412 39730
rect 27356 39676 27412 39678
rect 27468 39564 27524 39620
rect 25676 38050 25732 38052
rect 25676 37998 25678 38050
rect 25678 37998 25730 38050
rect 25730 37998 25732 38050
rect 25676 37996 25732 37998
rect 26460 38050 26516 38052
rect 26460 37998 26462 38050
rect 26462 37998 26514 38050
rect 26514 37998 26516 38050
rect 26460 37996 26516 37998
rect 26964 38050 27020 38052
rect 26964 37998 26966 38050
rect 26966 37998 27018 38050
rect 27018 37998 27020 38050
rect 26964 37996 27020 37998
rect 27244 38050 27300 38052
rect 27244 37998 27246 38050
rect 27246 37998 27298 38050
rect 27298 37998 27300 38050
rect 27244 37996 27300 37998
rect 27468 38780 27524 38836
rect 28364 40236 28420 40292
rect 28028 38780 28084 38836
rect 27804 37996 27860 38052
rect 27468 37884 27524 37940
rect 26236 37772 26292 37828
rect 27580 37772 27636 37828
rect 26236 37100 26292 37156
rect 26348 36988 26404 37044
rect 25676 35644 25732 35700
rect 25956 35868 26012 35924
rect 26124 35698 26180 35700
rect 26124 35646 26126 35698
rect 26126 35646 26178 35698
rect 26178 35646 26180 35698
rect 26124 35644 26180 35646
rect 26852 37042 26908 37044
rect 26852 36990 26854 37042
rect 26854 36990 26906 37042
rect 26906 36990 26908 37042
rect 26852 36988 26908 36990
rect 27132 36876 27188 36932
rect 27412 37266 27468 37268
rect 27412 37214 27414 37266
rect 27414 37214 27466 37266
rect 27466 37214 27468 37266
rect 27412 37212 27468 37214
rect 28812 40348 28868 40404
rect 29708 39564 29764 39620
rect 31612 41970 31668 41972
rect 31612 41918 31614 41970
rect 31614 41918 31666 41970
rect 31666 41918 31668 41970
rect 31612 41916 31668 41918
rect 30940 41298 30996 41300
rect 30940 41246 30942 41298
rect 30942 41246 30994 41298
rect 30994 41246 30996 41298
rect 30940 41244 30996 41246
rect 31164 40572 31220 40628
rect 32284 40460 32340 40516
rect 33628 41916 33684 41972
rect 32396 40348 32452 40404
rect 33292 41298 33348 41300
rect 33292 41246 33294 41298
rect 33294 41246 33346 41298
rect 33346 41246 33348 41298
rect 33292 41244 33348 41246
rect 30268 39618 30324 39620
rect 30268 39566 30270 39618
rect 30270 39566 30322 39618
rect 30322 39566 30324 39618
rect 30268 39564 30324 39566
rect 28700 38834 28756 38836
rect 28700 38782 28702 38834
rect 28702 38782 28754 38834
rect 28754 38782 28756 38834
rect 28700 38780 28756 38782
rect 33180 40572 33236 40628
rect 33423 40460 33479 40516
rect 33628 40348 33684 40404
rect 34300 40402 34356 40404
rect 34300 40350 34302 40402
rect 34302 40350 34354 40402
rect 34354 40350 34356 40402
rect 34300 40348 34356 40350
rect 32844 39564 32900 39620
rect 33740 39618 33796 39620
rect 33740 39566 33742 39618
rect 33742 39566 33794 39618
rect 33794 39566 33796 39618
rect 33740 39564 33796 39566
rect 31052 39004 31108 39060
rect 32396 39058 32452 39060
rect 32396 39006 32398 39058
rect 32398 39006 32450 39058
rect 32450 39006 32452 39058
rect 32396 39004 32452 39006
rect 32956 39004 33012 39060
rect 29708 38780 29764 38836
rect 28364 38668 28420 38724
rect 29540 38668 29596 38724
rect 29260 38050 29316 38052
rect 29260 37998 29262 38050
rect 29262 37998 29314 38050
rect 29314 37998 29316 38050
rect 29260 37996 29316 37998
rect 29036 37884 29092 37940
rect 27020 36428 27076 36484
rect 26908 35868 26964 35924
rect 26628 35810 26684 35812
rect 26628 35758 26630 35810
rect 26630 35758 26682 35810
rect 26682 35758 26684 35810
rect 26628 35756 26684 35758
rect 25116 35308 25172 35364
rect 25676 35308 25732 35364
rect 25956 35308 26012 35364
rect 26908 35308 26964 35364
rect 27020 34748 27076 34804
rect 24556 34130 24612 34132
rect 24556 34078 24558 34130
rect 24558 34078 24610 34130
rect 24610 34078 24612 34130
rect 24556 34076 24612 34078
rect 24220 33628 24276 33684
rect 25452 34130 25508 34132
rect 25452 34078 25454 34130
rect 25454 34078 25506 34130
rect 25506 34078 25508 34130
rect 25452 34076 25508 34078
rect 24780 33740 24836 33796
rect 25284 33628 25340 33684
rect 24444 33292 24500 33348
rect 25452 33404 25508 33460
rect 26124 33458 26180 33460
rect 26124 33406 26126 33458
rect 26126 33406 26178 33458
rect 26178 33406 26180 33458
rect 26124 33404 26180 33406
rect 24668 33068 24724 33124
rect 20636 30434 20692 30436
rect 20636 30382 20638 30434
rect 20638 30382 20690 30434
rect 20690 30382 20692 30434
rect 20636 30380 20692 30382
rect 21980 31778 22036 31780
rect 21980 31726 21982 31778
rect 21982 31726 22034 31778
rect 22034 31726 22036 31778
rect 21980 31724 22036 31726
rect 21196 30380 21252 30436
rect 21980 30604 22036 30660
rect 21644 30156 21700 30212
rect 22876 30994 22932 30996
rect 22876 30942 22878 30994
rect 22878 30942 22930 30994
rect 22930 30942 22932 30994
rect 22876 30940 22932 30942
rect 20524 28418 20580 28420
rect 20524 28366 20526 28418
rect 20526 28366 20578 28418
rect 20578 28366 20580 28418
rect 20524 28364 20580 28366
rect 20300 27132 20356 27188
rect 19852 27074 19908 27076
rect 19852 27022 19854 27074
rect 19854 27022 19906 27074
rect 19906 27022 19908 27074
rect 19852 27020 19908 27022
rect 16716 24220 16772 24276
rect 16268 23884 16324 23940
rect 17836 25340 17892 25396
rect 17836 25116 17892 25172
rect 17276 24722 17332 24724
rect 17276 24670 17278 24722
rect 17278 24670 17330 24722
rect 17330 24670 17332 24722
rect 17276 24668 17332 24670
rect 17164 23938 17220 23940
rect 17164 23886 17166 23938
rect 17166 23886 17218 23938
rect 17218 23886 17220 23938
rect 17164 23884 17220 23886
rect 14476 23154 14532 23156
rect 14476 23102 14478 23154
rect 14478 23102 14530 23154
rect 14530 23102 14532 23154
rect 14476 23100 14532 23102
rect 13692 22764 13748 22820
rect 13580 22370 13636 22372
rect 13580 22318 13582 22370
rect 13582 22318 13634 22370
rect 13634 22318 13636 22370
rect 13580 22316 13636 22318
rect 9660 21420 9716 21476
rect 8092 20636 8148 20692
rect 8092 20076 8148 20132
rect 8036 19906 8092 19908
rect 8036 19854 8038 19906
rect 8038 19854 8090 19906
rect 8090 19854 8092 19906
rect 8036 19852 8092 19854
rect 8764 20076 8820 20132
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 8428 19404 8484 19460
rect 8764 19292 8820 19348
rect 8372 19180 8428 19236
rect 8316 18508 8372 18564
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 7980 18060 8036 18116
rect 4684 18004 4740 18006
rect 8988 21308 9044 21364
rect 12124 21474 12180 21476
rect 12124 21422 12126 21474
rect 12126 21422 12178 21474
rect 12178 21422 12180 21474
rect 12124 21420 12180 21422
rect 8988 19852 9044 19908
rect 9436 19180 9492 19236
rect 9772 19458 9828 19460
rect 9772 19406 9774 19458
rect 9774 19406 9826 19458
rect 9826 19406 9828 19458
rect 9772 19404 9828 19406
rect 12012 20748 12068 20804
rect 10220 20524 10276 20580
rect 12236 20524 12292 20580
rect 11004 19404 11060 19460
rect 10892 18508 10948 18564
rect 10220 18413 10222 18452
rect 10222 18413 10274 18452
rect 10274 18413 10276 18452
rect 10220 18396 10276 18413
rect 10444 18284 10500 18340
rect 9100 18060 9156 18116
rect 10108 18060 10164 18116
rect 8540 17724 8596 17780
rect 9100 16940 9156 16996
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 8764 16828 8820 16884
rect 7980 15708 8036 15764
rect 8092 15148 8148 15204
rect 8876 16380 8932 16436
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 7532 14700 7588 14756
rect 8428 14700 8484 14756
rect 7644 13804 7700 13860
rect 7756 14364 7812 14420
rect 8764 14642 8820 14644
rect 8764 14590 8766 14642
rect 8766 14590 8818 14642
rect 8818 14590 8820 14642
rect 8764 14588 8820 14590
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 8428 13916 8484 13972
rect 8540 13804 8596 13860
rect 8092 13709 8094 13748
rect 8094 13709 8146 13748
rect 8146 13709 8148 13748
rect 8092 13692 8148 13709
rect 8092 13020 8148 13076
rect 7364 12908 7420 12964
rect 8652 13692 8708 13748
rect 8988 15820 9044 15876
rect 9100 15148 9156 15204
rect 10220 17778 10276 17780
rect 10220 17726 10222 17778
rect 10222 17726 10274 17778
rect 10274 17726 10276 17778
rect 10220 17724 10276 17726
rect 11676 19234 11732 19236
rect 11676 19182 11678 19234
rect 11678 19182 11730 19234
rect 11730 19182 11732 19234
rect 11676 19180 11732 19182
rect 12012 18450 12068 18452
rect 12012 18398 12014 18450
rect 12014 18398 12066 18450
rect 12066 18398 12068 18450
rect 12012 18396 12068 18398
rect 14252 21474 14308 21476
rect 14252 21422 14254 21474
rect 14254 21422 14306 21474
rect 14306 21422 14308 21474
rect 14252 21420 14308 21422
rect 13448 21084 13504 21140
rect 13580 20802 13636 20804
rect 13580 20750 13582 20802
rect 13582 20750 13634 20802
rect 13634 20750 13636 20802
rect 13580 20748 13636 20750
rect 12552 19628 12608 19684
rect 13804 19346 13860 19348
rect 13804 19294 13806 19346
rect 13806 19294 13858 19346
rect 13858 19294 13860 19346
rect 13804 19292 13860 19294
rect 12684 19180 12740 19236
rect 12348 18396 12404 18452
rect 11452 18284 11508 18340
rect 13468 19234 13524 19236
rect 13468 19182 13470 19234
rect 13470 19182 13522 19234
rect 13522 19182 13524 19234
rect 13468 19180 13524 19182
rect 12796 19122 12852 19124
rect 12796 19070 12798 19122
rect 12798 19070 12850 19122
rect 12850 19070 12852 19122
rect 12796 19068 12852 19070
rect 13804 19068 13860 19124
rect 14476 21196 14532 21252
rect 15148 22876 15204 22932
rect 14812 20076 14868 20132
rect 14140 17836 14196 17892
rect 11228 17724 11284 17780
rect 11564 17666 11620 17668
rect 11564 17614 11566 17666
rect 11566 17614 11618 17666
rect 11618 17614 11620 17666
rect 11564 17612 11620 17614
rect 12440 17388 12496 17444
rect 10444 16940 10500 16996
rect 12796 17052 12852 17108
rect 12124 16882 12180 16884
rect 12124 16830 12126 16882
rect 12126 16830 12178 16882
rect 12178 16830 12180 16882
rect 12124 16828 12180 16830
rect 10220 15820 10276 15876
rect 10556 15820 10612 15876
rect 11564 15538 11620 15540
rect 11564 15486 11566 15538
rect 11566 15486 11618 15538
rect 11618 15486 11620 15538
rect 11564 15484 11620 15486
rect 11452 15148 11508 15204
rect 11564 14588 11620 14644
rect 9660 13858 9716 13860
rect 9660 13806 9662 13858
rect 9662 13806 9714 13858
rect 9714 13806 9716 13858
rect 9660 13804 9716 13806
rect 11340 13692 11396 13748
rect 8540 13580 8596 13636
rect 8988 13020 9044 13076
rect 9436 12908 9492 12964
rect 8204 12124 8260 12180
rect 10220 12178 10276 12180
rect 10220 12126 10222 12178
rect 10222 12126 10274 12178
rect 10274 12126 10276 12178
rect 10220 12124 10276 12126
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 12552 15596 12608 15652
rect 11676 13580 11732 13636
rect 12012 15484 12068 15540
rect 13244 16940 13300 16996
rect 12908 16828 12964 16884
rect 12684 15484 12740 15540
rect 13468 16828 13524 16884
rect 13580 16492 13636 16548
rect 13468 15820 13524 15876
rect 12124 14364 12180 14420
rect 13132 13804 13188 13860
rect 14344 17666 14400 17668
rect 14344 17614 14346 17666
rect 14346 17614 14398 17666
rect 14398 17614 14400 17666
rect 14344 17612 14400 17614
rect 15372 21756 15428 21812
rect 16156 23100 16212 23156
rect 15708 21756 15764 21812
rect 15932 21644 15988 21700
rect 15708 21084 15764 21140
rect 15596 20972 15652 21028
rect 15036 20076 15092 20132
rect 15372 19628 15428 19684
rect 15932 21084 15988 21140
rect 16940 21084 16996 21140
rect 17612 20972 17668 21028
rect 19180 25228 19236 25284
rect 18060 23996 18116 24052
rect 18620 24050 18676 24052
rect 18620 23998 18622 24050
rect 18622 23998 18674 24050
rect 18674 23998 18676 24050
rect 18620 23996 18676 23998
rect 18956 23938 19012 23940
rect 18956 23886 18958 23938
rect 18958 23886 19010 23938
rect 19010 23886 19012 23938
rect 18956 23884 19012 23886
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20188 26684 20244 26740
rect 20044 26628 20100 26630
rect 20412 27020 20468 27076
rect 20412 26796 20468 26852
rect 20860 27244 20916 27300
rect 22204 28364 22260 28420
rect 21532 27804 21588 27860
rect 21308 27132 21364 27188
rect 20860 27074 20916 27076
rect 20860 27022 20862 27074
rect 20862 27022 20914 27074
rect 20914 27022 20916 27074
rect 20860 27020 20916 27022
rect 20524 26908 20580 26964
rect 21532 26908 21588 26964
rect 21420 26796 21476 26852
rect 20636 26460 20692 26516
rect 20188 25900 20244 25956
rect 20076 25394 20132 25396
rect 20076 25342 20078 25394
rect 20078 25342 20130 25394
rect 20130 25342 20132 25394
rect 20076 25340 20132 25342
rect 20524 25564 20580 25620
rect 20792 25900 20848 25956
rect 20188 25228 20244 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19404 23884 19460 23940
rect 19852 23938 19908 23940
rect 19852 23886 19854 23938
rect 19854 23886 19906 23938
rect 19906 23886 19908 23938
rect 19852 23884 19908 23886
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 17948 23212 18004 23268
rect 21084 23212 21140 23268
rect 21308 23212 21364 23268
rect 21196 23100 21252 23156
rect 23324 30828 23380 30884
rect 23212 29372 23268 29428
rect 23212 28588 23268 28644
rect 23100 28028 23156 28084
rect 22596 27298 22652 27300
rect 22596 27246 22598 27298
rect 22598 27246 22650 27298
rect 22650 27246 22652 27298
rect 22596 27244 22652 27246
rect 22652 27020 22708 27076
rect 21756 26460 21812 26516
rect 22148 26962 22204 26964
rect 22148 26910 22150 26962
rect 22150 26910 22202 26962
rect 22202 26910 22204 26962
rect 22148 26908 22204 26910
rect 21644 24556 21700 24612
rect 21644 23884 21700 23940
rect 22316 26514 22372 26516
rect 22316 26462 22318 26514
rect 22318 26462 22370 26514
rect 22370 26462 22372 26514
rect 22316 26460 22372 26462
rect 24332 32562 24388 32564
rect 24332 32510 24334 32562
rect 24334 32510 24386 32562
rect 24386 32510 24388 32562
rect 24332 32508 24388 32510
rect 27448 33346 27504 33348
rect 27448 33294 27450 33346
rect 27450 33294 27502 33346
rect 27502 33294 27504 33346
rect 27448 33292 27504 33294
rect 26572 33068 26628 33124
rect 25004 32956 25060 33012
rect 24892 32508 24948 32564
rect 24724 31890 24780 31892
rect 24724 31838 24726 31890
rect 24726 31838 24778 31890
rect 24778 31838 24780 31890
rect 24724 31836 24780 31838
rect 23548 31724 23604 31780
rect 23884 30210 23940 30212
rect 23884 30158 23886 30210
rect 23886 30158 23938 30210
rect 23938 30158 23940 30210
rect 23884 30156 23940 30158
rect 26460 32450 26516 32452
rect 26460 32398 26462 32450
rect 26462 32398 26514 32450
rect 26514 32398 26516 32450
rect 26460 32396 26516 32398
rect 27692 35698 27748 35700
rect 27692 35646 27694 35698
rect 27694 35646 27746 35698
rect 27746 35646 27748 35698
rect 27692 35644 27748 35646
rect 30268 36482 30324 36484
rect 30268 36430 30270 36482
rect 30270 36430 30322 36482
rect 30322 36430 30324 36482
rect 30268 36428 30324 36430
rect 29036 35756 29092 35812
rect 29596 36092 29652 36148
rect 29372 35644 29428 35700
rect 27916 35532 27972 35588
rect 30268 35532 30324 35588
rect 27972 35308 28028 35364
rect 28028 34748 28084 34804
rect 27692 31836 27748 31892
rect 27916 31890 27972 31892
rect 27916 31838 27918 31890
rect 27918 31838 27970 31890
rect 27970 31838 27972 31890
rect 27916 31836 27972 31838
rect 25452 31750 25508 31780
rect 25004 31388 25060 31444
rect 25452 31724 25454 31750
rect 25454 31724 25506 31750
rect 25506 31724 25508 31750
rect 25564 31276 25620 31332
rect 25228 30828 25284 30884
rect 25452 30828 25508 30884
rect 25788 31724 25844 31780
rect 27804 31724 27860 31780
rect 26012 31666 26068 31668
rect 26012 31614 26014 31666
rect 26014 31614 26066 31666
rect 26066 31614 26068 31666
rect 26012 31612 26068 31614
rect 26236 31500 26292 31556
rect 27244 31388 27300 31444
rect 26124 30716 26180 30772
rect 26348 30716 26404 30772
rect 23548 29932 23604 29988
rect 23884 29202 23940 29204
rect 23884 29150 23886 29202
rect 23886 29150 23938 29202
rect 23938 29150 23940 29202
rect 23884 29148 23940 29150
rect 23660 28476 23716 28532
rect 23548 28364 23604 28420
rect 23772 27916 23828 27972
rect 23772 27020 23828 27076
rect 25228 30210 25284 30212
rect 25228 30158 25230 30210
rect 25230 30158 25282 30210
rect 25282 30158 25284 30210
rect 25228 30156 25284 30158
rect 25788 30156 25844 30212
rect 25004 30044 25060 30100
rect 24556 29986 24612 29988
rect 24556 29934 24558 29986
rect 24558 29934 24610 29986
rect 24610 29934 24612 29986
rect 24556 29932 24612 29934
rect 24220 29426 24276 29428
rect 24220 29374 24222 29426
rect 24222 29374 24274 29426
rect 24274 29374 24276 29426
rect 24220 29372 24276 29374
rect 24220 29148 24276 29204
rect 24108 28642 24164 28644
rect 24108 28590 24110 28642
rect 24110 28590 24162 28642
rect 24162 28590 24164 28642
rect 24108 28588 24164 28590
rect 26460 30156 26516 30212
rect 25004 28812 25060 28868
rect 25116 29260 25172 29316
rect 23100 26290 23156 26292
rect 23100 26238 23102 26290
rect 23102 26238 23154 26290
rect 23154 26238 23156 26290
rect 23100 26236 23156 26238
rect 21980 25618 22036 25620
rect 21980 25566 21982 25618
rect 21982 25566 22034 25618
rect 22034 25566 22036 25618
rect 21980 25564 22036 25566
rect 23548 24556 23604 24612
rect 21868 23324 21924 23380
rect 21644 23212 21700 23268
rect 20860 22988 20916 23044
rect 21532 22988 21588 23044
rect 17948 21084 18004 21140
rect 19628 22764 19684 22820
rect 19871 22764 19927 22820
rect 20356 22764 20412 22820
rect 20748 22370 20804 22372
rect 20748 22318 20750 22370
rect 20750 22318 20802 22370
rect 20802 22318 20804 22370
rect 20748 22316 20804 22318
rect 21084 22316 21140 22372
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 18396 21756 18452 21812
rect 19292 21810 19348 21812
rect 19292 21758 19294 21810
rect 19294 21758 19346 21810
rect 19346 21758 19348 21810
rect 19292 21756 19348 21758
rect 19628 21756 19684 21812
rect 15820 20130 15876 20132
rect 15820 20078 15822 20130
rect 15822 20078 15874 20130
rect 15874 20078 15876 20130
rect 15820 20076 15876 20078
rect 15708 19292 15764 19348
rect 15372 17836 15428 17892
rect 14476 17052 14532 17108
rect 15988 19628 16044 19684
rect 14344 16098 14400 16100
rect 14344 16046 14346 16098
rect 14346 16046 14398 16098
rect 14398 16046 14400 16098
rect 14344 16044 14400 16046
rect 15932 18956 15988 19012
rect 16734 20018 16790 20020
rect 16734 19966 16736 20018
rect 16736 19966 16788 20018
rect 16788 19966 16790 20018
rect 16734 19964 16790 19966
rect 17276 20018 17332 20020
rect 17276 19966 17278 20018
rect 17278 19966 17330 20018
rect 17330 19966 17332 20018
rect 17276 19964 17332 19966
rect 16492 18956 16548 19012
rect 17108 19010 17164 19012
rect 17108 18958 17110 19010
rect 17110 18958 17162 19010
rect 17162 18958 17164 19010
rect 17108 18956 17164 18958
rect 14812 15314 14868 15316
rect 14812 15262 14814 15314
rect 14814 15262 14866 15314
rect 14866 15262 14868 15314
rect 17724 18060 17780 18116
rect 17724 16882 17780 16884
rect 17724 16830 17726 16882
rect 17726 16830 17778 16882
rect 17778 16830 17780 16882
rect 17724 16828 17780 16830
rect 14812 15260 14868 15262
rect 13692 14924 13748 14980
rect 16492 15260 16548 15316
rect 13468 14812 13524 14868
rect 13468 14530 13524 14532
rect 13468 14478 13470 14530
rect 13470 14478 13522 14530
rect 13522 14478 13524 14530
rect 13468 14476 13524 14478
rect 14588 14924 14644 14980
rect 16156 15036 16212 15092
rect 14344 14364 14400 14420
rect 13244 13692 13300 13748
rect 13804 13692 13860 13748
rect 13468 13244 13524 13300
rect 15596 14530 15652 14532
rect 15596 14478 15598 14530
rect 15598 14478 15650 14530
rect 15650 14478 15652 14530
rect 15596 14476 15652 14478
rect 15932 14588 15988 14644
rect 16044 14530 16100 14532
rect 16044 14478 16046 14530
rect 16046 14478 16098 14530
rect 16098 14478 16100 14530
rect 16044 14476 16100 14478
rect 15708 14252 15764 14308
rect 16044 13692 16100 13748
rect 17164 14252 17220 14308
rect 14476 13356 14532 13412
rect 16660 13468 16716 13524
rect 17052 13692 17108 13748
rect 17276 13746 17332 13748
rect 17276 13694 17278 13746
rect 17278 13694 17330 13746
rect 17330 13694 17332 13746
rect 17276 13692 17332 13694
rect 16156 12178 16212 12180
rect 16156 12126 16158 12178
rect 16158 12126 16210 12178
rect 16210 12126 16212 12178
rect 16156 12124 16212 12126
rect 17612 12124 17668 12180
rect 18508 20524 18564 20580
rect 18396 20076 18452 20132
rect 19012 21308 19068 21364
rect 19180 20188 19236 20244
rect 19292 20524 19348 20580
rect 18900 18060 18956 18116
rect 18172 17612 18228 17668
rect 18508 17666 18564 17668
rect 18508 17614 18510 17666
rect 18510 17614 18562 17666
rect 18562 17614 18564 17666
rect 18508 17612 18564 17614
rect 18060 16098 18116 16100
rect 18060 16046 18062 16098
rect 18062 16046 18114 16098
rect 18114 16046 18116 16098
rect 18060 16044 18116 16046
rect 18956 16828 19012 16884
rect 18228 15484 18284 15540
rect 18732 15484 18788 15540
rect 18396 15314 18452 15316
rect 18396 15262 18398 15314
rect 18398 15262 18450 15314
rect 18450 15262 18452 15314
rect 18396 15260 18452 15262
rect 18060 15148 18116 15204
rect 18172 15036 18228 15092
rect 18844 15202 18900 15204
rect 18844 15150 18846 15202
rect 18846 15150 18898 15202
rect 18898 15150 18900 15202
rect 18844 15148 18900 15150
rect 19180 16828 19236 16884
rect 18956 14924 19012 14980
rect 19404 17666 19460 17668
rect 19404 17614 19406 17666
rect 19406 17614 19458 17666
rect 19458 17614 19460 17666
rect 19404 17612 19460 17614
rect 21308 21532 21364 21588
rect 20207 20972 20263 21028
rect 20860 20860 20916 20916
rect 19684 20578 19740 20580
rect 19684 20526 19686 20578
rect 19686 20526 19738 20578
rect 19738 20526 19740 20578
rect 19684 20524 19740 20526
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19964 20188 20020 20244
rect 20524 20188 20580 20244
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19852 18508 19908 18564
rect 19292 15148 19348 15204
rect 21402 20914 21458 20916
rect 21402 20862 21404 20914
rect 21404 20862 21456 20914
rect 21456 20862 21458 20914
rect 21402 20860 21458 20862
rect 21756 23154 21812 23156
rect 21756 23102 21758 23154
rect 21758 23102 21810 23154
rect 21810 23102 21812 23154
rect 21756 23100 21812 23102
rect 21644 22316 21700 22372
rect 22652 23548 22708 23604
rect 21868 21196 21924 21252
rect 21644 20860 21700 20916
rect 21756 20748 21812 20804
rect 21476 19234 21532 19236
rect 21476 19182 21478 19234
rect 21478 19182 21530 19234
rect 21530 19182 21532 19234
rect 21476 19180 21532 19182
rect 21308 19122 21364 19124
rect 21308 19070 21310 19122
rect 21310 19070 21362 19122
rect 21362 19070 21364 19122
rect 21308 19068 21364 19070
rect 19628 18060 19684 18116
rect 19516 15372 19572 15428
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19852 17052 19908 17108
rect 19740 16882 19796 16884
rect 19740 16830 19742 16882
rect 19742 16830 19794 16882
rect 19794 16830 19796 16882
rect 19740 16828 19796 16830
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19852 15260 19908 15316
rect 19516 14924 19572 14980
rect 19628 14364 19684 14420
rect 20020 14364 20076 14420
rect 20300 14252 20356 14308
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 14028 11116 14084 11172
rect 16716 10610 16772 10612
rect 16716 10558 16718 10610
rect 16718 10558 16770 10610
rect 16770 10558 16772 10610
rect 16716 10556 16772 10558
rect 14812 10498 14868 10500
rect 14812 10446 14814 10498
rect 14814 10446 14866 10498
rect 14866 10446 14868 10498
rect 14812 10444 14868 10446
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 17108 11170 17164 11172
rect 17108 11118 17110 11170
rect 17110 11118 17162 11170
rect 17162 11118 17164 11170
rect 17108 11116 17164 11118
rect 21532 17724 21588 17780
rect 22148 21196 22204 21252
rect 22820 20914 22876 20916
rect 22820 20862 22822 20914
rect 22822 20862 22874 20914
rect 22874 20862 22876 20914
rect 22820 20860 22876 20862
rect 21756 19180 21812 19236
rect 21980 19292 22036 19348
rect 22204 19068 22260 19124
rect 23492 19740 23548 19796
rect 22820 19346 22876 19348
rect 22820 19294 22822 19346
rect 22822 19294 22874 19346
rect 22874 19294 22876 19346
rect 22820 19292 22876 19294
rect 23884 26684 23940 26740
rect 23772 26236 23828 26292
rect 23996 24444 24052 24500
rect 24444 28588 24500 28644
rect 24724 27858 24780 27860
rect 24724 27806 24726 27858
rect 24726 27806 24778 27858
rect 24778 27806 24780 27858
rect 24724 27804 24780 27806
rect 25564 28812 25620 28868
rect 25116 27356 25172 27412
rect 25564 27916 25620 27972
rect 25564 27468 25620 27524
rect 25676 27356 25732 27412
rect 26012 26908 26068 26964
rect 24444 23996 24500 24052
rect 24220 23436 24276 23492
rect 23772 22540 23828 22596
rect 24444 22594 24500 22596
rect 24444 22542 24446 22594
rect 24446 22542 24498 22594
rect 24498 22542 24500 22594
rect 24444 22540 24500 22542
rect 24556 21756 24612 21812
rect 24108 21586 24164 21588
rect 24108 21534 24110 21586
rect 24110 21534 24162 21586
rect 24162 21534 24164 21586
rect 24108 21532 24164 21534
rect 24332 21586 24388 21588
rect 24332 21534 24334 21586
rect 24334 21534 24386 21586
rect 24386 21534 24388 21586
rect 24332 21532 24388 21534
rect 25116 26796 25172 26852
rect 27132 30882 27188 30884
rect 27132 30830 27134 30882
rect 27134 30830 27186 30882
rect 27186 30830 27188 30882
rect 27132 30828 27188 30830
rect 26796 30156 26852 30212
rect 28252 34188 28308 34244
rect 28476 33404 28532 33460
rect 28028 31500 28084 31556
rect 27468 30994 27524 30996
rect 27468 30942 27470 30994
rect 27470 30942 27522 30994
rect 27522 30942 27524 30994
rect 27468 30940 27524 30942
rect 26572 30044 26628 30100
rect 28588 33292 28644 33348
rect 29484 33307 29540 33348
rect 29484 33292 29486 33307
rect 29486 33292 29538 33307
rect 29538 33292 29540 33307
rect 30044 33346 30100 33348
rect 30044 33294 30046 33346
rect 30046 33294 30098 33346
rect 30098 33294 30100 33346
rect 30044 33292 30100 33294
rect 29260 33068 29316 33124
rect 28364 32562 28420 32564
rect 28364 32510 28366 32562
rect 28366 32510 28418 32562
rect 28418 32510 28420 32562
rect 28364 32508 28420 32510
rect 28588 32508 28644 32564
rect 28140 31052 28196 31108
rect 27916 30716 27972 30772
rect 28476 30994 28532 30996
rect 28476 30942 28478 30994
rect 28478 30942 28530 30994
rect 28530 30942 28532 30994
rect 28476 30940 28532 30942
rect 29036 32562 29092 32564
rect 29036 32510 29038 32562
rect 29038 32510 29090 32562
rect 29090 32510 29092 32562
rect 29036 32508 29092 32510
rect 28868 32396 28924 32452
rect 31444 38722 31500 38724
rect 31444 38670 31446 38722
rect 31446 38670 31498 38722
rect 31498 38670 31500 38722
rect 31444 38668 31500 38670
rect 31948 38834 32004 38836
rect 31948 38782 31950 38834
rect 31950 38782 32002 38834
rect 32002 38782 32004 38834
rect 31948 38780 32004 38782
rect 33124 38834 33180 38836
rect 33124 38782 33126 38834
rect 33126 38782 33178 38834
rect 33178 38782 33180 38834
rect 33124 38780 33180 38782
rect 32060 38668 32116 38724
rect 30828 38108 30884 38164
rect 31836 38162 31892 38164
rect 31836 38110 31838 38162
rect 31838 38110 31890 38162
rect 31890 38110 31892 38162
rect 31836 38108 31892 38110
rect 31052 37660 31108 37716
rect 30828 37212 30884 37268
rect 30716 37100 30772 37156
rect 30548 36482 30604 36484
rect 30548 36430 30550 36482
rect 30550 36430 30602 36482
rect 30602 36430 30604 36482
rect 30548 36428 30604 36430
rect 32172 37436 32228 37492
rect 33180 37548 33236 37604
rect 31500 37100 31556 37156
rect 31052 36482 31108 36484
rect 31052 36430 31054 36482
rect 31054 36430 31106 36482
rect 31106 36430 31108 36482
rect 31052 36428 31108 36430
rect 31668 36482 31724 36484
rect 31668 36430 31670 36482
rect 31670 36430 31722 36482
rect 31722 36430 31724 36482
rect 31668 36428 31724 36430
rect 32340 37042 32396 37044
rect 32340 36990 32342 37042
rect 32342 36990 32394 37042
rect 32394 36990 32396 37042
rect 32340 36988 32396 36990
rect 33068 36876 33124 36932
rect 32956 36092 33012 36148
rect 32172 35868 32228 35924
rect 31836 35756 31892 35812
rect 30716 35644 30772 35700
rect 31052 35532 31108 35588
rect 31500 35586 31556 35588
rect 31500 35534 31502 35586
rect 31502 35534 31554 35586
rect 31554 35534 31556 35586
rect 31500 35532 31556 35534
rect 32060 35698 32116 35700
rect 32060 35646 32062 35698
rect 32062 35646 32114 35698
rect 32114 35646 32116 35698
rect 32060 35644 32116 35646
rect 33068 35756 33124 35812
rect 32396 35698 32452 35700
rect 32396 35646 32398 35698
rect 32398 35646 32450 35698
rect 32450 35646 32452 35698
rect 32396 35644 32452 35646
rect 33628 39004 33684 39060
rect 33404 38220 33460 38276
rect 34188 38220 34244 38276
rect 34524 39618 34580 39620
rect 34524 39566 34526 39618
rect 34526 39566 34578 39618
rect 34578 39566 34580 39618
rect 34524 39564 34580 39566
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 34972 39564 35028 39620
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35756 40460 35812 40516
rect 36092 40908 36148 40964
rect 35084 38780 35140 38836
rect 33628 37772 33684 37828
rect 33516 37266 33572 37268
rect 33516 37214 33518 37266
rect 33518 37214 33570 37266
rect 33570 37214 33572 37266
rect 33516 37212 33572 37214
rect 33180 36764 33236 36820
rect 34636 37884 34692 37940
rect 34860 37548 34916 37604
rect 33852 36988 33908 37044
rect 34300 36988 34356 37044
rect 33740 36652 33796 36708
rect 34860 36652 34916 36708
rect 34300 36540 34356 36596
rect 33516 36316 33572 36372
rect 33852 36204 33908 36260
rect 32172 35532 32228 35588
rect 33460 35586 33516 35588
rect 32396 35420 32452 35476
rect 33460 35534 33462 35586
rect 33462 35534 33514 35586
rect 33514 35534 33516 35586
rect 33460 35532 33516 35534
rect 34524 36540 34580 36596
rect 35420 38834 35476 38836
rect 35420 38782 35422 38834
rect 35422 38782 35474 38834
rect 35474 38782 35476 38834
rect 35420 38780 35476 38782
rect 36428 41186 36484 41188
rect 36428 41134 36430 41186
rect 36430 41134 36482 41186
rect 36482 41134 36484 41186
rect 36428 41132 36484 41134
rect 36540 40684 36596 40740
rect 36204 40572 36260 40628
rect 36876 40572 36932 40628
rect 37100 41132 37156 41188
rect 36316 39618 36372 39620
rect 36316 39566 36318 39618
rect 36318 39566 36370 39618
rect 36370 39566 36372 39618
rect 36316 39564 36372 39566
rect 36988 39618 37044 39620
rect 36988 39566 36990 39618
rect 36990 39566 37042 39618
rect 37042 39566 37044 39618
rect 36988 39564 37044 39566
rect 37772 41132 37828 41188
rect 37996 40962 38052 40964
rect 37996 40910 37998 40962
rect 37998 40910 38050 40962
rect 38050 40910 38052 40962
rect 37996 40908 38052 40910
rect 39788 41020 39844 41076
rect 37660 40348 37716 40404
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 36540 38050 36596 38052
rect 36540 37998 36542 38050
rect 36542 37998 36594 38050
rect 36594 37998 36596 38050
rect 36540 37996 36596 37998
rect 38612 40402 38668 40404
rect 38612 40350 38614 40402
rect 38614 40350 38666 40402
rect 38666 40350 38668 40402
rect 38612 40348 38668 40350
rect 40516 41074 40572 41076
rect 40516 41022 40518 41074
rect 40518 41022 40570 41074
rect 40570 41022 40572 41074
rect 40516 41020 40572 41022
rect 39900 40348 39956 40404
rect 39452 39676 39508 39732
rect 40124 40290 40180 40292
rect 40124 40238 40126 40290
rect 40126 40238 40178 40290
rect 40178 40238 40180 40290
rect 40124 40236 40180 40238
rect 39564 39590 39620 39620
rect 39452 39004 39508 39060
rect 39564 39564 39566 39590
rect 39566 39564 39618 39590
rect 39618 39564 39620 39590
rect 39452 38817 39454 38836
rect 39454 38817 39506 38836
rect 39506 38817 39508 38836
rect 39452 38780 39508 38817
rect 39340 38556 39396 38612
rect 37436 38050 37492 38052
rect 37436 37998 37438 38050
rect 37438 37998 37490 38050
rect 37490 37998 37492 38050
rect 37436 37996 37492 37998
rect 38668 38050 38724 38052
rect 38668 37998 38670 38050
rect 38670 37998 38722 38050
rect 38722 37998 38724 38050
rect 38668 37996 38724 37998
rect 37100 37938 37156 37940
rect 37100 37886 37102 37938
rect 37102 37886 37154 37938
rect 37154 37886 37156 37938
rect 37100 37884 37156 37886
rect 35868 37772 35924 37828
rect 36372 37826 36428 37828
rect 36372 37774 36374 37826
rect 36374 37774 36426 37826
rect 36426 37774 36428 37826
rect 36372 37772 36428 37774
rect 35868 37266 35924 37268
rect 35868 37214 35870 37266
rect 35870 37214 35922 37266
rect 35922 37214 35924 37266
rect 35868 37212 35924 37214
rect 35532 36988 35588 37044
rect 36540 37212 36596 37268
rect 36204 37154 36260 37156
rect 36204 37102 36206 37154
rect 36206 37102 36258 37154
rect 36258 37102 36260 37154
rect 36204 37100 36260 37102
rect 36092 36988 36148 37044
rect 37212 37100 37268 37156
rect 37436 37212 37492 37268
rect 36652 36988 36708 37044
rect 36988 36988 37044 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35084 36540 35140 36596
rect 34412 36204 34468 36260
rect 34412 35868 34468 35924
rect 33964 35532 34020 35588
rect 34132 35420 34188 35476
rect 30380 34188 30436 34244
rect 30492 34636 30548 34692
rect 31220 34690 31276 34692
rect 31220 34638 31222 34690
rect 31222 34638 31274 34690
rect 31274 34638 31276 34690
rect 31220 34636 31276 34638
rect 31948 34636 32004 34692
rect 33068 34860 33124 34916
rect 32172 34188 32228 34244
rect 31500 33404 31556 33460
rect 31276 33346 31332 33348
rect 31276 33294 31278 33346
rect 31278 33294 31330 33346
rect 31330 33294 31332 33346
rect 31276 33292 31332 33294
rect 30492 32284 30548 32340
rect 30604 32562 30660 32564
rect 30604 32510 30606 32562
rect 30606 32510 30658 32562
rect 30658 32510 30660 32562
rect 30604 32508 30660 32510
rect 31052 32620 31108 32676
rect 30604 32172 30660 32228
rect 29652 31836 29708 31892
rect 29484 31778 29540 31780
rect 29484 31726 29486 31778
rect 29486 31726 29538 31778
rect 29538 31726 29540 31778
rect 29484 31724 29540 31726
rect 29372 31500 29428 31556
rect 28980 31164 29036 31220
rect 29596 31106 29652 31108
rect 29596 31054 29598 31106
rect 29598 31054 29650 31106
rect 29650 31054 29652 31106
rect 29596 31052 29652 31054
rect 28084 30434 28140 30436
rect 28084 30382 28086 30434
rect 28086 30382 28138 30434
rect 28138 30382 28140 30434
rect 28084 30380 28140 30382
rect 27244 30175 27300 30212
rect 27244 30156 27246 30175
rect 27246 30156 27298 30175
rect 27298 30156 27300 30175
rect 26796 28627 26852 28644
rect 26796 28588 26798 28627
rect 26798 28588 26850 28627
rect 26850 28588 26852 28627
rect 27580 28627 27636 28644
rect 27580 28588 27582 28627
rect 27582 28588 27634 28627
rect 27634 28588 27636 28627
rect 26460 28364 26516 28420
rect 26348 27468 26404 27524
rect 26348 27074 26404 27076
rect 26348 27022 26350 27074
rect 26350 27022 26402 27074
rect 26402 27022 26404 27074
rect 26348 27020 26404 27022
rect 24780 25228 24836 25284
rect 25564 25228 25620 25284
rect 26124 25228 26180 25284
rect 25900 25116 25956 25172
rect 25340 24050 25396 24052
rect 25340 23998 25342 24050
rect 25342 23998 25394 24050
rect 25394 23998 25396 24050
rect 25340 23996 25396 23998
rect 27356 28364 27412 28420
rect 26572 27468 26628 27524
rect 27244 27468 27300 27524
rect 26684 27356 26740 27412
rect 26572 26908 26628 26964
rect 27020 27020 27076 27076
rect 27356 27244 27412 27300
rect 26460 24498 26516 24500
rect 26460 24446 26462 24498
rect 26462 24446 26514 24498
rect 26514 24446 26516 24498
rect 26460 24444 26516 24446
rect 25452 23548 25508 23604
rect 27468 25452 27524 25508
rect 26908 23660 26964 23716
rect 25900 23042 25956 23044
rect 25900 22990 25902 23042
rect 25902 22990 25954 23042
rect 25954 22990 25956 23042
rect 25900 22988 25956 22990
rect 25452 22540 25508 22596
rect 26684 22370 26740 22372
rect 26348 21868 26404 21924
rect 26684 22318 26686 22370
rect 26686 22318 26738 22370
rect 26738 22318 26740 22370
rect 26684 22316 26740 22318
rect 26460 21532 26516 21588
rect 25228 21420 25284 21476
rect 25116 20802 25172 20804
rect 25116 20750 25118 20802
rect 25118 20750 25170 20802
rect 25170 20750 25172 20802
rect 25116 20748 25172 20750
rect 23660 19628 23716 19684
rect 24276 20018 24332 20020
rect 24276 19966 24278 20018
rect 24278 19966 24330 20018
rect 24330 19966 24332 20018
rect 24276 19964 24332 19966
rect 22540 18508 22596 18564
rect 23996 19740 24052 19796
rect 22876 18450 22932 18452
rect 22204 17948 22260 18004
rect 20860 17666 20916 17668
rect 20860 17614 20862 17666
rect 20862 17614 20914 17666
rect 20914 17614 20916 17666
rect 20860 17612 20916 17614
rect 22876 18398 22878 18450
rect 22878 18398 22930 18450
rect 22930 18398 22932 18450
rect 22876 18396 22932 18398
rect 24724 19740 24780 19796
rect 24220 19628 24276 19684
rect 23996 18450 24052 18452
rect 23996 18398 23998 18450
rect 23998 18398 24050 18450
rect 24050 18398 24052 18450
rect 23996 18396 24052 18398
rect 22204 17500 22260 17556
rect 21532 17052 21588 17108
rect 23118 17612 23174 17668
rect 22428 17388 22484 17444
rect 24108 19292 24164 19348
rect 23754 18338 23810 18340
rect 23754 18286 23756 18338
rect 23756 18286 23808 18338
rect 23808 18286 23810 18338
rect 23754 18284 23810 18286
rect 23660 17724 23716 17780
rect 23100 16156 23156 16212
rect 22876 16098 22932 16100
rect 22876 16046 22878 16098
rect 22878 16046 22930 16098
rect 22930 16046 22932 16098
rect 22876 16044 22932 16046
rect 24108 17666 24164 17668
rect 24108 17614 24110 17666
rect 24110 17614 24162 17666
rect 24162 17614 24164 17666
rect 24108 17612 24164 17614
rect 23996 16882 24052 16884
rect 23996 16830 23998 16882
rect 23998 16830 24050 16882
rect 24050 16830 24052 16882
rect 23996 16828 24052 16830
rect 25396 21026 25452 21028
rect 25396 20974 25398 21026
rect 25398 20974 25450 21026
rect 25450 20974 25452 21026
rect 25396 20972 25452 20974
rect 26684 20860 26740 20916
rect 26796 21868 26852 21924
rect 27468 25116 27524 25172
rect 27244 23826 27300 23828
rect 27244 23774 27246 23826
rect 27246 23774 27298 23826
rect 27298 23774 27300 23826
rect 27244 23772 27300 23774
rect 27468 22764 27524 22820
rect 26348 20412 26404 20468
rect 24500 18172 24556 18228
rect 24332 17836 24388 17892
rect 24444 17948 24500 18004
rect 24556 17724 24612 17780
rect 24500 17052 24556 17108
rect 24780 18396 24836 18452
rect 25452 18450 25508 18452
rect 25452 18398 25454 18450
rect 25454 18398 25506 18450
rect 25506 18398 25508 18450
rect 25452 18396 25508 18398
rect 25116 18284 25172 18340
rect 25452 17836 25508 17892
rect 24220 16716 24276 16772
rect 24668 16492 24724 16548
rect 23884 16268 23940 16324
rect 24892 16268 24948 16324
rect 23660 16210 23716 16212
rect 23660 16158 23662 16210
rect 23662 16158 23714 16210
rect 23714 16158 23716 16210
rect 23660 16156 23716 16158
rect 23324 16044 23380 16100
rect 23772 15484 23828 15540
rect 24276 15538 24332 15540
rect 24276 15486 24278 15538
rect 24278 15486 24330 15538
rect 24330 15486 24332 15538
rect 24276 15484 24332 15486
rect 21756 15314 21812 15316
rect 21756 15262 21758 15314
rect 21758 15262 21810 15314
rect 21810 15262 21812 15314
rect 21756 15260 21812 15262
rect 21196 14588 21252 14644
rect 23100 15148 23156 15204
rect 21420 14588 21476 14644
rect 21308 13916 21364 13972
rect 20748 12348 20804 12404
rect 18620 11564 18676 11620
rect 18396 11452 18452 11508
rect 19852 11564 19908 11620
rect 21868 13692 21924 13748
rect 24444 15148 24500 15204
rect 22988 14924 23044 14980
rect 22652 14306 22708 14308
rect 22652 14254 22654 14306
rect 22654 14254 22706 14306
rect 22706 14254 22708 14306
rect 22652 14252 22708 14254
rect 23100 13916 23156 13972
rect 23212 13634 23268 13636
rect 23212 13582 23214 13634
rect 23214 13582 23266 13634
rect 23266 13582 23268 13634
rect 23212 13580 23268 13582
rect 25452 17052 25508 17108
rect 25340 16828 25396 16884
rect 27356 20748 27412 20804
rect 26348 20018 26404 20020
rect 26348 19966 26350 20018
rect 26350 19966 26402 20018
rect 26402 19966 26404 20018
rect 26348 19964 26404 19966
rect 27020 19964 27076 20020
rect 27132 20076 27188 20132
rect 28028 28252 28084 28308
rect 27804 27132 27860 27188
rect 29260 30994 29316 30996
rect 29260 30942 29262 30994
rect 29262 30942 29314 30994
rect 29314 30942 29316 30994
rect 29260 30940 29316 30942
rect 30268 31612 30324 31668
rect 31276 31724 31332 31780
rect 31948 33292 32004 33348
rect 34300 34914 34356 34916
rect 34300 34862 34302 34914
rect 34302 34862 34354 34914
rect 34354 34862 34356 34914
rect 34300 34860 34356 34862
rect 33516 34111 33518 34132
rect 33518 34111 33570 34132
rect 33570 34111 33572 34132
rect 33516 34076 33572 34111
rect 32396 33516 32452 33572
rect 32284 33404 32340 33460
rect 31836 32620 31892 32676
rect 31724 32562 31780 32564
rect 31724 32510 31726 32562
rect 31726 32510 31778 32562
rect 31778 32510 31780 32562
rect 31724 32508 31780 32510
rect 31982 32284 32038 32340
rect 31144 31164 31200 31220
rect 30492 31052 30548 31108
rect 30156 30828 30212 30884
rect 28812 28588 28868 28644
rect 29820 28476 29876 28532
rect 29148 28364 29204 28420
rect 28700 27244 28756 27300
rect 30268 28252 30324 28308
rect 29652 27132 29708 27188
rect 30268 27186 30324 27188
rect 30268 27134 30270 27186
rect 30270 27134 30322 27186
rect 30322 27134 30324 27186
rect 30268 27132 30324 27134
rect 29148 26908 29204 26964
rect 28588 26460 28644 26516
rect 29708 26908 29764 26964
rect 29372 26012 29428 26068
rect 27804 25506 27860 25508
rect 27804 25454 27806 25506
rect 27806 25454 27858 25506
rect 27858 25454 27860 25506
rect 27804 25452 27860 25454
rect 28476 25228 28532 25284
rect 27692 23772 27748 23828
rect 27692 22764 27748 22820
rect 28308 22988 28364 23044
rect 28364 21868 28420 21924
rect 28644 24834 28700 24836
rect 28644 24782 28646 24834
rect 28646 24782 28698 24834
rect 28698 24782 28700 24834
rect 28644 24780 28700 24782
rect 29148 24444 29204 24500
rect 28700 23996 28756 24052
rect 29484 26460 29540 26516
rect 29260 23996 29316 24052
rect 29764 25394 29820 25396
rect 29764 25342 29766 25394
rect 29766 25342 29818 25394
rect 29818 25342 29820 25394
rect 29764 25340 29820 25342
rect 29148 23660 29204 23716
rect 28812 23324 28868 23380
rect 28812 22876 28868 22932
rect 28588 22316 28644 22372
rect 28700 21644 28756 21700
rect 27692 20802 27748 20804
rect 27692 20750 27694 20802
rect 27694 20750 27746 20802
rect 27746 20750 27748 20802
rect 27692 20748 27748 20750
rect 27468 20412 27524 20468
rect 28644 20412 28700 20468
rect 28028 20076 28084 20132
rect 25788 18284 25844 18340
rect 25788 17724 25844 17780
rect 26012 17836 26068 17892
rect 26012 16882 26068 16884
rect 26012 16830 26014 16882
rect 26014 16830 26066 16882
rect 26066 16830 26068 16882
rect 26012 16828 26068 16830
rect 26124 17666 26180 17668
rect 26124 17614 26126 17666
rect 26126 17614 26178 17666
rect 26178 17614 26180 17666
rect 26124 17612 26180 17614
rect 25900 15484 25956 15540
rect 23996 13746 24052 13748
rect 23996 13694 23998 13746
rect 23998 13694 24050 13746
rect 24050 13694 24052 13746
rect 23996 13692 24052 13694
rect 24948 13916 25004 13972
rect 24444 13634 24500 13636
rect 24444 13582 24446 13634
rect 24446 13582 24498 13634
rect 24498 13582 24500 13634
rect 24444 13580 24500 13582
rect 20636 11506 20692 11508
rect 20636 11454 20638 11506
rect 20638 11454 20690 11506
rect 20690 11454 20692 11506
rect 20636 11452 20692 11454
rect 18060 11116 18116 11172
rect 17388 10498 17444 10500
rect 17388 10446 17390 10498
rect 17390 10446 17442 10498
rect 17442 10446 17444 10498
rect 17388 10444 17444 10446
rect 17836 10610 17892 10612
rect 17836 10558 17838 10610
rect 17838 10558 17890 10610
rect 17890 10558 17892 10610
rect 17836 10556 17892 10558
rect 16940 9548 16996 9604
rect 16324 8988 16380 9044
rect 16492 8876 16548 8932
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 17948 9996 18004 10052
rect 18620 9772 18676 9828
rect 18732 9996 18788 10052
rect 17836 9548 17892 9604
rect 17948 9100 18004 9156
rect 17780 8818 17836 8820
rect 17780 8766 17782 8818
rect 17782 8766 17834 8818
rect 17834 8766 17836 8818
rect 17780 8764 17836 8766
rect 18620 8876 18676 8932
rect 18620 8652 18676 8708
rect 16940 7474 16996 7476
rect 16940 7422 16942 7474
rect 16942 7422 16994 7474
rect 16994 7422 16996 7474
rect 18956 9212 19012 9268
rect 19292 9660 19348 9716
rect 19292 9100 19348 9156
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19740 9938 19796 9940
rect 19740 9886 19742 9938
rect 19742 9886 19794 9938
rect 19794 9886 19796 9938
rect 19740 9884 19796 9886
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 18844 9042 18900 9044
rect 18844 8990 18846 9042
rect 18846 8990 18898 9042
rect 18898 8990 18900 9042
rect 18844 8988 18900 8990
rect 16940 7420 16996 7422
rect 17724 7420 17780 7476
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 15148 5852 15204 5908
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 16492 5906 16548 5908
rect 16492 5854 16494 5906
rect 16494 5854 16546 5906
rect 16546 5854 16548 5906
rect 16492 5852 16548 5854
rect 16940 5964 16996 6020
rect 16604 5740 16660 5796
rect 16772 5682 16828 5684
rect 16772 5630 16774 5682
rect 16774 5630 16826 5682
rect 16826 5630 16828 5682
rect 16772 5628 16828 5630
rect 17724 6076 17780 6132
rect 17612 5964 17668 6020
rect 17388 5794 17444 5796
rect 17388 5742 17390 5794
rect 17390 5742 17442 5794
rect 17442 5742 17444 5794
rect 17388 5740 17444 5742
rect 17500 4956 17556 5012
rect 19740 8876 19796 8932
rect 19180 8652 19236 8708
rect 19068 8316 19124 8372
rect 18844 7868 18900 7924
rect 20076 8652 20132 8708
rect 22316 11618 22372 11620
rect 22316 11566 22318 11618
rect 22318 11566 22370 11618
rect 22370 11566 22372 11618
rect 22316 11564 22372 11566
rect 22428 11452 22484 11508
rect 23660 11788 23716 11844
rect 22652 10780 22708 10836
rect 21644 9884 21700 9940
rect 21308 9798 21364 9828
rect 21308 9772 21310 9798
rect 21310 9772 21362 9798
rect 21362 9772 21364 9798
rect 21196 8652 21252 8708
rect 18956 7308 19012 7364
rect 18508 6860 18564 6916
rect 18620 6748 18676 6804
rect 18396 6076 18452 6132
rect 18620 6188 18676 6244
rect 17836 5852 17892 5908
rect 17836 5628 17892 5684
rect 18620 5794 18676 5796
rect 18620 5742 18622 5794
rect 18622 5742 18674 5794
rect 18674 5742 18676 5794
rect 18620 5740 18676 5742
rect 18284 5180 18340 5236
rect 18060 5068 18116 5124
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 17948 4301 17950 4340
rect 17950 4301 18002 4340
rect 18002 4301 18004 4340
rect 17948 4284 18004 4301
rect 18732 5122 18788 5124
rect 18732 5070 18734 5122
rect 18734 5070 18786 5122
rect 18786 5070 18788 5122
rect 18732 5068 18788 5070
rect 18284 4956 18340 5012
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 21532 8204 21588 8260
rect 19068 6636 19124 6692
rect 19292 6188 19348 6244
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19516 5852 19572 5908
rect 20636 6690 20692 6692
rect 20636 6638 20638 6690
rect 20638 6638 20690 6690
rect 20690 6638 20692 6690
rect 20636 6636 20692 6638
rect 20392 6524 20448 6580
rect 20636 5964 20692 6020
rect 20412 5794 20468 5796
rect 20412 5742 20414 5794
rect 20414 5742 20466 5794
rect 20466 5742 20468 5794
rect 20412 5740 20468 5742
rect 25788 15260 25844 15316
rect 25340 12738 25396 12740
rect 25340 12686 25342 12738
rect 25342 12686 25394 12738
rect 25394 12686 25396 12738
rect 25340 12684 25396 12686
rect 25228 12290 25284 12292
rect 25228 12238 25230 12290
rect 25230 12238 25282 12290
rect 25282 12238 25284 12290
rect 25228 12236 25284 12238
rect 24556 11788 24612 11844
rect 24780 11900 24836 11956
rect 24444 10834 24500 10836
rect 24444 10782 24446 10834
rect 24446 10782 24498 10834
rect 24498 10782 24500 10834
rect 24444 10780 24500 10782
rect 22316 10050 22372 10052
rect 22316 9998 22318 10050
rect 22318 9998 22370 10050
rect 22370 9998 22372 10050
rect 22316 9996 22372 9998
rect 23436 9884 23492 9940
rect 23324 9266 23380 9268
rect 23324 9214 23326 9266
rect 23326 9214 23378 9266
rect 23378 9214 23380 9266
rect 23324 9212 23380 9214
rect 23324 8092 23380 8148
rect 21756 7362 21812 7364
rect 21756 7310 21758 7362
rect 21758 7310 21810 7362
rect 21810 7310 21812 7362
rect 21756 7308 21812 7310
rect 22316 7474 22372 7476
rect 22316 7422 22318 7474
rect 22318 7422 22370 7474
rect 22370 7422 22372 7474
rect 22316 7420 22372 7422
rect 22316 6914 22372 6916
rect 22316 6862 22318 6914
rect 22318 6862 22370 6914
rect 22370 6862 22372 6914
rect 22316 6860 22372 6862
rect 22092 6748 22148 6804
rect 22316 5852 22372 5908
rect 24556 10220 24612 10276
rect 25396 11788 25452 11844
rect 25340 11564 25396 11620
rect 24780 10108 24836 10164
rect 24108 9660 24164 9716
rect 25452 9996 25508 10052
rect 24780 8428 24836 8484
rect 23660 6524 23716 6580
rect 23996 8204 24052 8260
rect 24220 8204 24276 8260
rect 24984 8258 25040 8260
rect 24984 8206 24986 8258
rect 24986 8206 25038 8258
rect 25038 8206 25040 8258
rect 24984 8204 25040 8206
rect 24444 6663 24500 6692
rect 24444 6636 24446 6663
rect 24446 6636 24498 6663
rect 24498 6636 24500 6663
rect 24108 6524 24164 6580
rect 24444 6412 24500 6468
rect 23436 5906 23492 5908
rect 23436 5854 23438 5906
rect 23438 5854 23490 5906
rect 23490 5854 23492 5906
rect 23436 5852 23492 5854
rect 20188 4956 20244 5012
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 17500 3554 17556 3556
rect 17500 3502 17502 3554
rect 17502 3502 17554 3554
rect 17554 3502 17556 3554
rect 17500 3500 17556 3502
rect 19516 4060 19572 4116
rect 19516 3500 19572 3556
rect 22316 5180 22372 5236
rect 21532 5122 21588 5124
rect 21532 5070 21534 5122
rect 21534 5070 21586 5122
rect 21586 5070 21588 5122
rect 21532 5068 21588 5070
rect 21756 5122 21812 5124
rect 21756 5070 21758 5122
rect 21758 5070 21810 5122
rect 21810 5070 21812 5122
rect 21756 5068 21812 5070
rect 21364 4898 21420 4900
rect 21364 4846 21366 4898
rect 21366 4846 21418 4898
rect 21418 4846 21420 4898
rect 21364 4844 21420 4846
rect 22204 4844 22260 4900
rect 22876 4508 22932 4564
rect 22540 4301 22542 4340
rect 22542 4301 22594 4340
rect 22594 4301 22596 4340
rect 22540 4284 22596 4301
rect 21420 4226 21476 4228
rect 21420 4174 21422 4226
rect 21422 4174 21474 4226
rect 21474 4174 21476 4226
rect 21420 4172 21476 4174
rect 22428 4226 22484 4228
rect 22428 4174 22430 4226
rect 22430 4174 22482 4226
rect 22482 4174 22484 4226
rect 22428 4172 22484 4174
rect 22876 4060 22932 4116
rect 22540 3724 22596 3780
rect 22988 3554 23044 3556
rect 22988 3502 22990 3554
rect 22990 3502 23042 3554
rect 23042 3502 23044 3554
rect 22988 3500 23044 3502
rect 26012 16604 26068 16660
rect 28140 19964 28196 20020
rect 26908 19180 26964 19236
rect 26572 18450 26628 18452
rect 26572 18398 26574 18450
rect 26574 18398 26626 18450
rect 26626 18398 26628 18450
rect 26572 18396 26628 18398
rect 26796 18338 26852 18340
rect 26796 18286 26798 18338
rect 26798 18286 26850 18338
rect 26850 18286 26852 18338
rect 26796 18284 26852 18286
rect 26460 18172 26516 18228
rect 27244 18172 27300 18228
rect 27356 18396 27412 18452
rect 26236 16604 26292 16660
rect 26572 18060 26628 18116
rect 27132 17948 27188 18004
rect 27020 17500 27076 17556
rect 26908 16882 26964 16884
rect 26908 16830 26910 16882
rect 26910 16830 26962 16882
rect 26962 16830 26964 16882
rect 26908 16828 26964 16830
rect 26908 16604 26964 16660
rect 26796 16098 26852 16100
rect 26796 16046 26798 16098
rect 26798 16046 26850 16098
rect 26850 16046 26852 16098
rect 26796 16044 26852 16046
rect 26908 16044 26964 16100
rect 27804 18284 27860 18340
rect 27580 18060 27636 18116
rect 28140 18844 28196 18900
rect 27916 17948 27972 18004
rect 27244 17052 27300 17108
rect 27465 16940 27521 16996
rect 27916 17052 27972 17108
rect 28364 19628 28420 19684
rect 28924 20076 28980 20132
rect 29372 23100 29428 23156
rect 29260 21868 29316 21924
rect 29540 22540 29596 22596
rect 32396 32060 32452 32116
rect 32956 32284 33012 32340
rect 30604 30828 30660 30884
rect 31108 30994 31164 30996
rect 31108 30942 31110 30994
rect 31110 30942 31162 30994
rect 31162 30942 31164 30994
rect 31724 31052 31780 31108
rect 31108 30940 31164 30942
rect 30828 30828 30884 30884
rect 31948 31724 32004 31780
rect 32172 31778 32228 31780
rect 32172 31726 32174 31778
rect 32174 31726 32226 31778
rect 32226 31726 32228 31778
rect 32172 31724 32228 31726
rect 33404 32284 33460 32340
rect 34692 35980 34748 36036
rect 34692 35810 34748 35812
rect 34692 35758 34694 35810
rect 34694 35758 34746 35810
rect 34746 35758 34748 35810
rect 34692 35756 34748 35758
rect 34972 35420 35028 35476
rect 35196 36316 35252 36372
rect 35476 35698 35532 35700
rect 35476 35646 35478 35698
rect 35478 35646 35530 35698
rect 35530 35646 35532 35698
rect 35476 35644 35532 35646
rect 35532 35420 35588 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34636 34076 34692 34132
rect 35924 35420 35980 35476
rect 35756 35084 35812 35140
rect 35084 33852 35140 33908
rect 37044 35474 37100 35476
rect 37044 35422 37046 35474
rect 37046 35422 37098 35474
rect 37098 35422 37100 35474
rect 37044 35420 37100 35422
rect 34020 32674 34076 32676
rect 34020 32622 34022 32674
rect 34022 32622 34074 32674
rect 34074 32622 34076 32674
rect 34020 32620 34076 32622
rect 33740 31836 33796 31892
rect 32732 31052 32788 31108
rect 31836 30828 31892 30884
rect 32172 30828 32228 30884
rect 32284 30940 32340 30996
rect 30828 30380 30884 30436
rect 31612 30210 31668 30212
rect 31612 30158 31614 30210
rect 31614 30158 31666 30210
rect 31666 30158 31668 30210
rect 31612 30156 31668 30158
rect 32732 30434 32788 30436
rect 32732 30382 32734 30434
rect 32734 30382 32786 30434
rect 32786 30382 32788 30434
rect 32732 30380 32788 30382
rect 33180 30994 33236 30996
rect 33180 30942 33182 30994
rect 33182 30942 33234 30994
rect 33234 30942 33236 30994
rect 33180 30940 33236 30942
rect 33348 30994 33404 30996
rect 33348 30942 33350 30994
rect 33350 30942 33402 30994
rect 33402 30942 33404 30994
rect 33348 30940 33404 30942
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35084 33516 35140 33572
rect 34412 33068 34468 33124
rect 34748 33180 34804 33236
rect 34580 32844 34636 32900
rect 34300 32284 34356 32340
rect 34300 32060 34356 32116
rect 33852 30940 33908 30996
rect 33740 30770 33796 30772
rect 33740 30718 33742 30770
rect 33742 30718 33794 30770
rect 33794 30718 33796 30770
rect 33740 30716 33796 30718
rect 33516 30380 33572 30436
rect 33068 30156 33124 30212
rect 34188 30994 34244 30996
rect 34188 30942 34190 30994
rect 34190 30942 34242 30994
rect 34242 30942 34244 30994
rect 34188 30940 34244 30942
rect 34972 33292 35028 33348
rect 35532 32620 35588 32676
rect 35644 32844 35700 32900
rect 35196 32396 35252 32452
rect 35644 32508 35700 32564
rect 34860 31836 34916 31892
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35868 32284 35924 32340
rect 35756 31948 35812 32004
rect 35308 31778 35364 31780
rect 35308 31726 35310 31778
rect 35310 31726 35362 31778
rect 35362 31726 35364 31778
rect 35308 31724 35364 31726
rect 35532 30940 35588 30996
rect 35644 31724 35700 31780
rect 36484 33122 36540 33124
rect 36484 33070 36486 33122
rect 36486 33070 36538 33122
rect 36538 33070 36540 33122
rect 36484 33068 36540 33070
rect 37100 35026 37156 35028
rect 37100 34974 37102 35026
rect 37102 34974 37154 35026
rect 37154 34974 37156 35026
rect 37100 34972 37156 34974
rect 37212 34300 37268 34356
rect 37324 34972 37380 35028
rect 36764 33516 36820 33572
rect 37212 34106 37214 34132
rect 37214 34106 37266 34132
rect 37266 34106 37268 34132
rect 37884 37266 37940 37268
rect 37884 37214 37886 37266
rect 37886 37214 37938 37266
rect 37938 37214 37940 37266
rect 37884 37212 37940 37214
rect 38220 37212 38276 37268
rect 37548 37042 37604 37044
rect 37548 36990 37550 37042
rect 37550 36990 37602 37042
rect 37602 36990 37604 37042
rect 37548 36988 37604 36990
rect 39228 37266 39284 37268
rect 39228 37214 39230 37266
rect 39230 37214 39282 37266
rect 39282 37214 39284 37266
rect 39228 37212 39284 37214
rect 39788 38556 39844 38612
rect 40012 40124 40068 40180
rect 40012 38668 40068 38724
rect 40292 38610 40348 38612
rect 40292 38558 40294 38610
rect 40294 38558 40346 38610
rect 40346 38558 40348 38610
rect 40292 38556 40348 38558
rect 39340 36988 39396 37044
rect 39900 36988 39956 37044
rect 37996 36594 38052 36596
rect 37996 36542 37998 36594
rect 37998 36542 38050 36594
rect 38050 36542 38052 36594
rect 37996 36540 38052 36542
rect 39788 36316 39844 36372
rect 37884 36092 37940 36148
rect 40012 35756 40068 35812
rect 39452 35586 39508 35588
rect 39452 35534 39454 35586
rect 39454 35534 39506 35586
rect 39506 35534 39508 35586
rect 39452 35532 39508 35534
rect 37884 34188 37940 34244
rect 37212 34076 37268 34106
rect 37436 34076 37492 34132
rect 36988 33404 37044 33460
rect 37324 33852 37380 33908
rect 37044 33234 37100 33236
rect 37044 33182 37046 33234
rect 37046 33182 37098 33234
rect 37098 33182 37100 33234
rect 37044 33180 37100 33182
rect 37548 33404 37604 33460
rect 38332 33628 38388 33684
rect 37884 33516 37940 33572
rect 38108 33346 38164 33348
rect 38108 33294 38110 33346
rect 38110 33294 38162 33346
rect 38162 33294 38164 33346
rect 38108 33292 38164 33294
rect 36652 32956 36708 33012
rect 35980 31836 36036 31892
rect 37996 32956 38052 33012
rect 39004 33628 39060 33684
rect 38892 33292 38948 33348
rect 39452 33346 39508 33348
rect 39452 33294 39454 33346
rect 39454 33294 39506 33346
rect 39506 33294 39508 33346
rect 39452 33292 39508 33294
rect 38836 32786 38892 32788
rect 38836 32734 38838 32786
rect 38838 32734 38890 32786
rect 38890 32734 38892 32786
rect 38836 32732 38892 32734
rect 39788 34076 39844 34132
rect 39788 33292 39844 33348
rect 41020 40348 41076 40404
rect 42028 40572 42084 40628
rect 42812 40572 42868 40628
rect 41580 40290 41636 40292
rect 41580 40238 41582 40290
rect 41582 40238 41634 40290
rect 41634 40238 41636 40290
rect 41580 40236 41636 40238
rect 41356 40124 41412 40180
rect 41356 39730 41412 39732
rect 41356 39678 41358 39730
rect 41358 39678 41410 39730
rect 41410 39678 41412 39730
rect 41356 39676 41412 39678
rect 41244 39564 41300 39620
rect 40908 39452 40964 39508
rect 40572 39340 40628 39396
rect 40908 38780 40964 38836
rect 41356 38780 41412 38836
rect 41020 38722 41076 38724
rect 41020 38670 41022 38722
rect 41022 38670 41074 38722
rect 41074 38670 41076 38722
rect 41020 38668 41076 38670
rect 41580 38668 41636 38724
rect 41916 38444 41972 38500
rect 41468 37212 41524 37268
rect 41692 37266 41748 37268
rect 41692 37214 41694 37266
rect 41694 37214 41746 37266
rect 41746 37214 41748 37266
rect 41692 37212 41748 37214
rect 40460 36652 40516 36708
rect 42028 36876 42084 36932
rect 40516 36370 40572 36372
rect 40516 36318 40518 36370
rect 40518 36318 40570 36370
rect 40570 36318 40572 36370
rect 40516 36316 40572 36318
rect 41020 36454 41076 36484
rect 41020 36428 41022 36454
rect 41022 36428 41074 36454
rect 41074 36428 41076 36454
rect 40908 35644 40964 35700
rect 42028 35980 42084 36036
rect 41580 35586 41636 35588
rect 41580 35534 41582 35586
rect 41582 35534 41634 35586
rect 41634 35534 41636 35586
rect 41580 35532 41636 35534
rect 41356 35196 41412 35252
rect 40236 34972 40292 35028
rect 40684 35026 40740 35028
rect 40684 34974 40686 35026
rect 40686 34974 40738 35026
rect 40738 34974 40740 35026
rect 40684 34972 40740 34974
rect 40124 34188 40180 34244
rect 38668 32562 38724 32564
rect 38668 32510 38670 32562
rect 38670 32510 38722 32562
rect 38722 32510 38724 32562
rect 40348 34748 40404 34804
rect 40236 32732 40292 32788
rect 42588 34802 42644 34804
rect 42588 34750 42590 34802
rect 42590 34750 42642 34802
rect 42642 34750 42644 34802
rect 42588 34748 42644 34750
rect 41580 34188 41636 34244
rect 40796 34130 40852 34132
rect 40796 34078 40798 34130
rect 40798 34078 40850 34130
rect 40850 34078 40852 34130
rect 40796 34076 40852 34078
rect 43036 39788 43092 39844
rect 43484 40124 43540 40180
rect 43932 39842 43988 39844
rect 43932 39790 43934 39842
rect 43934 39790 43986 39842
rect 43986 39790 43988 39842
rect 43932 39788 43988 39790
rect 43372 39676 43428 39732
rect 43260 39506 43316 39508
rect 43260 39454 43262 39506
rect 43262 39454 43314 39506
rect 43314 39454 43316 39506
rect 43260 39452 43316 39454
rect 42924 38220 42980 38276
rect 43372 38556 43428 38612
rect 43036 37212 43092 37268
rect 43148 36316 43204 36372
rect 43148 35868 43204 35924
rect 43708 38834 43764 38836
rect 43708 38782 43710 38834
rect 43710 38782 43762 38834
rect 43762 38782 43764 38834
rect 43708 38780 43764 38782
rect 43708 38274 43764 38276
rect 43708 38222 43710 38274
rect 43710 38222 43762 38274
rect 43762 38222 43764 38274
rect 43708 38220 43764 38222
rect 43596 36876 43652 36932
rect 43820 35868 43876 35924
rect 38668 32508 38724 32510
rect 38108 31724 38164 31780
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 36316 29260 36372 29316
rect 31052 28476 31108 28532
rect 30828 28364 30884 28420
rect 31388 28364 31444 28420
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 31612 28476 31668 28532
rect 31164 28082 31220 28084
rect 31164 28030 31166 28082
rect 31166 28030 31218 28082
rect 31218 28030 31220 28082
rect 31164 28028 31220 28030
rect 31612 27132 31668 27188
rect 34524 28588 34580 28644
rect 35420 28642 35476 28644
rect 30940 26124 30996 26180
rect 30604 26066 30660 26068
rect 30604 26014 30606 26066
rect 30606 26014 30658 26066
rect 30658 26014 30660 26066
rect 30604 26012 30660 26014
rect 30716 25618 30772 25620
rect 30716 25566 30718 25618
rect 30718 25566 30770 25618
rect 30770 25566 30772 25618
rect 30716 25564 30772 25566
rect 32060 28028 32116 28084
rect 32508 27244 32564 27300
rect 32172 27186 32228 27188
rect 32172 27134 32174 27186
rect 32174 27134 32226 27186
rect 32226 27134 32228 27186
rect 32172 27132 32228 27134
rect 33180 27020 33236 27076
rect 32060 25564 32116 25620
rect 31948 24780 32004 24836
rect 30156 24050 30212 24052
rect 30156 23998 30158 24050
rect 30158 23998 30210 24050
rect 30210 23998 30212 24050
rect 30156 23996 30212 23998
rect 31052 23996 31108 24052
rect 29932 23212 29988 23268
rect 30808 23154 30864 23156
rect 30808 23102 30810 23154
rect 30810 23102 30862 23154
rect 30862 23102 30864 23154
rect 30808 23100 30864 23102
rect 30808 22540 30864 22596
rect 29932 22370 29988 22372
rect 29932 22318 29934 22370
rect 29934 22318 29986 22370
rect 29986 22318 29988 22370
rect 29932 22316 29988 22318
rect 30604 22316 30660 22372
rect 29596 21980 29652 22036
rect 29764 21756 29820 21812
rect 29372 21420 29428 21476
rect 28812 19404 28868 19460
rect 28700 18844 28756 18900
rect 28252 18508 28308 18564
rect 28252 18338 28308 18340
rect 28252 18286 28254 18338
rect 28254 18286 28306 18338
rect 28306 18286 28308 18338
rect 28252 18284 28308 18286
rect 28140 18172 28196 18228
rect 28028 16940 28084 16996
rect 28812 18450 28868 18452
rect 28812 18398 28814 18450
rect 28814 18398 28866 18450
rect 28866 18398 28868 18450
rect 28812 18396 28868 18398
rect 28700 18284 28756 18340
rect 28476 17052 28532 17108
rect 28588 17164 28644 17220
rect 27692 16716 27748 16772
rect 27468 16604 27524 16660
rect 27580 16492 27636 16548
rect 27468 16156 27524 16212
rect 27804 16492 27860 16548
rect 27804 16044 27860 16100
rect 26124 15820 26180 15876
rect 27468 15372 27524 15428
rect 26124 15314 26180 15316
rect 26124 15262 26126 15314
rect 26126 15262 26178 15314
rect 26178 15262 26180 15314
rect 26124 15260 26180 15262
rect 26012 15148 26068 15204
rect 26460 14476 26516 14532
rect 26516 14306 26572 14308
rect 26516 14254 26518 14306
rect 26518 14254 26570 14306
rect 26570 14254 26572 14306
rect 26516 14252 26572 14254
rect 27244 14530 27300 14532
rect 27244 14478 27246 14530
rect 27246 14478 27298 14530
rect 27298 14478 27300 14530
rect 27244 14476 27300 14478
rect 27580 15202 27636 15204
rect 27580 15150 27582 15202
rect 27582 15150 27634 15202
rect 27634 15150 27636 15202
rect 27580 15148 27636 15150
rect 28364 16098 28420 16100
rect 28364 16046 28366 16098
rect 28366 16046 28418 16098
rect 28418 16046 28420 16098
rect 28364 16044 28420 16046
rect 28028 15874 28084 15876
rect 28028 15822 28030 15874
rect 28030 15822 28082 15874
rect 28082 15822 28084 15874
rect 28028 15820 28084 15822
rect 28700 15260 28756 15316
rect 28140 14924 28196 14980
rect 29260 18620 29316 18676
rect 29148 18060 29204 18116
rect 30044 21980 30100 22036
rect 30380 21586 30436 21588
rect 30380 21534 30382 21586
rect 30382 21534 30434 21586
rect 30434 21534 30436 21586
rect 30380 21532 30436 21534
rect 30716 21308 30772 21364
rect 29708 20802 29764 20804
rect 29708 20750 29710 20802
rect 29710 20750 29762 20802
rect 29762 20750 29764 20802
rect 29708 20748 29764 20750
rect 29596 19964 29652 20020
rect 30380 20748 30436 20804
rect 29932 20130 29988 20132
rect 29932 20078 29934 20130
rect 29934 20078 29986 20130
rect 29986 20078 29988 20130
rect 29932 20076 29988 20078
rect 29820 19740 29876 19796
rect 30156 19852 30212 19908
rect 30156 19180 30212 19236
rect 29484 18284 29540 18340
rect 29372 17164 29428 17220
rect 29596 17666 29652 17668
rect 29596 17614 29598 17666
rect 29598 17614 29650 17666
rect 29650 17614 29652 17666
rect 29596 17612 29652 17614
rect 30492 20076 30548 20132
rect 30716 20018 30772 20020
rect 30716 19966 30718 20018
rect 30718 19966 30770 20018
rect 30770 19966 30772 20018
rect 30716 19964 30772 19966
rect 30716 18508 30772 18564
rect 30380 17666 30436 17668
rect 30380 17614 30382 17666
rect 30382 17614 30434 17666
rect 30434 17614 30436 17666
rect 30380 17612 30436 17614
rect 30828 18620 30884 18676
rect 30548 17612 30604 17668
rect 30156 17052 30212 17108
rect 29820 16940 29876 16996
rect 29708 16716 29764 16772
rect 29148 16098 29204 16100
rect 29148 16046 29150 16098
rect 29150 16046 29202 16098
rect 29202 16046 29204 16098
rect 29148 16044 29204 16046
rect 29036 15484 29092 15540
rect 29932 16268 29988 16324
rect 29596 16210 29652 16212
rect 29596 16158 29598 16210
rect 29598 16158 29650 16210
rect 29650 16158 29652 16210
rect 29596 16156 29652 16158
rect 29484 15932 29540 15988
rect 29820 15372 29876 15428
rect 28924 14588 28980 14644
rect 29484 14588 29540 14644
rect 28140 14252 28196 14308
rect 28588 14476 28644 14532
rect 26908 13692 26964 13748
rect 27692 13746 27748 13748
rect 27692 13694 27694 13746
rect 27694 13694 27746 13746
rect 27746 13694 27748 13746
rect 27692 13692 27748 13694
rect 28476 13132 28532 13188
rect 25564 8540 25620 8596
rect 25228 8428 25284 8484
rect 27356 12796 27412 12852
rect 26572 12290 26628 12292
rect 26572 12238 26574 12290
rect 26574 12238 26626 12290
rect 26626 12238 26628 12290
rect 26572 12236 26628 12238
rect 26142 11954 26198 11956
rect 26142 11902 26144 11954
rect 26144 11902 26196 11954
rect 26196 11902 26198 11954
rect 26142 11900 26198 11902
rect 26012 11676 26068 11732
rect 28252 12684 28308 12740
rect 27244 12012 27300 12068
rect 27020 11676 27076 11732
rect 26740 11564 26796 11620
rect 27244 10498 27300 10500
rect 27244 10446 27246 10498
rect 27246 10446 27298 10498
rect 27298 10446 27300 10498
rect 27244 10444 27300 10446
rect 30492 16882 30548 16884
rect 30492 16830 30494 16882
rect 30494 16830 30546 16882
rect 30546 16830 30548 16882
rect 30492 16828 30548 16830
rect 30828 16882 30884 16884
rect 30828 16830 30830 16882
rect 30830 16830 30882 16882
rect 30882 16830 30884 16882
rect 30828 16828 30884 16830
rect 30604 15932 30660 15988
rect 30492 15372 30548 15428
rect 30604 14924 30660 14980
rect 31388 23436 31444 23492
rect 33068 26290 33124 26292
rect 33068 26238 33070 26290
rect 33070 26238 33122 26290
rect 33122 26238 33124 26290
rect 33068 26236 33124 26238
rect 34076 27132 34132 27188
rect 33628 27074 33684 27076
rect 33628 27022 33630 27074
rect 33630 27022 33682 27074
rect 33682 27022 33684 27074
rect 33628 27020 33684 27022
rect 35420 28590 35422 28642
rect 35422 28590 35474 28642
rect 35474 28590 35476 28642
rect 35420 28588 35476 28590
rect 35980 28476 36036 28532
rect 36260 28418 36316 28420
rect 36260 28366 36262 28418
rect 36262 28366 36314 28418
rect 36314 28366 36316 28418
rect 36260 28364 36316 28366
rect 36428 28252 36484 28308
rect 35756 28028 35812 28084
rect 33628 26290 33684 26292
rect 33628 26238 33630 26290
rect 33630 26238 33682 26290
rect 33682 26238 33684 26290
rect 33628 26236 33684 26238
rect 32508 25340 32564 25396
rect 32396 24108 32452 24164
rect 31500 23100 31556 23156
rect 31500 22876 31556 22932
rect 31612 21756 31668 21812
rect 31332 20578 31388 20580
rect 31332 20526 31334 20578
rect 31334 20526 31386 20578
rect 31386 20526 31388 20578
rect 31332 20524 31388 20526
rect 31388 19852 31444 19908
rect 31388 18508 31444 18564
rect 32172 23212 32228 23268
rect 32060 23154 32116 23156
rect 32060 23102 32062 23154
rect 32062 23102 32114 23154
rect 32114 23102 32116 23154
rect 32060 23100 32116 23102
rect 39564 31778 39620 31780
rect 39564 31726 39566 31778
rect 39566 31726 39618 31778
rect 39618 31726 39620 31778
rect 39564 31724 39620 31726
rect 42252 31890 42308 31892
rect 42252 31838 42254 31890
rect 42254 31838 42306 31890
rect 42306 31838 42308 31890
rect 42252 31836 42308 31838
rect 40012 30716 40068 30772
rect 40460 30322 40516 30324
rect 40460 30270 40462 30322
rect 40462 30270 40514 30322
rect 40514 30270 40516 30322
rect 40460 30268 40516 30270
rect 36876 29426 36932 29428
rect 36876 29374 36878 29426
rect 36878 29374 36930 29426
rect 36930 29374 36932 29426
rect 36876 29372 36932 29374
rect 37212 29260 37268 29316
rect 37324 29372 37380 29428
rect 36708 28588 36764 28644
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35868 27468 35924 27524
rect 35084 26796 35140 26852
rect 36652 28364 36708 28420
rect 34748 26066 34804 26068
rect 34748 26014 34750 26066
rect 34750 26014 34802 26066
rect 34802 26014 34804 26066
rect 34748 26012 34804 26014
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34636 25676 34692 25732
rect 34972 25394 35028 25396
rect 34972 25342 34974 25394
rect 34974 25342 35026 25394
rect 35026 25342 35028 25394
rect 34972 25340 35028 25342
rect 33292 23996 33348 24052
rect 33628 24050 33684 24052
rect 33628 23998 33630 24050
rect 33630 23998 33682 24050
rect 33682 23998 33684 24050
rect 33628 23996 33684 23998
rect 32732 23324 32788 23380
rect 33572 23378 33628 23380
rect 33572 23326 33574 23378
rect 33574 23326 33626 23378
rect 33626 23326 33628 23378
rect 33572 23324 33628 23326
rect 32508 23100 32564 23156
rect 33292 23154 33348 23156
rect 33292 23102 33294 23154
rect 33294 23102 33346 23154
rect 33346 23102 33348 23154
rect 33292 23100 33348 23102
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35532 23938 35588 23940
rect 35532 23886 35534 23938
rect 35534 23886 35586 23938
rect 35586 23886 35588 23938
rect 35532 23884 35588 23886
rect 36316 27186 36372 27188
rect 36316 27134 36318 27186
rect 36318 27134 36370 27186
rect 36370 27134 36372 27186
rect 36316 27132 36372 27134
rect 36652 27020 36708 27076
rect 36876 28252 36932 28308
rect 36988 27468 37044 27524
rect 36876 27132 36932 27188
rect 36092 26908 36148 26964
rect 36988 26908 37044 26964
rect 37212 28476 37268 28532
rect 37436 28476 37492 28532
rect 37548 27804 37604 27860
rect 37772 29260 37828 29316
rect 37884 28642 37940 28644
rect 37884 28590 37886 28642
rect 37886 28590 37938 28642
rect 37938 28590 37940 28642
rect 37884 28588 37940 28590
rect 37996 27298 38052 27300
rect 37996 27246 37998 27298
rect 37998 27246 38050 27298
rect 38050 27246 38052 27298
rect 37996 27244 38052 27246
rect 37324 26348 37380 26404
rect 38668 28754 38724 28756
rect 38668 28702 38670 28754
rect 38670 28702 38722 28754
rect 38722 28702 38724 28754
rect 38668 28700 38724 28702
rect 38556 28476 38612 28532
rect 39340 29314 39396 29316
rect 39340 29262 39342 29314
rect 39342 29262 39394 29314
rect 39394 29262 39396 29314
rect 39340 29260 39396 29262
rect 38892 28028 38948 28084
rect 39676 27858 39732 27860
rect 39676 27806 39678 27858
rect 39678 27806 39730 27858
rect 39730 27806 39732 27858
rect 39676 27804 39732 27806
rect 38556 27020 38612 27076
rect 39676 27074 39732 27076
rect 39676 27022 39678 27074
rect 39678 27022 39730 27074
rect 39730 27022 39732 27074
rect 39676 27020 39732 27022
rect 37100 25564 37156 25620
rect 36540 25506 36596 25508
rect 36540 25454 36542 25506
rect 36542 25454 36594 25506
rect 36594 25454 36596 25506
rect 36540 25452 36596 25454
rect 36316 25228 36372 25284
rect 31836 22316 31892 22372
rect 33852 22316 33908 22372
rect 32060 21644 32116 21700
rect 32340 21980 32396 22036
rect 33292 22092 33348 22148
rect 32172 21532 32228 21588
rect 32956 21756 33012 21812
rect 32060 21084 32116 21140
rect 31724 20748 31780 20804
rect 32508 20802 32564 20804
rect 32508 20750 32510 20802
rect 32510 20750 32562 20802
rect 32562 20750 32564 20802
rect 32508 20748 32564 20750
rect 33852 22146 33908 22148
rect 33852 22094 33854 22146
rect 33854 22094 33906 22146
rect 33906 22094 33908 22146
rect 33852 22092 33908 22094
rect 33740 21084 33796 21140
rect 34860 23154 34916 23156
rect 34860 23102 34862 23154
rect 34862 23102 34914 23154
rect 34914 23102 34916 23154
rect 34860 23100 34916 23102
rect 35532 23100 35588 23156
rect 36092 24108 36148 24164
rect 35980 24050 36036 24052
rect 35980 23998 35982 24050
rect 35982 23998 36034 24050
rect 36034 23998 36036 24050
rect 35980 23996 36036 23998
rect 36988 25340 37044 25396
rect 37100 25228 37156 25284
rect 37436 25676 37492 25732
rect 37436 25228 37492 25284
rect 36316 23938 36372 23940
rect 36316 23886 36318 23938
rect 36318 23886 36370 23938
rect 36370 23886 36372 23938
rect 36316 23884 36372 23886
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35084 22370 35140 22372
rect 35084 22318 35086 22370
rect 35086 22318 35138 22370
rect 35138 22318 35140 22370
rect 35084 22316 35140 22318
rect 34860 21532 34916 21588
rect 32956 20748 33012 20804
rect 33516 20748 33572 20804
rect 32172 19740 32228 19796
rect 33404 18956 33460 19012
rect 31724 18508 31780 18564
rect 32060 18620 32116 18676
rect 33908 20524 33964 20580
rect 34748 20300 34804 20356
rect 34076 20018 34132 20020
rect 34076 19966 34078 20018
rect 34078 19966 34130 20018
rect 34130 19966 34132 20018
rect 34076 19964 34132 19966
rect 33740 18956 33796 19012
rect 32396 18226 32452 18228
rect 32396 18174 32398 18226
rect 32398 18174 32450 18226
rect 32450 18174 32452 18226
rect 32396 18172 32452 18174
rect 31724 17948 31780 18004
rect 31836 17724 31892 17780
rect 31724 17500 31780 17556
rect 31164 17052 31220 17108
rect 31052 16268 31108 16324
rect 31052 15314 31108 15316
rect 31052 15262 31054 15314
rect 31054 15262 31106 15314
rect 31106 15262 31108 15314
rect 31052 15260 31108 15262
rect 30828 15036 30884 15092
rect 30604 14418 30660 14420
rect 30604 14366 30606 14418
rect 30606 14366 30658 14418
rect 30658 14366 30660 14418
rect 30604 14364 30660 14366
rect 29372 13186 29428 13188
rect 29372 13134 29374 13186
rect 29374 13134 29426 13186
rect 29426 13134 29428 13186
rect 29372 13132 29428 13134
rect 30604 13468 30660 13524
rect 29708 12684 29764 12740
rect 28868 12402 28924 12404
rect 28868 12350 28870 12402
rect 28870 12350 28922 12402
rect 28922 12350 28924 12402
rect 28868 12348 28924 12350
rect 28476 10498 28532 10500
rect 28476 10446 28478 10498
rect 28478 10446 28530 10498
rect 28530 10446 28532 10498
rect 28476 10444 28532 10446
rect 26012 10220 26068 10276
rect 27112 10220 27168 10276
rect 25676 8316 25732 8372
rect 25770 8146 25826 8148
rect 25770 8094 25772 8146
rect 25772 8094 25824 8146
rect 25824 8094 25826 8146
rect 25770 8092 25826 8094
rect 26236 9548 26292 9604
rect 26684 8316 26740 8372
rect 26012 8092 26068 8148
rect 25900 7868 25956 7924
rect 26684 7980 26740 8036
rect 27188 8092 27244 8148
rect 27020 7868 27076 7924
rect 26236 7532 26292 7588
rect 25900 6972 25956 7028
rect 25340 5964 25396 6020
rect 25004 5852 25060 5908
rect 25788 6578 25844 6580
rect 25788 6526 25790 6578
rect 25790 6526 25842 6578
rect 25842 6526 25844 6578
rect 25788 6524 25844 6526
rect 26031 6412 26087 6468
rect 27188 7868 27244 7924
rect 26908 6972 26964 7028
rect 27636 8034 27692 8036
rect 27636 7982 27638 8034
rect 27638 7982 27690 8034
rect 27690 7982 27692 8034
rect 27636 7980 27692 7982
rect 29148 8876 29204 8932
rect 29260 8258 29316 8260
rect 29260 8206 29262 8258
rect 29262 8206 29314 8258
rect 29314 8206 29316 8258
rect 29260 8204 29316 8206
rect 28812 8092 28868 8148
rect 28644 7980 28700 8036
rect 30604 13186 30660 13188
rect 30604 13134 30606 13186
rect 30606 13134 30658 13186
rect 30658 13134 30660 13186
rect 30604 13132 30660 13134
rect 31388 16828 31444 16884
rect 31612 16882 31668 16884
rect 31612 16830 31614 16882
rect 31614 16830 31666 16882
rect 31666 16830 31668 16882
rect 31612 16828 31668 16830
rect 31500 16604 31556 16660
rect 31500 15260 31556 15316
rect 31388 15202 31444 15204
rect 31388 15150 31390 15202
rect 31390 15150 31442 15202
rect 31442 15150 31444 15202
rect 31388 15148 31444 15150
rect 32172 17500 32228 17556
rect 32284 17388 32340 17444
rect 32060 16828 32116 16884
rect 31948 16770 32004 16772
rect 31948 16718 31950 16770
rect 31950 16718 32002 16770
rect 32002 16718 32004 16770
rect 31948 16716 32004 16718
rect 31836 16604 31892 16660
rect 31948 16492 32004 16548
rect 32004 15426 32060 15428
rect 32004 15374 32006 15426
rect 32006 15374 32058 15426
rect 32058 15374 32060 15426
rect 32004 15372 32060 15374
rect 31332 14642 31388 14644
rect 31332 14590 31334 14642
rect 31334 14590 31386 14642
rect 31386 14590 31388 14642
rect 31332 14588 31388 14590
rect 31164 14364 31220 14420
rect 31052 13356 31108 13412
rect 30940 13244 30996 13300
rect 31500 13020 31556 13076
rect 31164 12738 31220 12740
rect 31164 12686 31166 12738
rect 31166 12686 31218 12738
rect 31218 12686 31220 12738
rect 31164 12684 31220 12686
rect 29820 11004 29876 11060
rect 30268 10108 30324 10164
rect 30604 9660 30660 9716
rect 30940 8988 30996 9044
rect 29708 8876 29764 8932
rect 29820 8316 29876 8372
rect 27244 6972 27300 7028
rect 25452 5852 25508 5908
rect 26216 5906 26272 5908
rect 26216 5854 26218 5906
rect 26218 5854 26270 5906
rect 26270 5854 26272 5906
rect 26216 5852 26272 5854
rect 28364 6972 28420 7028
rect 28252 6748 28308 6804
rect 28120 6690 28176 6692
rect 28120 6638 28122 6690
rect 28122 6638 28174 6690
rect 28174 6638 28176 6690
rect 28120 6636 28176 6638
rect 27244 6300 27300 6356
rect 25788 5068 25844 5124
rect 26796 5068 26852 5124
rect 24332 4396 24388 4452
rect 29932 8204 29988 8260
rect 29484 7532 29540 7588
rect 30156 7868 30212 7924
rect 29372 7474 29428 7476
rect 29372 7422 29374 7474
rect 29374 7422 29426 7474
rect 29426 7422 29428 7474
rect 29372 7420 29428 7422
rect 28644 6748 28700 6804
rect 29372 6636 29428 6692
rect 27692 6076 27748 6132
rect 30044 7586 30100 7588
rect 30044 7534 30046 7586
rect 30046 7534 30098 7586
rect 30098 7534 30100 7586
rect 30044 7532 30100 7534
rect 28568 5906 28624 5908
rect 28568 5854 28570 5906
rect 28570 5854 28622 5906
rect 28622 5854 28624 5906
rect 28568 5852 28624 5854
rect 27468 5180 27524 5236
rect 28028 5122 28084 5124
rect 28028 5070 28030 5122
rect 28030 5070 28082 5122
rect 28082 5070 28084 5122
rect 28028 5068 28084 5070
rect 27244 4508 27300 4564
rect 25564 3778 25620 3780
rect 25564 3726 25566 3778
rect 25566 3726 25618 3778
rect 25618 3726 25620 3778
rect 25564 3724 25620 3726
rect 28700 4450 28756 4452
rect 28700 4398 28702 4450
rect 28702 4398 28754 4450
rect 28754 4398 28756 4450
rect 28700 4396 28756 4398
rect 29652 6690 29708 6692
rect 29652 6638 29654 6690
rect 29654 6638 29706 6690
rect 29706 6638 29708 6690
rect 29652 6636 29708 6638
rect 31724 13522 31780 13524
rect 31724 13470 31726 13522
rect 31726 13470 31778 13522
rect 31778 13470 31780 13522
rect 31724 13468 31780 13470
rect 31724 13244 31780 13300
rect 31724 11564 31780 11620
rect 31836 12124 31892 12180
rect 31724 11340 31780 11396
rect 32844 17666 32900 17668
rect 32844 17614 32846 17666
rect 32846 17614 32898 17666
rect 32898 17614 32900 17666
rect 32844 17612 32900 17614
rect 33180 17442 33236 17444
rect 33180 17390 33182 17442
rect 33182 17390 33234 17442
rect 33234 17390 33236 17442
rect 33180 17388 33236 17390
rect 32508 16268 32564 16324
rect 34020 19010 34076 19012
rect 34020 18958 34022 19010
rect 34022 18958 34074 19010
rect 34074 18958 34076 19010
rect 34020 18956 34076 18958
rect 35644 21756 35700 21812
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 20914 35252 20916
rect 35196 20862 35198 20914
rect 35198 20862 35250 20914
rect 35250 20862 35252 20914
rect 35196 20860 35252 20862
rect 35084 19964 35140 20020
rect 35980 22930 36036 22932
rect 35980 22878 35982 22930
rect 35982 22878 36034 22930
rect 36034 22878 36036 22930
rect 35980 22876 36036 22878
rect 35960 21756 36016 21812
rect 35756 20860 35812 20916
rect 35644 20524 35700 20580
rect 35812 20300 35868 20356
rect 35868 19964 35924 20020
rect 35532 19852 35588 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35980 19292 36036 19348
rect 34300 17836 34356 17892
rect 33852 17724 33908 17780
rect 32396 15372 32452 15428
rect 32284 12962 32340 12964
rect 32284 12910 32286 12962
rect 32286 12910 32338 12962
rect 32338 12910 32340 12962
rect 32284 12908 32340 12910
rect 32956 15314 33012 15316
rect 32956 15262 32958 15314
rect 32958 15262 33010 15314
rect 33010 15262 33012 15314
rect 32956 15260 33012 15262
rect 32956 13468 33012 13524
rect 34076 17500 34132 17556
rect 35868 18508 35924 18564
rect 35756 18284 35812 18340
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35588 18060 35644 18116
rect 34804 17836 34860 17892
rect 34972 17724 35028 17780
rect 35420 17666 35476 17668
rect 35420 17614 35422 17666
rect 35422 17614 35474 17666
rect 35474 17614 35476 17666
rect 35420 17612 35476 17614
rect 37772 26402 37828 26404
rect 37772 26350 37774 26402
rect 37774 26350 37826 26402
rect 37826 26350 37828 26402
rect 37772 26348 37828 26350
rect 37548 24668 37604 24724
rect 37660 26124 37716 26180
rect 37996 25452 38052 25508
rect 38556 26348 38612 26404
rect 41020 28028 41076 28084
rect 39788 25228 39844 25284
rect 39900 25340 39956 25396
rect 39676 25004 39732 25060
rect 38220 23996 38276 24052
rect 37548 23436 37604 23492
rect 38108 23436 38164 23492
rect 37100 22988 37156 23044
rect 36204 22594 36260 22596
rect 36204 22542 36206 22594
rect 36206 22542 36258 22594
rect 36258 22542 36260 22594
rect 36204 22540 36260 22542
rect 36988 22370 37044 22372
rect 36988 22318 36990 22370
rect 36990 22318 37042 22370
rect 37042 22318 37044 22370
rect 36988 22316 37044 22318
rect 38108 22652 38164 22708
rect 38332 22540 38388 22596
rect 38220 22428 38276 22484
rect 37772 21756 37828 21812
rect 39116 24722 39172 24724
rect 39116 24670 39118 24722
rect 39118 24670 39170 24722
rect 39170 24670 39172 24722
rect 39116 24668 39172 24670
rect 39992 24722 40048 24724
rect 39992 24670 39994 24722
rect 39994 24670 40046 24722
rect 40046 24670 40048 24722
rect 39992 24668 40048 24670
rect 38556 22876 38612 22932
rect 38668 22652 38724 22708
rect 38668 22482 38724 22484
rect 38668 22430 38670 22482
rect 38670 22430 38722 22482
rect 38722 22430 38724 22482
rect 38668 22428 38724 22430
rect 38892 22652 38948 22708
rect 39004 22540 39060 22596
rect 38556 21756 38612 21812
rect 39676 23884 39732 23940
rect 39116 21756 39172 21812
rect 39564 21532 39620 21588
rect 38444 20076 38500 20132
rect 37156 19292 37212 19348
rect 36988 19180 37044 19236
rect 36988 18508 37044 18564
rect 38780 20636 38836 20692
rect 38668 20018 38724 20020
rect 38668 19966 38670 20018
rect 38670 19966 38722 20018
rect 38722 19966 38724 20018
rect 38668 19964 38724 19966
rect 37772 19292 37828 19348
rect 38668 19292 38724 19348
rect 38780 19180 38836 19236
rect 37660 18620 37716 18676
rect 36204 18450 36260 18452
rect 36204 18398 36206 18450
rect 36206 18398 36258 18450
rect 36258 18398 36260 18450
rect 36204 18396 36260 18398
rect 35868 17612 35924 17668
rect 36092 17666 36148 17668
rect 36092 17614 36094 17666
rect 36094 17614 36146 17666
rect 36146 17614 36148 17666
rect 36092 17612 36148 17614
rect 34300 17052 34356 17108
rect 34188 16828 34244 16884
rect 34524 15986 34580 15988
rect 34524 15934 34526 15986
rect 34526 15934 34578 15986
rect 34578 15934 34580 15986
rect 34524 15932 34580 15934
rect 33292 13468 33348 13524
rect 33628 13356 33684 13412
rect 33460 12908 33516 12964
rect 33068 12684 33124 12740
rect 31612 10108 31668 10164
rect 31948 9042 32004 9044
rect 31948 8990 31950 9042
rect 31950 8990 32002 9042
rect 32002 8990 32004 9042
rect 31948 8988 32004 8990
rect 31164 8370 31220 8372
rect 31164 8318 31166 8370
rect 31166 8318 31218 8370
rect 31218 8318 31220 8370
rect 31164 8316 31220 8318
rect 34804 17106 34860 17108
rect 34804 17054 34806 17106
rect 34806 17054 34858 17106
rect 34858 17054 34860 17106
rect 34804 17052 34860 17054
rect 34972 16828 35028 16884
rect 35980 17106 36036 17108
rect 35980 17054 35982 17106
rect 35982 17054 36034 17106
rect 36034 17054 36036 17106
rect 35980 17052 36036 17054
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35644 16882 35700 16884
rect 35644 16830 35646 16882
rect 35646 16830 35698 16882
rect 35698 16830 35700 16882
rect 35644 16828 35700 16830
rect 35308 15874 35364 15876
rect 35308 15822 35310 15874
rect 35310 15822 35362 15874
rect 35362 15822 35364 15874
rect 35308 15820 35364 15822
rect 35532 15090 35588 15092
rect 35532 15038 35534 15090
rect 35534 15038 35586 15090
rect 35586 15038 35588 15090
rect 35532 15036 35588 15038
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 14530 35252 14532
rect 35196 14478 35198 14530
rect 35198 14478 35250 14530
rect 35250 14478 35252 14530
rect 35196 14476 35252 14478
rect 35980 14476 36036 14532
rect 35700 14252 35756 14308
rect 35868 14418 35924 14420
rect 35868 14366 35870 14418
rect 35870 14366 35922 14418
rect 35922 14366 35924 14418
rect 35868 14364 35924 14366
rect 33740 12796 33796 12852
rect 32284 11228 32340 11284
rect 32508 11394 32564 11396
rect 32508 11342 32510 11394
rect 32510 11342 32562 11394
rect 32562 11342 32564 11394
rect 32508 11340 32564 11342
rect 33068 11340 33124 11396
rect 32396 11116 32452 11172
rect 32508 11004 32564 11060
rect 32620 10668 32676 10724
rect 32620 10332 32676 10388
rect 32172 9324 32228 9380
rect 32956 8876 33012 8932
rect 31948 8092 32004 8148
rect 31052 7532 31108 7588
rect 30156 6412 30212 6468
rect 29596 5852 29652 5908
rect 31668 6466 31724 6468
rect 31668 6414 31670 6466
rect 31670 6414 31722 6466
rect 31722 6414 31724 6466
rect 31668 6412 31724 6414
rect 32284 8204 32340 8260
rect 32172 6076 32228 6132
rect 28364 3724 28420 3780
rect 29036 4284 29092 4340
rect 30268 4338 30324 4340
rect 24108 3500 24164 3556
rect 24556 3526 24612 3556
rect 24556 3500 24558 3526
rect 24558 3500 24610 3526
rect 24610 3500 24612 3526
rect 30268 4286 30270 4338
rect 30270 4286 30322 4338
rect 30322 4286 30324 4338
rect 30268 4284 30324 4286
rect 29278 3778 29334 3780
rect 29278 3726 29280 3778
rect 29280 3726 29332 3778
rect 29332 3726 29334 3778
rect 29278 3724 29334 3726
rect 33852 12348 33908 12404
rect 34076 13468 34132 13524
rect 34356 12962 34412 12964
rect 34356 12910 34358 12962
rect 34358 12910 34410 12962
rect 34410 12910 34412 12962
rect 34356 12908 34412 12910
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35868 13468 35924 13524
rect 35980 14252 36036 14308
rect 35980 13580 36036 13636
rect 36092 13916 36148 13972
rect 35420 12908 35476 12964
rect 34972 12684 35028 12740
rect 35102 12460 35158 12516
rect 35756 12962 35812 12964
rect 35756 12910 35758 12962
rect 35758 12910 35810 12962
rect 35810 12910 35812 12962
rect 35756 12908 35812 12910
rect 36092 13020 36148 13076
rect 35420 12236 35476 12292
rect 35980 12908 36036 12964
rect 37548 18396 37604 18452
rect 36764 18060 36820 18116
rect 36316 17836 36372 17892
rect 37212 17890 37268 17892
rect 37212 17838 37214 17890
rect 37214 17838 37266 17890
rect 37266 17838 37268 17890
rect 37212 17836 37268 17838
rect 38668 17836 38724 17892
rect 40012 21980 40068 22036
rect 39564 19852 39620 19908
rect 40236 24892 40292 24948
rect 40348 25676 40404 25732
rect 40236 23884 40292 23940
rect 40460 25452 40516 25508
rect 40796 25618 40852 25620
rect 40796 25566 40798 25618
rect 40798 25566 40850 25618
rect 40850 25566 40852 25618
rect 40796 25564 40852 25566
rect 40684 25340 40740 25396
rect 40908 25340 40964 25396
rect 40684 25004 40740 25060
rect 41244 29260 41300 29316
rect 41916 30716 41972 30772
rect 43148 32956 43204 33012
rect 43484 35586 43540 35588
rect 43484 35534 43486 35586
rect 43486 35534 43538 35586
rect 43538 35534 43540 35586
rect 43484 35532 43540 35534
rect 43260 31836 43316 31892
rect 42700 30770 42756 30772
rect 42700 30718 42702 30770
rect 42702 30718 42754 30770
rect 42754 30718 42756 30770
rect 42700 30716 42756 30718
rect 42924 30268 42980 30324
rect 41692 28812 41748 28868
rect 41356 28700 41412 28756
rect 41244 28588 41300 28644
rect 41244 27244 41300 27300
rect 41020 24050 41076 24052
rect 41020 23998 41022 24050
rect 41022 23998 41074 24050
rect 41074 23998 41076 24050
rect 41020 23996 41076 23998
rect 40460 23212 40516 23268
rect 41692 27244 41748 27300
rect 41356 23117 41358 23156
rect 41358 23117 41410 23156
rect 41410 23117 41412 23156
rect 41356 23100 41412 23117
rect 42140 27020 42196 27076
rect 43372 29650 43428 29652
rect 43372 29598 43374 29650
rect 43374 29598 43426 29650
rect 43426 29598 43428 29650
rect 43372 29596 43428 29598
rect 43596 28812 43652 28868
rect 43484 28588 43540 28644
rect 43708 26908 43764 26964
rect 41692 24892 41748 24948
rect 42700 25394 42756 25396
rect 42700 25342 42702 25394
rect 42702 25342 42754 25394
rect 42754 25342 42756 25394
rect 42700 25340 42756 25342
rect 42364 24946 42420 24948
rect 42364 24894 42366 24946
rect 42366 24894 42418 24946
rect 42418 24894 42420 24946
rect 42364 24892 42420 24894
rect 43820 26572 43876 26628
rect 44044 26348 44100 26404
rect 44268 26236 44324 26292
rect 43820 25506 43876 25508
rect 43820 25454 43822 25506
rect 43822 25454 43874 25506
rect 43874 25454 43876 25506
rect 43820 25452 43876 25454
rect 41916 23436 41972 23492
rect 43036 23212 43092 23268
rect 40572 22652 40628 22708
rect 40124 21308 40180 21364
rect 40124 20802 40180 20804
rect 40124 20750 40126 20802
rect 40126 20750 40178 20802
rect 40178 20750 40180 20802
rect 40124 20748 40180 20750
rect 40124 20412 40180 20468
rect 43036 22764 43092 22820
rect 42252 22652 42308 22708
rect 42924 22594 42980 22596
rect 42924 22542 42926 22594
rect 42926 22542 42978 22594
rect 42978 22542 42980 22594
rect 42924 22540 42980 22542
rect 42140 21644 42196 21700
rect 41132 21586 41188 21588
rect 41132 21534 41134 21586
rect 41134 21534 41186 21586
rect 41186 21534 41188 21586
rect 41132 21532 41188 21534
rect 41300 20802 41356 20804
rect 41300 20750 41302 20802
rect 41302 20750 41354 20802
rect 41354 20750 41356 20802
rect 41300 20748 41356 20750
rect 40796 20690 40852 20692
rect 40796 20638 40798 20690
rect 40798 20638 40850 20690
rect 40850 20638 40852 20690
rect 40796 20636 40852 20638
rect 39770 19458 39826 19460
rect 39770 19406 39772 19458
rect 39772 19406 39824 19458
rect 39824 19406 39826 19458
rect 39770 19404 39826 19406
rect 40124 19852 40180 19908
rect 39452 19180 39508 19236
rect 39340 18396 39396 18452
rect 39788 18450 39844 18452
rect 39788 18398 39790 18450
rect 39790 18398 39842 18450
rect 39842 18398 39844 18450
rect 39788 18396 39844 18398
rect 39788 17164 39844 17220
rect 39116 16828 39172 16884
rect 36540 15820 36596 15876
rect 36372 15484 36428 15540
rect 36372 15202 36428 15204
rect 36372 15150 36374 15202
rect 36374 15150 36426 15202
rect 36426 15150 36428 15202
rect 36372 15148 36428 15150
rect 36764 15314 36820 15316
rect 36764 15262 36766 15314
rect 36766 15262 36818 15314
rect 36818 15262 36820 15314
rect 36764 15260 36820 15262
rect 38444 16156 38500 16212
rect 36372 14530 36428 14532
rect 36372 14478 36374 14530
rect 36374 14478 36426 14530
rect 36426 14478 36428 14530
rect 36372 14476 36428 14478
rect 35084 12178 35140 12180
rect 35084 12126 35086 12178
rect 35086 12126 35138 12178
rect 35138 12126 35140 12178
rect 35084 12124 35140 12126
rect 33964 12012 34020 12068
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35644 12236 35700 12292
rect 34300 11452 34356 11508
rect 33944 11116 34000 11172
rect 34188 10610 34244 10612
rect 34188 10558 34190 10610
rect 34190 10558 34242 10610
rect 34242 10558 34244 10610
rect 34188 10556 34244 10558
rect 34076 8764 34132 8820
rect 34860 11340 34916 11396
rect 34412 10668 34468 10724
rect 34636 10668 34692 10724
rect 35084 10332 35140 10388
rect 36148 12738 36204 12740
rect 36148 12686 36150 12738
rect 36150 12686 36202 12738
rect 36202 12686 36204 12738
rect 36148 12684 36204 12686
rect 36092 12460 36148 12516
rect 36428 12402 36484 12404
rect 36428 12350 36430 12402
rect 36430 12350 36482 12402
rect 36482 12350 36484 12402
rect 36428 12348 36484 12350
rect 35868 11506 35924 11508
rect 35868 11454 35870 11506
rect 35870 11454 35922 11506
rect 35922 11454 35924 11506
rect 35868 11452 35924 11454
rect 35980 11379 36036 11396
rect 35980 11340 35982 11379
rect 35982 11340 36034 11379
rect 36034 11340 36036 11379
rect 36204 11394 36260 11396
rect 36204 11342 36206 11394
rect 36206 11342 36258 11394
rect 36258 11342 36260 11394
rect 36204 11340 36260 11342
rect 35644 10444 35700 10500
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 9826 35252 9828
rect 35196 9774 35198 9826
rect 35198 9774 35250 9826
rect 35250 9774 35252 9826
rect 35196 9772 35252 9774
rect 35532 9436 35588 9492
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35868 9212 35924 9268
rect 36876 15036 36932 15092
rect 37212 15314 37268 15316
rect 37212 15262 37214 15314
rect 37214 15262 37266 15314
rect 37266 15262 37268 15314
rect 37212 15260 37268 15262
rect 37100 14700 37156 14756
rect 36988 14418 37044 14420
rect 36988 14366 36990 14418
rect 36990 14366 37042 14418
rect 37042 14366 37044 14418
rect 36988 14364 37044 14366
rect 39340 16156 39396 16212
rect 40236 19740 40292 19796
rect 40796 19404 40852 19460
rect 40516 19292 40572 19348
rect 41132 19794 41188 19796
rect 41132 19742 41134 19794
rect 41134 19742 41186 19794
rect 41186 19742 41188 19794
rect 41132 19740 41188 19742
rect 40908 19234 40964 19236
rect 40908 19182 40910 19234
rect 40910 19182 40962 19234
rect 40962 19182 40964 19234
rect 40908 19180 40964 19182
rect 40684 19122 40740 19124
rect 40684 19070 40686 19122
rect 40686 19070 40738 19122
rect 40738 19070 40740 19122
rect 40684 19068 40740 19070
rect 40796 18450 40852 18452
rect 40796 18398 40798 18450
rect 40798 18398 40850 18450
rect 40850 18398 40852 18450
rect 40796 18396 40852 18398
rect 40684 18060 40740 18116
rect 40012 17612 40068 17668
rect 41076 17164 41132 17220
rect 41860 19964 41916 20020
rect 43372 23436 43428 23492
rect 43484 23146 43486 23156
rect 43486 23146 43538 23156
rect 43538 23146 43540 23156
rect 43484 23100 43540 23146
rect 43932 24498 43988 24500
rect 43932 24446 43934 24498
rect 43934 24446 43986 24498
rect 43986 24446 43988 24498
rect 43932 24444 43988 24446
rect 44156 25900 44212 25956
rect 44380 26572 44436 26628
rect 44380 25452 44436 25508
rect 44380 24668 44436 24724
rect 43820 23212 43876 23268
rect 43596 22764 43652 22820
rect 43148 20802 43204 20804
rect 43148 20750 43150 20802
rect 43150 20750 43202 20802
rect 43202 20750 43204 20802
rect 43148 20748 43204 20750
rect 41804 19292 41860 19348
rect 42700 18620 42756 18676
rect 42812 18284 42868 18340
rect 42812 17724 42868 17780
rect 41692 17052 41748 17108
rect 41692 16882 41748 16884
rect 41692 16830 41694 16882
rect 41694 16830 41746 16882
rect 41746 16830 41748 16882
rect 42364 16994 42420 16996
rect 42364 16942 42366 16994
rect 42366 16942 42418 16994
rect 42418 16942 42420 16994
rect 42364 16940 42420 16942
rect 44492 24444 44548 24500
rect 43148 19292 43204 19348
rect 43484 21644 43540 21700
rect 43036 18396 43092 18452
rect 43148 19068 43204 19124
rect 41692 16828 41748 16830
rect 43372 19794 43428 19796
rect 43372 19742 43374 19794
rect 43374 19742 43426 19794
rect 43426 19742 43428 19794
rect 43372 19740 43428 19742
rect 44268 20748 44324 20804
rect 43596 19628 43652 19684
rect 43708 20018 43764 20020
rect 43708 19966 43710 20018
rect 43710 19966 43762 20018
rect 43762 19966 43764 20018
rect 43708 19964 43764 19966
rect 43708 19516 43764 19572
rect 44044 19906 44100 19908
rect 44044 19854 44046 19906
rect 44046 19854 44098 19906
rect 44098 19854 44100 19906
rect 44044 19852 44100 19854
rect 43260 18620 43316 18676
rect 43484 18620 43540 18676
rect 43596 18396 43652 18452
rect 42924 17106 42980 17108
rect 42924 17054 42926 17106
rect 42926 17054 42978 17106
rect 42978 17054 42980 17106
rect 42924 17052 42980 17054
rect 43820 18284 43876 18340
rect 43932 17778 43988 17780
rect 43932 17726 43934 17778
rect 43934 17726 43986 17778
rect 43986 17726 43988 17778
rect 43932 17724 43988 17726
rect 43820 17164 43876 17220
rect 43148 16940 43204 16996
rect 42812 16828 42868 16884
rect 43540 16268 43596 16324
rect 39900 16156 39956 16212
rect 40292 16210 40348 16212
rect 40292 16158 40294 16210
rect 40294 16158 40346 16210
rect 40346 16158 40348 16210
rect 40292 16156 40348 16158
rect 37324 13916 37380 13972
rect 37660 15148 37716 15204
rect 37772 14700 37828 14756
rect 37996 14700 38052 14756
rect 39116 15986 39172 15988
rect 39116 15934 39118 15986
rect 39118 15934 39170 15986
rect 39170 15934 39172 15986
rect 39116 15932 39172 15934
rect 41468 15932 41524 15988
rect 40796 15260 40852 15316
rect 38780 14754 38836 14756
rect 38780 14702 38782 14754
rect 38782 14702 38834 14754
rect 38834 14702 38836 14754
rect 38780 14700 38836 14702
rect 37902 14418 37958 14420
rect 37902 14366 37904 14418
rect 37904 14366 37956 14418
rect 37956 14366 37958 14418
rect 37902 14364 37958 14366
rect 39116 14364 39172 14420
rect 37660 13916 37716 13972
rect 38780 13634 38836 13636
rect 38780 13582 38782 13634
rect 38782 13582 38834 13634
rect 38834 13582 38836 13634
rect 38780 13580 38836 13582
rect 37100 12850 37156 12852
rect 37100 12798 37102 12850
rect 37102 12798 37154 12850
rect 37154 12798 37156 12850
rect 37100 12796 37156 12798
rect 37324 12153 37326 12180
rect 37326 12153 37378 12180
rect 37378 12153 37380 12180
rect 37324 12124 37380 12153
rect 39788 12962 39844 12964
rect 39788 12910 39790 12962
rect 39790 12910 39842 12962
rect 39842 12910 39844 12962
rect 39788 12908 39844 12910
rect 37772 12124 37828 12180
rect 38892 12796 38948 12852
rect 37212 11228 37268 11284
rect 36652 10780 36708 10836
rect 36316 10050 36372 10052
rect 36316 9998 36318 10050
rect 36318 9998 36370 10050
rect 36370 9998 36372 10050
rect 36316 9996 36372 9998
rect 36540 9996 36596 10052
rect 34412 8092 34468 8148
rect 34188 7420 34244 7476
rect 33740 6076 33796 6132
rect 33908 5906 33964 5908
rect 33908 5854 33910 5906
rect 33910 5854 33962 5906
rect 33962 5854 33964 5906
rect 33908 5852 33964 5854
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34748 6300 34804 6356
rect 35252 6188 35308 6244
rect 35420 6636 35476 6692
rect 34654 5682 34710 5684
rect 34654 5630 34656 5682
rect 34656 5630 34708 5682
rect 34708 5630 34710 5682
rect 34654 5628 34710 5630
rect 33740 5122 33796 5124
rect 33740 5070 33742 5122
rect 33742 5070 33794 5122
rect 33794 5070 33796 5122
rect 33740 5068 33796 5070
rect 33628 4284 33684 4340
rect 35756 7474 35812 7476
rect 35756 7422 35758 7474
rect 35758 7422 35810 7474
rect 35810 7422 35812 7474
rect 35756 7420 35812 7422
rect 36204 8930 36260 8932
rect 36204 8878 36206 8930
rect 36206 8878 36258 8930
rect 36258 8878 36260 8930
rect 36204 8876 36260 8878
rect 36652 8764 36708 8820
rect 36092 7980 36148 8036
rect 36540 8316 36596 8372
rect 35644 6524 35700 6580
rect 35756 6412 35812 6468
rect 35532 5964 35588 6020
rect 35663 5906 35719 5908
rect 35663 5854 35665 5906
rect 35665 5854 35717 5906
rect 35717 5854 35719 5906
rect 35663 5852 35719 5854
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 36540 6076 36596 6132
rect 35868 5516 35924 5572
rect 36316 5122 36372 5124
rect 36316 5070 36318 5122
rect 36318 5070 36370 5122
rect 36370 5070 36372 5122
rect 36316 5068 36372 5070
rect 36652 5068 36708 5124
rect 34860 4508 34916 4564
rect 36092 4508 36148 4564
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 37324 8988 37380 9044
rect 37212 8316 37268 8372
rect 37212 7980 37268 8036
rect 36988 7756 37044 7812
rect 36876 7532 36932 7588
rect 37100 7644 37156 7700
rect 36988 6690 37044 6692
rect 36988 6638 36990 6690
rect 36990 6638 37042 6690
rect 37042 6638 37044 6690
rect 36988 6636 37044 6638
rect 37324 7644 37380 7700
rect 37324 6748 37380 6804
rect 37548 8230 37604 8260
rect 37548 8204 37550 8230
rect 37550 8204 37602 8230
rect 37602 8204 37604 8230
rect 38780 10610 38836 10612
rect 38780 10558 38782 10610
rect 38782 10558 38834 10610
rect 38834 10558 38836 10610
rect 38780 10556 38836 10558
rect 37996 9266 38052 9268
rect 37996 9214 37998 9266
rect 37998 9214 38050 9266
rect 38050 9214 38052 9266
rect 37996 9212 38052 9214
rect 37884 8316 37940 8372
rect 40460 13746 40516 13748
rect 40460 13694 40462 13746
rect 40462 13694 40514 13746
rect 40514 13694 40516 13746
rect 40460 13692 40516 13694
rect 40124 13020 40180 13076
rect 41188 13970 41244 13972
rect 41188 13918 41190 13970
rect 41190 13918 41242 13970
rect 41242 13918 41244 13970
rect 41188 13916 41244 13918
rect 43652 15538 43708 15540
rect 43652 15486 43654 15538
rect 43654 15486 43706 15538
rect 43706 15486 43708 15538
rect 43652 15484 43708 15486
rect 41580 15036 41636 15092
rect 41468 13858 41524 13860
rect 41468 13806 41470 13858
rect 41470 13806 41522 13858
rect 41522 13806 41524 13858
rect 41468 13804 41524 13806
rect 41636 14140 41692 14196
rect 42382 15090 42438 15092
rect 42382 15038 42384 15090
rect 42384 15038 42436 15090
rect 42436 15038 42438 15090
rect 42382 15036 42438 15038
rect 42140 14812 42196 14868
rect 43036 15202 43092 15204
rect 43036 15150 43038 15202
rect 43038 15150 43090 15202
rect 43090 15150 43092 15202
rect 43036 15148 43092 15150
rect 42140 14252 42196 14308
rect 43372 15036 43428 15092
rect 43148 13916 43204 13972
rect 42906 13746 42962 13748
rect 42906 13694 42908 13746
rect 42908 13694 42960 13746
rect 42960 13694 42962 13746
rect 42906 13692 42962 13694
rect 41804 13468 41860 13524
rect 43260 13356 43316 13412
rect 41356 13074 41412 13076
rect 41356 13022 41358 13074
rect 41358 13022 41410 13074
rect 41410 13022 41412 13074
rect 41356 13020 41412 13022
rect 40572 12962 40628 12964
rect 40572 12910 40574 12962
rect 40574 12910 40626 12962
rect 40626 12910 40628 12962
rect 40572 12908 40628 12910
rect 40908 12178 40964 12180
rect 40908 12126 40910 12178
rect 40910 12126 40962 12178
rect 40962 12126 40964 12178
rect 40908 12124 40964 12126
rect 39788 11228 39844 11284
rect 39452 10668 39508 10724
rect 39340 10220 39396 10276
rect 39676 10610 39732 10612
rect 39676 10558 39678 10610
rect 39678 10558 39730 10610
rect 39730 10558 39732 10610
rect 39676 10556 39732 10558
rect 40012 10668 40068 10724
rect 41468 11282 41524 11284
rect 41468 11230 41470 11282
rect 41470 11230 41522 11282
rect 41522 11230 41524 11282
rect 41468 11228 41524 11230
rect 44492 20748 44548 20804
rect 44380 19516 44436 19572
rect 44212 18450 44268 18452
rect 44212 18398 44214 18450
rect 44214 18398 44266 18450
rect 44266 18398 44268 18450
rect 44212 18396 44268 18398
rect 44380 16268 44436 16324
rect 44212 16210 44268 16212
rect 44212 16158 44214 16210
rect 44214 16158 44266 16210
rect 44266 16158 44268 16210
rect 44212 16156 44268 16158
rect 43596 14812 43652 14868
rect 44100 14306 44156 14308
rect 44100 14254 44102 14306
rect 44102 14254 44154 14306
rect 44154 14254 44156 14306
rect 44100 14252 44156 14254
rect 43484 14140 43540 14196
rect 43484 13804 43540 13860
rect 43484 13468 43540 13524
rect 43652 13356 43708 13412
rect 41692 12178 41748 12180
rect 41692 12126 41694 12178
rect 41694 12126 41746 12178
rect 41746 12126 41748 12178
rect 41692 12124 41748 12126
rect 41711 11788 41767 11844
rect 44380 12796 44436 12852
rect 43260 11788 43316 11844
rect 43932 12124 43988 12180
rect 43932 11618 43988 11620
rect 43932 11566 43934 11618
rect 43934 11566 43986 11618
rect 43986 11566 43988 11618
rect 43932 11564 43988 11566
rect 41020 10668 41076 10724
rect 41244 10610 41300 10612
rect 41244 10558 41246 10610
rect 41246 10558 41298 10610
rect 41298 10558 41300 10610
rect 41244 10556 41300 10558
rect 39228 8204 39284 8260
rect 39004 8092 39060 8148
rect 37996 7868 38052 7924
rect 37772 7644 37828 7700
rect 37996 7532 38052 7588
rect 39452 9660 39508 9716
rect 39900 9826 39956 9828
rect 39900 9774 39902 9826
rect 39902 9774 39954 9826
rect 39954 9774 39956 9826
rect 39900 9772 39956 9774
rect 39452 9042 39508 9044
rect 39452 8990 39454 9042
rect 39454 8990 39506 9042
rect 39506 8990 39508 9042
rect 39452 8988 39508 8990
rect 39900 8428 39956 8484
rect 39788 8258 39844 8260
rect 39788 8206 39790 8258
rect 39790 8206 39842 8258
rect 39842 8206 39844 8258
rect 39788 8204 39844 8206
rect 39564 7868 39620 7924
rect 37884 7308 37940 7364
rect 38444 7362 38500 7364
rect 38444 7310 38446 7362
rect 38446 7310 38498 7362
rect 38498 7310 38500 7362
rect 38444 7308 38500 7310
rect 37660 7196 37716 7252
rect 37548 6860 37604 6916
rect 40180 9772 40236 9828
rect 40460 9660 40516 9716
rect 40348 9212 40404 9268
rect 42588 9714 42644 9716
rect 42588 9662 42590 9714
rect 42590 9662 42642 9714
rect 42642 9662 42644 9714
rect 42588 9660 42644 9662
rect 41020 8930 41076 8932
rect 41020 8878 41022 8930
rect 41022 8878 41074 8930
rect 41074 8878 41076 8930
rect 41020 8876 41076 8878
rect 40684 8428 40740 8484
rect 40908 8204 40964 8260
rect 41692 8034 41748 8036
rect 41692 7982 41694 8034
rect 41694 7982 41746 8034
rect 41746 7982 41748 8034
rect 41692 7980 41748 7982
rect 42252 7474 42308 7476
rect 42252 7422 42254 7474
rect 42254 7422 42306 7474
rect 42306 7422 42308 7474
rect 42252 7420 42308 7422
rect 40124 7196 40180 7252
rect 43540 11394 43596 11396
rect 43540 11342 43542 11394
rect 43542 11342 43594 11394
rect 43594 11342 43596 11394
rect 43540 11340 43596 11342
rect 42980 11170 43036 11172
rect 42980 11118 42982 11170
rect 42982 11118 43034 11170
rect 43034 11118 43036 11170
rect 42980 11116 43036 11118
rect 43932 10610 43988 10612
rect 43932 10558 43934 10610
rect 43934 10558 43986 10610
rect 43986 10558 43988 10610
rect 43932 10556 43988 10558
rect 43820 10108 43876 10164
rect 42924 9660 42980 9716
rect 44268 11394 44324 11396
rect 44268 11342 44270 11394
rect 44270 11342 44322 11394
rect 44322 11342 44324 11394
rect 44268 11340 44324 11342
rect 44380 11116 44436 11172
rect 43932 9602 43988 9604
rect 43932 9550 43934 9602
rect 43934 9550 43986 9602
rect 43986 9550 43988 9602
rect 43932 9548 43988 9550
rect 44268 9436 44324 9492
rect 43092 8988 43148 9044
rect 43708 9042 43764 9044
rect 43708 8990 43710 9042
rect 43710 8990 43762 9042
rect 43762 8990 43764 9042
rect 43708 8988 43764 8990
rect 42812 7532 42868 7588
rect 43820 8876 43876 8932
rect 43820 7437 43822 7476
rect 43822 7437 43874 7476
rect 43874 7437 43876 7476
rect 43820 7420 43876 7437
rect 42924 7308 42980 7364
rect 43708 7362 43764 7364
rect 43708 7310 43710 7362
rect 43710 7310 43762 7362
rect 43762 7310 43764 7362
rect 43708 7308 43764 7310
rect 38892 6860 38948 6916
rect 37660 6524 37716 6580
rect 39228 6636 39284 6692
rect 38780 5740 38836 5796
rect 38892 5852 38948 5908
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 37660 5122 37716 5124
rect 37660 5070 37662 5122
rect 37662 5070 37714 5122
rect 37714 5070 37716 5122
rect 37660 5068 37716 5070
rect 38780 5068 38836 5124
rect 38500 4844 38556 4900
rect 37231 4508 37287 4564
rect 38332 4172 38388 4228
rect 38556 4284 38612 4340
rect 41356 6578 41412 6580
rect 41356 6526 41358 6578
rect 41358 6526 41410 6578
rect 41410 6526 41412 6578
rect 41356 6524 41412 6526
rect 43036 6524 43092 6580
rect 40124 6466 40180 6468
rect 40124 6414 40126 6466
rect 40126 6414 40178 6466
rect 40178 6414 40180 6466
rect 40124 6412 40180 6414
rect 39564 6188 39620 6244
rect 39340 5852 39396 5908
rect 39676 6076 39732 6132
rect 39116 4284 39172 4340
rect 40908 6076 40964 6132
rect 41692 5964 41748 6020
rect 41244 5869 41246 5908
rect 41246 5869 41298 5908
rect 41298 5869 41300 5908
rect 41244 5852 41300 5869
rect 40236 5740 40292 5796
rect 39900 5180 39956 5236
rect 40684 5122 40740 5124
rect 40684 5070 40686 5122
rect 40686 5070 40738 5122
rect 40738 5070 40740 5122
rect 40684 5068 40740 5070
rect 40348 4956 40404 5012
rect 40348 4338 40404 4340
rect 40348 4286 40350 4338
rect 40350 4286 40402 4338
rect 40402 4286 40404 4338
rect 40348 4284 40404 4286
rect 41356 4226 41412 4228
rect 41356 4174 41358 4226
rect 41358 4174 41410 4226
rect 41410 4174 41412 4226
rect 41356 4172 41412 4174
rect 42700 5794 42756 5796
rect 42700 5742 42702 5794
rect 42702 5742 42754 5794
rect 42754 5742 42756 5794
rect 42700 5740 42756 5742
rect 43148 6412 43204 6468
rect 43932 5346 43988 5348
rect 43932 5294 43934 5346
rect 43934 5294 43986 5346
rect 43986 5294 43988 5346
rect 43932 5292 43988 5294
rect 42140 4956 42196 5012
rect 42588 5010 42644 5012
rect 42588 4958 42590 5010
rect 42590 4958 42642 5010
rect 42642 4958 42644 5010
rect 42588 4956 42644 4958
rect 44268 6076 44324 6132
rect 44268 5404 44324 5460
rect 42140 3388 42196 3444
rect 43932 4172 43988 4228
rect 42700 3388 42756 3444
rect 36876 2716 36932 2772
<< metal3 >>
rect 45200 43092 46000 43120
rect 41682 43036 41692 43092
rect 41748 43036 46000 43092
rect 45200 43008 46000 43036
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 31602 41916 31612 41972
rect 31668 41916 33628 41972
rect 33684 41916 33694 41972
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 30930 41244 30940 41300
rect 30996 41244 33292 41300
rect 33348 41244 33358 41300
rect 24658 41132 24668 41188
rect 24724 41132 26012 41188
rect 26068 41132 26078 41188
rect 36418 41132 36428 41188
rect 36484 41132 37100 41188
rect 37156 41132 37772 41188
rect 37828 41132 37838 41188
rect 24770 41020 24780 41076
rect 24836 41020 25732 41076
rect 25788 41020 25798 41076
rect 39778 41020 39788 41076
rect 39844 41020 40516 41076
rect 40572 41020 40582 41076
rect 26226 40908 26236 40964
rect 26292 40908 28644 40964
rect 28700 40908 28710 40964
rect 36082 40908 36092 40964
rect 36148 40908 37996 40964
rect 38052 40908 38062 40964
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 35756 40684 36540 40740
rect 36596 40684 36606 40740
rect 31154 40572 31164 40628
rect 31220 40572 33180 40628
rect 33236 40572 33246 40628
rect 35756 40516 35812 40684
rect 36194 40572 36204 40628
rect 36260 40572 36876 40628
rect 36932 40572 37716 40628
rect 42018 40572 42028 40628
rect 42084 40572 42812 40628
rect 42868 40572 42878 40628
rect 32274 40460 32284 40516
rect 32340 40460 33423 40516
rect 33479 40460 35756 40516
rect 35812 40460 35822 40516
rect 37660 40404 37716 40572
rect 23202 40348 23212 40404
rect 23268 40348 23940 40404
rect 23996 40348 24006 40404
rect 25106 40348 25116 40404
rect 25172 40348 28812 40404
rect 28868 40348 28878 40404
rect 32386 40348 32396 40404
rect 32452 40348 33628 40404
rect 33684 40348 34300 40404
rect 34356 40348 34366 40404
rect 37650 40348 37660 40404
rect 37716 40348 38612 40404
rect 38668 40348 38678 40404
rect 39890 40348 39900 40404
rect 39956 40348 41020 40404
rect 41076 40348 41086 40404
rect 24434 40236 24444 40292
rect 24500 40236 25900 40292
rect 25956 40236 25966 40292
rect 27010 40236 27020 40292
rect 27076 40236 28364 40292
rect 28420 40236 28430 40292
rect 40114 40236 40124 40292
rect 40180 40236 41580 40292
rect 41636 40236 41646 40292
rect 23090 40124 23100 40180
rect 23156 40124 23436 40180
rect 23492 40124 23502 40180
rect 40002 40124 40012 40180
rect 40068 40124 41356 40180
rect 41412 40124 43484 40180
rect 43540 40124 43550 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 43026 39788 43036 39844
rect 43092 39788 43932 39844
rect 43988 39788 43998 39844
rect 45200 39732 46000 39760
rect 24322 39676 24332 39732
rect 24388 39676 27356 39732
rect 27412 39676 27422 39732
rect 39442 39676 39452 39732
rect 39508 39676 41356 39732
rect 41412 39676 41422 39732
rect 43362 39676 43372 39732
rect 43428 39676 46000 39732
rect 45200 39648 46000 39676
rect 20738 39564 20748 39620
rect 20804 39564 24108 39620
rect 24164 39564 27468 39620
rect 27524 39564 27534 39620
rect 29698 39564 29708 39620
rect 29764 39564 30268 39620
rect 30324 39564 30334 39620
rect 32834 39564 32844 39620
rect 32900 39564 33740 39620
rect 33796 39564 34524 39620
rect 34580 39564 34590 39620
rect 34962 39564 34972 39620
rect 35028 39564 36316 39620
rect 36372 39564 36988 39620
rect 37044 39564 37054 39620
rect 39554 39564 39564 39620
rect 39620 39564 41244 39620
rect 41300 39564 41310 39620
rect 22638 39452 22648 39508
rect 22704 39452 23548 39508
rect 23604 39452 23614 39508
rect 40572 39396 40628 39564
rect 40898 39452 40908 39508
rect 40964 39452 43260 39508
rect 43316 39452 43326 39508
rect 40562 39340 40572 39396
rect 40628 39340 40638 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 21522 39116 21532 39172
rect 21588 39116 22988 39172
rect 23044 39116 23054 39172
rect 31042 39004 31052 39060
rect 31108 39004 32396 39060
rect 32452 39004 32462 39060
rect 32946 39004 32956 39060
rect 33012 39004 33628 39060
rect 33684 39004 39452 39060
rect 39508 39004 39518 39060
rect 23426 38892 23436 38948
rect 23492 38892 24332 38948
rect 24388 38892 24398 38948
rect 19730 38780 19740 38836
rect 19796 38780 20748 38836
rect 20804 38780 20814 38836
rect 27458 38780 27468 38836
rect 27524 38780 28028 38836
rect 28084 38780 28700 38836
rect 28756 38780 29708 38836
rect 29764 38780 29774 38836
rect 31938 38780 31948 38836
rect 32004 38780 33124 38836
rect 33180 38780 33190 38836
rect 35074 38780 35084 38836
rect 35140 38780 35420 38836
rect 35476 38780 35486 38836
rect 39442 38780 39452 38836
rect 39508 38780 40908 38836
rect 40964 38780 40974 38836
rect 41346 38780 41356 38836
rect 41412 38780 43708 38836
rect 43764 38780 43774 38836
rect 20178 38668 20188 38724
rect 20244 38668 21868 38724
rect 21924 38668 21934 38724
rect 28354 38668 28364 38724
rect 28420 38668 29540 38724
rect 29596 38668 29606 38724
rect 31434 38668 31444 38724
rect 31500 38668 32060 38724
rect 32116 38668 32126 38724
rect 40002 38668 40012 38724
rect 40068 38668 41020 38724
rect 41076 38668 41580 38724
rect 41636 38668 41646 38724
rect 39330 38556 39340 38612
rect 39396 38556 39788 38612
rect 39844 38556 39854 38612
rect 40282 38556 40292 38612
rect 40348 38556 43372 38612
rect 43428 38556 43438 38612
rect 39788 38500 39844 38556
rect 39788 38444 41916 38500
rect 41972 38444 41982 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 33394 38220 33404 38276
rect 33460 38220 34188 38276
rect 34244 38220 34254 38276
rect 42914 38220 42924 38276
rect 42980 38220 43708 38276
rect 43764 38220 43774 38276
rect 24098 38108 24108 38164
rect 24164 38108 30828 38164
rect 30884 38108 31836 38164
rect 31892 38108 31902 38164
rect 20738 37996 20748 38052
rect 20804 37996 22988 38052
rect 23044 37996 23660 38052
rect 23716 37996 23828 38052
rect 23884 37996 23894 38052
rect 24434 37996 24444 38052
rect 24500 37996 25676 38052
rect 25732 37996 25742 38052
rect 26450 37996 26460 38052
rect 26516 37996 26964 38052
rect 27020 37996 27030 38052
rect 27234 37996 27244 38052
rect 27300 37996 27804 38052
rect 27860 37996 29260 38052
rect 29316 37996 29326 38052
rect 36530 37996 36540 38052
rect 36596 37996 37436 38052
rect 37492 37996 38668 38052
rect 38724 37996 38734 38052
rect 24444 37940 24500 37996
rect 23426 37884 23436 37940
rect 23492 37884 24500 37940
rect 24994 37884 25004 37940
rect 25060 37884 27468 37940
rect 27524 37884 29036 37940
rect 29092 37884 29102 37940
rect 34626 37884 34636 37940
rect 34692 37884 37100 37940
rect 37156 37884 37166 37940
rect 22306 37772 22316 37828
rect 22372 37772 26236 37828
rect 26292 37772 26302 37828
rect 27570 37772 27580 37828
rect 27636 37772 33628 37828
rect 33684 37772 33694 37828
rect 35858 37772 35868 37828
rect 35924 37772 36372 37828
rect 36428 37772 36438 37828
rect 31042 37660 31052 37716
rect 31108 37660 31118 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 21970 37548 21980 37604
rect 22036 37548 23940 37604
rect 23996 37548 24006 37604
rect 20178 37324 20188 37380
rect 20244 37324 21532 37380
rect 21588 37324 22652 37380
rect 22708 37324 22718 37380
rect 22306 37212 22316 37268
rect 22372 37212 23100 37268
rect 23156 37212 23436 37268
rect 23492 37212 23502 37268
rect 27402 37212 27412 37268
rect 27468 37212 30828 37268
rect 30884 37212 30894 37268
rect 20626 37100 20636 37156
rect 20692 37100 21644 37156
rect 21700 37100 22876 37156
rect 22932 37100 22942 37156
rect 26226 37100 26236 37156
rect 26292 37100 30716 37156
rect 30772 37100 30782 37156
rect 31052 37044 31108 37660
rect 33170 37548 33180 37604
rect 33236 37548 34412 37604
rect 34468 37548 34860 37604
rect 34916 37548 34926 37604
rect 32162 37436 32172 37492
rect 32228 37436 33124 37492
rect 31490 37100 31500 37156
rect 31556 37100 32900 37156
rect 20514 36988 20524 37044
rect 20580 36988 21868 37044
rect 21924 36988 21934 37044
rect 22642 36988 22652 37044
rect 22708 36988 24108 37044
rect 24164 36988 24174 37044
rect 26338 36988 26348 37044
rect 26404 36988 26852 37044
rect 26908 36988 26918 37044
rect 31052 36988 32340 37044
rect 32396 36988 32406 37044
rect 27020 36876 27132 36932
rect 27188 36876 27198 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 22138 36540 22148 36596
rect 22204 36540 22988 36596
rect 23044 36540 23054 36596
rect 27020 36484 27076 36876
rect 32844 36820 32900 37100
rect 33068 37044 33124 37436
rect 33506 37212 33516 37268
rect 33572 37212 34524 37268
rect 34580 37212 35868 37268
rect 35924 37212 35934 37268
rect 36530 37212 36540 37268
rect 36596 37212 37436 37268
rect 37492 37212 37884 37268
rect 37940 37212 37950 37268
rect 38210 37212 38220 37268
rect 38276 37212 39228 37268
rect 39284 37212 41468 37268
rect 41524 37212 41534 37268
rect 41682 37212 41692 37268
rect 41748 37212 43036 37268
rect 43092 37212 43102 37268
rect 36194 37100 36204 37156
rect 36260 37100 37212 37156
rect 37268 37100 37278 37156
rect 36988 37044 37044 37100
rect 33068 36988 33852 37044
rect 33908 36988 33918 37044
rect 34290 36988 34300 37044
rect 34356 36988 35532 37044
rect 35588 36988 36092 37044
rect 36148 36988 36652 37044
rect 36708 36988 36718 37044
rect 36978 36988 36988 37044
rect 37044 36988 37054 37044
rect 37538 36988 37548 37044
rect 37604 36988 39340 37044
rect 39396 36988 39900 37044
rect 39956 36988 39966 37044
rect 33068 36932 33124 36988
rect 33058 36876 33068 36932
rect 33124 36876 33134 36932
rect 42018 36876 42028 36932
rect 42084 36876 43596 36932
rect 43652 36876 43662 36932
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 32844 36764 33180 36820
rect 33236 36764 33246 36820
rect 33730 36652 33740 36708
rect 33796 36652 34860 36708
rect 34916 36652 34926 36708
rect 38612 36652 40460 36708
rect 40516 36652 40526 36708
rect 38612 36596 38668 36652
rect 34290 36540 34300 36596
rect 34356 36540 34524 36596
rect 34580 36540 34590 36596
rect 35074 36540 35084 36596
rect 35140 36540 37996 36596
rect 38052 36540 38668 36596
rect 21746 36428 21756 36484
rect 21812 36428 21980 36484
rect 22036 36428 22764 36484
rect 22820 36428 22830 36484
rect 27010 36428 27020 36484
rect 27076 36428 27086 36484
rect 30258 36428 30268 36484
rect 30324 36428 30548 36484
rect 30604 36428 30614 36484
rect 31042 36428 31052 36484
rect 31108 36428 31668 36484
rect 31724 36428 41020 36484
rect 41076 36428 41086 36484
rect 45200 36372 46000 36400
rect 21858 36316 21868 36372
rect 21924 36316 23268 36372
rect 23324 36316 23334 36372
rect 33506 36316 33516 36372
rect 33572 36316 35196 36372
rect 35252 36316 35262 36372
rect 39778 36316 39788 36372
rect 39844 36316 40516 36372
rect 40572 36316 40582 36372
rect 43138 36316 43148 36372
rect 43204 36316 46000 36372
rect 33852 36260 33908 36316
rect 45200 36288 46000 36316
rect 33842 36204 33852 36260
rect 33908 36204 33918 36260
rect 34374 36204 34412 36260
rect 34468 36204 34478 36260
rect 29586 36092 29596 36148
rect 29652 36092 32956 36148
rect 33012 36092 37884 36148
rect 37940 36092 37950 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 34682 35980 34692 36036
rect 34748 35980 42028 36036
rect 42084 35980 42094 36036
rect 25946 35868 25956 35924
rect 26012 35868 26908 35924
rect 26964 35868 26974 35924
rect 32162 35868 32172 35924
rect 32228 35868 34412 35924
rect 34468 35868 34478 35924
rect 43138 35868 43148 35924
rect 43204 35868 43820 35924
rect 43876 35868 43886 35924
rect 26618 35756 26628 35812
rect 26684 35756 29036 35812
rect 29092 35756 29102 35812
rect 31826 35756 31836 35812
rect 31892 35756 33068 35812
rect 33124 35756 33134 35812
rect 34682 35756 34692 35812
rect 34748 35756 40012 35812
rect 40068 35756 40078 35812
rect 10414 35644 10424 35700
rect 10480 35644 11116 35700
rect 11172 35644 12572 35700
rect 12628 35644 12638 35700
rect 23426 35644 23436 35700
rect 23492 35644 25676 35700
rect 25732 35644 26124 35700
rect 26180 35644 26190 35700
rect 27682 35644 27692 35700
rect 27748 35644 29372 35700
rect 29428 35644 29438 35700
rect 30706 35644 30716 35700
rect 30772 35644 32060 35700
rect 32116 35644 32126 35700
rect 32386 35644 32396 35700
rect 32452 35644 35476 35700
rect 35532 35644 35542 35700
rect 40898 35644 40908 35700
rect 40964 35644 43540 35700
rect 43484 35588 43540 35644
rect 27906 35532 27916 35588
rect 27972 35532 27982 35588
rect 30258 35532 30268 35588
rect 30324 35532 31052 35588
rect 31108 35532 31500 35588
rect 31556 35532 32172 35588
rect 32228 35532 32238 35588
rect 33450 35532 33460 35588
rect 33516 35532 33964 35588
rect 34020 35532 35588 35588
rect 39442 35532 39452 35588
rect 39508 35532 41580 35588
rect 41636 35532 41646 35588
rect 43474 35532 43484 35588
rect 43540 35532 43550 35588
rect 27916 35476 27972 35532
rect 35532 35476 35588 35532
rect 27916 35420 28196 35476
rect 32386 35420 32396 35476
rect 32452 35420 34132 35476
rect 34188 35420 34972 35476
rect 35028 35420 35038 35476
rect 35522 35420 35532 35476
rect 35588 35420 35598 35476
rect 35914 35420 35924 35476
rect 35980 35420 37044 35476
rect 37100 35420 37110 35476
rect 10322 35308 10332 35364
rect 10388 35308 11695 35364
rect 11751 35308 11761 35364
rect 21410 35308 21420 35364
rect 21476 35308 22092 35364
rect 22148 35308 22158 35364
rect 23258 35308 23268 35364
rect 23324 35308 25116 35364
rect 25172 35308 25676 35364
rect 25732 35308 25956 35364
rect 26012 35308 26022 35364
rect 26898 35308 26908 35364
rect 26964 35308 27972 35364
rect 28028 35308 28038 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 10994 35196 11004 35252
rect 11060 35196 11452 35252
rect 11508 35196 11518 35252
rect 28140 35140 28196 35420
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 41346 35196 41356 35252
rect 41412 35196 41422 35252
rect 9090 35084 9100 35140
rect 9156 35084 12012 35140
rect 12068 35084 13356 35140
rect 13412 35084 13422 35140
rect 28140 35084 35756 35140
rect 35812 35084 35822 35140
rect 37090 34972 37100 35028
rect 37156 34972 37324 35028
rect 37380 34972 37390 35028
rect 40226 34972 40236 35028
rect 40292 34972 40684 35028
rect 40740 34972 40750 35028
rect 17378 34860 17388 34916
rect 17444 34860 18620 34916
rect 18676 34860 18686 34916
rect 33058 34860 33068 34916
rect 33124 34860 34300 34916
rect 34356 34860 34366 34916
rect 41356 34804 41412 35196
rect 27010 34748 27020 34804
rect 27076 34748 28028 34804
rect 28084 34748 28094 34804
rect 40338 34748 40348 34804
rect 40404 34748 42588 34804
rect 42644 34748 42654 34804
rect 13010 34636 13020 34692
rect 13076 34636 13692 34692
rect 13748 34636 13758 34692
rect 30482 34636 30492 34692
rect 30548 34636 31220 34692
rect 31276 34636 31948 34692
rect 32004 34636 32014 34692
rect 10994 34524 11004 34580
rect 11060 34524 11788 34580
rect 11844 34524 11854 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 37202 34300 37212 34356
rect 37268 34300 37278 34356
rect 37212 34244 37268 34300
rect 28242 34188 28252 34244
rect 28308 34188 30380 34244
rect 30436 34188 32172 34244
rect 32228 34188 37884 34244
rect 37940 34188 37950 34244
rect 40114 34188 40124 34244
rect 40180 34188 41580 34244
rect 41636 34188 41646 34244
rect 9884 34076 10668 34132
rect 10724 34076 10734 34132
rect 10994 34076 11004 34132
rect 11060 34076 13020 34132
rect 13076 34076 13086 34132
rect 24546 34076 24556 34132
rect 24612 34076 25452 34132
rect 25508 34076 25518 34132
rect 33506 34076 33516 34132
rect 33572 34076 34636 34132
rect 34692 34076 34702 34132
rect 37202 34076 37212 34132
rect 37268 34076 37436 34132
rect 37492 34076 37502 34132
rect 39778 34076 39788 34132
rect 39844 34076 40796 34132
rect 40852 34076 40862 34132
rect 9884 33908 9940 34076
rect 9874 33852 9884 33908
rect 9940 33852 9950 33908
rect 35074 33852 35084 33908
rect 35140 33852 37324 33908
rect 37380 33852 37390 33908
rect 11106 33740 11116 33796
rect 11172 33740 12292 33796
rect 12348 33740 12358 33796
rect 14018 33740 14028 33796
rect 14084 33740 14812 33796
rect 14868 33740 18172 33796
rect 18228 33740 18238 33796
rect 24742 33740 24780 33796
rect 24836 33740 24846 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 13122 33628 13132 33684
rect 13188 33628 15820 33684
rect 15876 33628 17276 33684
rect 17332 33628 17342 33684
rect 24210 33628 24220 33684
rect 24276 33628 25284 33684
rect 25340 33628 25350 33684
rect 38322 33628 38332 33684
rect 38388 33628 39004 33684
rect 39060 33628 39070 33684
rect 16762 33516 16772 33572
rect 16828 33516 18284 33572
rect 18340 33516 18350 33572
rect 32386 33516 32396 33572
rect 32452 33516 35084 33572
rect 35140 33516 35150 33572
rect 36754 33516 36764 33572
rect 36820 33516 37884 33572
rect 37940 33516 37950 33572
rect 9762 33404 9772 33460
rect 9828 33404 11788 33460
rect 11844 33404 11854 33460
rect 12898 33404 12908 33460
rect 12964 33404 16156 33460
rect 16212 33404 17780 33460
rect 25442 33404 25452 33460
rect 25508 33404 26124 33460
rect 26180 33404 28476 33460
rect 28532 33404 28542 33460
rect 31490 33404 31500 33460
rect 31556 33404 32284 33460
rect 32340 33404 32350 33460
rect 36978 33404 36988 33460
rect 37044 33404 37548 33460
rect 37604 33404 37614 33460
rect 17724 33348 17780 33404
rect 6066 33292 6076 33348
rect 6132 33292 8652 33348
rect 8708 33292 9100 33348
rect 9156 33292 9166 33348
rect 15922 33292 15932 33348
rect 15988 33292 17052 33348
rect 17108 33292 17118 33348
rect 17724 33292 18396 33348
rect 18452 33292 18462 33348
rect 24434 33292 24444 33348
rect 24500 33292 27448 33348
rect 27504 33292 27514 33348
rect 28578 33292 28588 33348
rect 28644 33292 29484 33348
rect 29540 33292 29550 33348
rect 30034 33292 30044 33348
rect 30100 33292 31276 33348
rect 31332 33292 31948 33348
rect 32004 33292 32014 33348
rect 34962 33292 34972 33348
rect 35028 33292 38108 33348
rect 38164 33292 38892 33348
rect 38948 33292 39452 33348
rect 39508 33292 39788 33348
rect 39844 33292 39854 33348
rect 12450 33180 12460 33236
rect 12516 33180 18172 33236
rect 18228 33180 18238 33236
rect 34738 33180 34748 33236
rect 34804 33180 37044 33236
rect 37100 33180 37110 33236
rect 17938 33068 17948 33124
rect 18004 33068 19964 33124
rect 20020 33068 20748 33124
rect 20804 33068 20814 33124
rect 24658 33068 24668 33124
rect 24724 33068 26572 33124
rect 26628 33068 29260 33124
rect 29316 33068 29326 33124
rect 34402 33068 34412 33124
rect 34468 33068 36484 33124
rect 36540 33068 36550 33124
rect 45200 33012 46000 33040
rect 24770 32956 24780 33012
rect 24836 32956 25004 33012
rect 25060 32956 25070 33012
rect 36642 32956 36652 33012
rect 36708 32956 37996 33012
rect 38052 32956 38062 33012
rect 43138 32956 43148 33012
rect 43204 32956 46000 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 45200 32928 46000 32956
rect 34570 32844 34580 32900
rect 34636 32844 35644 32900
rect 35700 32844 35710 32900
rect 38826 32732 38836 32788
rect 38892 32732 40236 32788
rect 40292 32732 40302 32788
rect 16594 32620 16604 32676
rect 16660 32620 17724 32676
rect 17780 32620 19292 32676
rect 19348 32620 19358 32676
rect 31042 32620 31052 32676
rect 31108 32620 31836 32676
rect 31892 32620 31902 32676
rect 34010 32620 34020 32676
rect 34076 32620 35532 32676
rect 35588 32620 35598 32676
rect 9650 32508 9660 32564
rect 9716 32508 10332 32564
rect 10388 32508 10398 32564
rect 18162 32508 18172 32564
rect 18228 32508 21644 32564
rect 21700 32508 21710 32564
rect 24322 32508 24332 32564
rect 24388 32508 24892 32564
rect 24948 32508 24958 32564
rect 28354 32508 28364 32564
rect 28420 32508 28588 32564
rect 28644 32508 29036 32564
rect 29092 32508 29102 32564
rect 30594 32508 30604 32564
rect 30660 32508 31724 32564
rect 31780 32508 31790 32564
rect 35634 32508 35644 32564
rect 35700 32508 38668 32564
rect 38724 32508 38734 32564
rect 26450 32396 26460 32452
rect 26516 32396 28868 32452
rect 28924 32396 28934 32452
rect 35186 32396 35196 32452
rect 35252 32396 35644 32452
rect 35700 32396 35710 32452
rect 8306 32284 8316 32340
rect 8372 32284 12460 32340
rect 12516 32284 12526 32340
rect 15026 32284 15036 32340
rect 15092 32284 17444 32340
rect 17500 32284 17510 32340
rect 30454 32284 30492 32340
rect 30548 32284 30558 32340
rect 31972 32284 31982 32340
rect 32038 32284 32956 32340
rect 33012 32284 33404 32340
rect 33460 32284 33470 32340
rect 34290 32284 34300 32340
rect 34356 32284 35868 32340
rect 35924 32284 35934 32340
rect 30594 32172 30604 32228
rect 30660 32172 30670 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 24714 31836 24724 31892
rect 24780 31836 27692 31892
rect 27748 31836 27758 31892
rect 27906 31836 27916 31892
rect 27972 31836 29652 31892
rect 29708 31836 29718 31892
rect 15586 31724 15596 31780
rect 15652 31724 16268 31780
rect 16324 31724 17612 31780
rect 17668 31724 17678 31780
rect 19618 31724 19628 31780
rect 19684 31724 21980 31780
rect 22036 31724 22046 31780
rect 23538 31724 23548 31780
rect 23604 31724 25452 31780
rect 25508 31724 25788 31780
rect 25844 31724 25854 31780
rect 26852 31724 27804 31780
rect 27860 31724 29484 31780
rect 29540 31724 29550 31780
rect 26852 31668 26908 31724
rect 30604 31668 30660 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 32386 32060 32396 32116
rect 32452 32060 34300 32116
rect 34356 32060 35028 32116
rect 34972 32004 35028 32060
rect 34972 31948 35756 32004
rect 35812 31948 35822 32004
rect 33730 31836 33740 31892
rect 33796 31836 34860 31892
rect 34916 31836 34926 31892
rect 35308 31836 35980 31892
rect 36036 31836 36046 31892
rect 42242 31836 42252 31892
rect 42308 31836 43260 31892
rect 43316 31836 43326 31892
rect 35308 31780 35364 31836
rect 31266 31724 31276 31780
rect 31332 31724 31948 31780
rect 32004 31724 32172 31780
rect 32228 31724 32238 31780
rect 35298 31724 35308 31780
rect 35364 31724 35374 31780
rect 35606 31724 35644 31780
rect 35700 31724 35710 31780
rect 38098 31724 38108 31780
rect 38164 31724 39564 31780
rect 39620 31724 39630 31780
rect 26002 31612 26012 31668
rect 26068 31612 26908 31668
rect 30258 31612 30268 31668
rect 30324 31612 30660 31668
rect 26226 31500 26236 31556
rect 26292 31500 28028 31556
rect 28084 31500 29372 31556
rect 29428 31500 29438 31556
rect 24994 31388 25004 31444
rect 25060 31388 27244 31444
rect 27300 31388 27310 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 30268 31332 30324 31612
rect 25554 31276 25564 31332
rect 25620 31276 30324 31332
rect 28970 31164 28980 31220
rect 29036 31164 31144 31220
rect 31200 31164 31210 31220
rect 28130 31052 28140 31108
rect 28196 31052 29596 31108
rect 29652 31052 29662 31108
rect 30454 31052 30492 31108
rect 30548 31052 30558 31108
rect 31714 31052 31724 31108
rect 31780 31052 32732 31108
rect 32788 31052 34244 31108
rect 31724 30996 31780 31052
rect 34188 30996 34244 31052
rect 22866 30940 22876 30996
rect 22932 30940 27468 30996
rect 27524 30940 27534 30996
rect 28466 30940 28476 30996
rect 28532 30940 29260 30996
rect 29316 30940 29326 30996
rect 31098 30940 31108 30996
rect 31164 30940 31780 30996
rect 32274 30940 32284 30996
rect 32340 30940 33180 30996
rect 33236 30940 33246 30996
rect 33338 30940 33348 30996
rect 33404 30940 33852 30996
rect 33908 30940 33918 30996
rect 34178 30940 34188 30996
rect 34244 30940 35532 30996
rect 35588 30940 35598 30996
rect 23314 30828 23324 30884
rect 23380 30828 25228 30884
rect 25284 30828 25452 30884
rect 25508 30828 25518 30884
rect 27122 30828 27132 30884
rect 27188 30828 30156 30884
rect 30212 30828 30604 30884
rect 30660 30828 30670 30884
rect 30818 30828 30828 30884
rect 30884 30828 31836 30884
rect 31892 30828 32172 30884
rect 32228 30828 32238 30884
rect 26114 30716 26124 30772
rect 26180 30716 26348 30772
rect 26404 30716 27916 30772
rect 27972 30716 27982 30772
rect 33730 30716 33740 30772
rect 33796 30716 40012 30772
rect 40068 30716 40078 30772
rect 41906 30716 41916 30772
rect 41972 30716 42700 30772
rect 42756 30716 42766 30772
rect 16716 30604 17836 30660
rect 17892 30604 21980 30660
rect 22036 30604 22046 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 16716 30548 16772 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 13906 30492 13916 30548
rect 13972 30492 15148 30548
rect 15204 30492 15214 30548
rect 16706 30492 16716 30548
rect 16772 30492 16782 30548
rect 20066 30380 20076 30436
rect 20132 30380 20636 30436
rect 20692 30380 21196 30436
rect 21252 30380 21262 30436
rect 28074 30380 28084 30436
rect 28140 30380 30828 30436
rect 30884 30380 30894 30436
rect 32722 30380 32732 30436
rect 32788 30380 33516 30436
rect 33572 30380 33582 30436
rect 17714 30268 17724 30324
rect 17780 30268 18676 30324
rect 40450 30268 40460 30324
rect 40516 30268 42924 30324
rect 42980 30268 42990 30324
rect 14802 30156 14812 30212
rect 14868 30156 16044 30212
rect 16100 30156 16110 30212
rect 18620 29988 18676 30268
rect 19898 30156 19908 30212
rect 19964 30156 21644 30212
rect 21700 30156 21710 30212
rect 23874 30156 23884 30212
rect 23940 30156 25228 30212
rect 25284 30156 25294 30212
rect 25778 30156 25788 30212
rect 25844 30156 26460 30212
rect 26516 30156 26796 30212
rect 26852 30156 27244 30212
rect 27300 30156 27310 30212
rect 31602 30156 31612 30212
rect 31668 30156 33068 30212
rect 33124 30156 33134 30212
rect 24994 30044 25004 30100
rect 25060 30044 26572 30100
rect 26628 30044 26638 30100
rect 18610 29932 18620 29988
rect 18676 29932 18686 29988
rect 23538 29932 23548 29988
rect 23604 29932 24556 29988
rect 24612 29932 24622 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 45200 29652 46000 29680
rect 43362 29596 43372 29652
rect 43428 29596 46000 29652
rect 45200 29568 46000 29596
rect 19730 29484 19740 29540
rect 19796 29484 20300 29540
rect 20356 29484 20366 29540
rect 23202 29372 23212 29428
rect 23268 29372 24220 29428
rect 24276 29372 24286 29428
rect 36866 29372 36876 29428
rect 36932 29372 37324 29428
rect 37380 29372 37390 29428
rect 17826 29260 17836 29316
rect 17892 29260 18956 29316
rect 19012 29260 25116 29316
rect 25172 29260 25182 29316
rect 36306 29260 36316 29316
rect 36372 29260 37212 29316
rect 37268 29260 37772 29316
rect 37828 29260 37838 29316
rect 39330 29260 39340 29316
rect 39396 29260 41244 29316
rect 41300 29260 41310 29316
rect 12674 29148 12684 29204
rect 12740 29148 13468 29204
rect 13524 29148 17052 29204
rect 17108 29148 17118 29204
rect 23874 29148 23884 29204
rect 23940 29148 24220 29204
rect 24276 29148 24286 29204
rect 15148 29092 15204 29148
rect 15138 29036 15148 29092
rect 15204 29036 15214 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 23660 28812 25004 28868
rect 25060 28812 25564 28868
rect 25620 28812 25630 28868
rect 41682 28812 41692 28868
rect 41748 28812 43596 28868
rect 43652 28812 43662 28868
rect 23202 28588 23212 28644
rect 23268 28588 23492 28644
rect 23436 28420 23492 28588
rect 23660 28532 23716 28812
rect 38658 28700 38668 28756
rect 38724 28700 41356 28756
rect 41412 28700 41422 28756
rect 24098 28588 24108 28644
rect 24164 28588 24444 28644
rect 24500 28588 24510 28644
rect 26786 28588 26796 28644
rect 26852 28588 27580 28644
rect 27636 28588 28812 28644
rect 28868 28588 28878 28644
rect 34514 28588 34524 28644
rect 34580 28588 35420 28644
rect 35476 28588 35486 28644
rect 36698 28588 36708 28644
rect 36764 28588 37884 28644
rect 37940 28588 37950 28644
rect 41234 28588 41244 28644
rect 41300 28588 43484 28644
rect 43540 28588 43550 28644
rect 23650 28476 23660 28532
rect 23716 28476 23726 28532
rect 29810 28476 29820 28532
rect 29876 28476 31052 28532
rect 31108 28476 31612 28532
rect 31668 28476 31678 28532
rect 35970 28476 35980 28532
rect 36036 28476 37212 28532
rect 37268 28476 37278 28532
rect 37426 28476 37436 28532
rect 37492 28476 38556 28532
rect 38612 28476 38622 28532
rect 20514 28364 20524 28420
rect 20580 28364 22204 28420
rect 22260 28364 22270 28420
rect 23436 28364 23548 28420
rect 23604 28364 23614 28420
rect 26450 28364 26460 28420
rect 26516 28364 27356 28420
rect 27412 28364 27422 28420
rect 29138 28364 29148 28420
rect 29204 28364 30828 28420
rect 30884 28364 31388 28420
rect 31444 28364 31454 28420
rect 36250 28364 36260 28420
rect 36316 28364 36652 28420
rect 36708 28364 36718 28420
rect 28018 28252 28028 28308
rect 28084 28252 30268 28308
rect 30324 28252 30334 28308
rect 36418 28252 36428 28308
rect 36484 28252 36876 28308
rect 36932 28252 36942 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 23090 28028 23100 28084
rect 23156 28028 23166 28084
rect 31154 28028 31164 28084
rect 31220 28028 32060 28084
rect 32116 28028 35756 28084
rect 35812 28028 35822 28084
rect 38882 28028 38892 28084
rect 38948 28028 41020 28084
rect 41076 28028 41086 28084
rect 23100 27860 23156 28028
rect 23762 27916 23772 27972
rect 23828 27916 25564 27972
rect 25620 27916 25630 27972
rect 10434 27804 10444 27860
rect 10500 27804 11788 27860
rect 11844 27804 12796 27860
rect 12852 27804 12862 27860
rect 21522 27804 21532 27860
rect 21588 27804 24724 27860
rect 24780 27804 24790 27860
rect 37538 27804 37548 27860
rect 37604 27804 39676 27860
rect 39732 27804 39742 27860
rect 25554 27468 25564 27524
rect 25620 27468 26348 27524
rect 26404 27468 26414 27524
rect 26562 27468 26572 27524
rect 26628 27468 27244 27524
rect 27300 27468 27310 27524
rect 35858 27468 35868 27524
rect 35924 27468 36988 27524
rect 37044 27468 37054 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 25106 27356 25116 27412
rect 25172 27356 25182 27412
rect 25666 27356 25676 27412
rect 25732 27356 26684 27412
rect 26740 27356 26750 27412
rect 14130 27244 14140 27300
rect 14196 27244 18844 27300
rect 18900 27244 18910 27300
rect 20850 27244 20860 27300
rect 20916 27244 22596 27300
rect 22652 27244 22662 27300
rect 25116 27188 25172 27356
rect 27346 27244 27356 27300
rect 27412 27244 28700 27300
rect 28756 27244 28766 27300
rect 32498 27244 32508 27300
rect 32564 27244 37996 27300
rect 38052 27244 41244 27300
rect 41300 27244 41310 27300
rect 41682 27244 41692 27300
rect 41748 27244 43708 27300
rect 14578 27132 14588 27188
rect 14644 27132 15596 27188
rect 15652 27132 15662 27188
rect 19058 27132 19068 27188
rect 19124 27132 20300 27188
rect 20356 27132 21308 27188
rect 21364 27132 21374 27188
rect 25116 27132 27804 27188
rect 27860 27132 27870 27188
rect 29642 27132 29652 27188
rect 29708 27132 30268 27188
rect 30324 27132 30334 27188
rect 31602 27132 31612 27188
rect 31668 27132 32172 27188
rect 32228 27132 32238 27188
rect 34066 27132 34076 27188
rect 34132 27132 36316 27188
rect 36372 27132 36876 27188
rect 36932 27132 36942 27188
rect 14466 27020 14476 27076
rect 14532 27020 15148 27076
rect 19842 27020 19852 27076
rect 19908 27020 20412 27076
rect 20468 27020 20860 27076
rect 20916 27020 20926 27076
rect 22642 27020 22652 27076
rect 22708 27020 23772 27076
rect 23828 27020 23838 27076
rect 15092 26964 15148 27020
rect 15092 26908 20524 26964
rect 20580 26908 20590 26964
rect 21522 26908 21532 26964
rect 21588 26908 22148 26964
rect 22204 26908 22214 26964
rect 25116 26852 25172 27132
rect 26338 27020 26348 27076
rect 26404 27020 27020 27076
rect 27076 27020 27086 27076
rect 33170 27020 33180 27076
rect 33236 27020 33628 27076
rect 33684 27020 33694 27076
rect 35084 27020 36652 27076
rect 36708 27020 36718 27076
rect 38546 27020 38556 27076
rect 38612 27020 39676 27076
rect 39732 27020 42140 27076
rect 42196 27020 42206 27076
rect 26002 26908 26012 26964
rect 26068 26908 26572 26964
rect 26628 26908 26638 26964
rect 29138 26908 29148 26964
rect 29204 26908 29708 26964
rect 29764 26908 29774 26964
rect 35084 26852 35140 27020
rect 36082 26908 36092 26964
rect 36148 26908 36988 26964
rect 37044 26908 37054 26964
rect 43652 26908 43708 27244
rect 43764 26908 43774 26964
rect 20402 26796 20412 26852
rect 20468 26796 21420 26852
rect 21476 26796 21486 26852
rect 25106 26796 25116 26852
rect 25172 26796 25182 26852
rect 35074 26796 35084 26852
rect 35140 26796 35150 26852
rect 20178 26684 20188 26740
rect 20244 26684 23884 26740
rect 23940 26684 23950 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 43810 26572 43820 26628
rect 43876 26572 44380 26628
rect 44436 26572 44446 26628
rect 20626 26460 20636 26516
rect 20692 26460 21756 26516
rect 21812 26460 22316 26516
rect 22372 26460 28588 26516
rect 28644 26460 29484 26516
rect 29540 26460 29550 26516
rect 37314 26348 37324 26404
rect 37380 26348 37772 26404
rect 37828 26348 38556 26404
rect 38612 26348 38622 26404
rect 44034 26348 44044 26404
rect 44100 26348 44110 26404
rect 10210 26236 10220 26292
rect 10276 26236 12684 26292
rect 12740 26236 17836 26292
rect 17892 26236 18732 26292
rect 18788 26236 18798 26292
rect 23090 26236 23100 26292
rect 23156 26236 23772 26292
rect 23828 26236 23838 26292
rect 33058 26236 33068 26292
rect 33124 26236 33628 26292
rect 33684 26236 33694 26292
rect 30930 26124 30940 26180
rect 30996 26124 37660 26180
rect 37716 26124 37726 26180
rect 29362 26012 29372 26068
rect 29428 26012 30604 26068
rect 30660 26012 30670 26068
rect 34738 26012 34748 26068
rect 34804 26012 38668 26068
rect 20178 25900 20188 25956
rect 20244 25900 20792 25956
rect 20848 25900 20858 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 38612 25732 38668 26012
rect 44044 25956 44100 26348
rect 45200 26292 46000 26320
rect 44258 26236 44268 26292
rect 44324 26236 46000 26292
rect 45200 26208 46000 26236
rect 44044 25900 44156 25956
rect 44212 25900 44222 25956
rect 34626 25676 34636 25732
rect 34692 25676 37436 25732
rect 37492 25676 37502 25732
rect 38612 25676 40348 25732
rect 40404 25676 40414 25732
rect 20514 25564 20524 25620
rect 20580 25564 21980 25620
rect 22036 25564 22046 25620
rect 30706 25564 30716 25620
rect 30772 25564 32060 25620
rect 32116 25564 32126 25620
rect 37090 25564 37100 25620
rect 37156 25564 40796 25620
rect 40852 25564 40862 25620
rect 11106 25452 11116 25508
rect 11172 25452 13020 25508
rect 13076 25452 13086 25508
rect 27458 25452 27468 25508
rect 27524 25452 27804 25508
rect 27860 25452 27870 25508
rect 36530 25452 36540 25508
rect 36596 25452 37996 25508
rect 38052 25452 38062 25508
rect 40450 25452 40460 25508
rect 40516 25452 43820 25508
rect 43876 25452 44380 25508
rect 44436 25452 44446 25508
rect 12338 25340 12348 25396
rect 12404 25340 13356 25396
rect 13412 25340 13422 25396
rect 17826 25340 17836 25396
rect 17892 25340 20076 25396
rect 20132 25340 29764 25396
rect 29820 25340 29830 25396
rect 32498 25340 32508 25396
rect 32564 25340 34972 25396
rect 35028 25340 36988 25396
rect 37044 25340 37054 25396
rect 39890 25340 39900 25396
rect 39956 25340 40684 25396
rect 40740 25340 40750 25396
rect 40898 25340 40908 25396
rect 40964 25340 42700 25396
rect 42756 25340 42766 25396
rect 9874 25228 9884 25284
rect 9940 25228 10332 25284
rect 10388 25228 11228 25284
rect 11284 25228 11294 25284
rect 11442 25228 11452 25284
rect 11508 25228 12236 25284
rect 12292 25228 12302 25284
rect 19170 25228 19180 25284
rect 19236 25228 20188 25284
rect 20244 25228 20254 25284
rect 24770 25228 24780 25284
rect 24836 25228 25564 25284
rect 25620 25228 25630 25284
rect 26114 25228 26124 25284
rect 26180 25228 28476 25284
rect 28532 25228 28542 25284
rect 36306 25228 36316 25284
rect 36372 25228 37100 25284
rect 37156 25228 37166 25284
rect 37426 25228 37436 25284
rect 37492 25228 39788 25284
rect 39844 25228 39854 25284
rect 10882 25116 10892 25172
rect 10948 25116 17836 25172
rect 17892 25116 17902 25172
rect 25890 25116 25900 25172
rect 25956 25116 27468 25172
rect 27524 25116 27534 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 15138 25004 15148 25060
rect 15204 25004 16604 25060
rect 16660 25004 16670 25060
rect 39666 25004 39676 25060
rect 39732 25004 40684 25060
rect 40740 25004 40750 25060
rect 40226 24892 40236 24948
rect 40292 24892 41692 24948
rect 41748 24892 42364 24948
rect 42420 24892 42430 24948
rect 28634 24780 28644 24836
rect 28700 24780 31948 24836
rect 32004 24780 32014 24836
rect 16818 24668 16828 24724
rect 16884 24668 17276 24724
rect 17332 24668 17342 24724
rect 37538 24668 37548 24724
rect 37604 24668 39116 24724
rect 39172 24668 39182 24724
rect 39982 24668 39992 24724
rect 40048 24668 44380 24724
rect 44436 24668 44446 24724
rect 21634 24556 21644 24612
rect 21700 24556 23548 24612
rect 23604 24556 23614 24612
rect 23986 24444 23996 24500
rect 24052 24444 26460 24500
rect 26516 24444 29148 24500
rect 29204 24444 29214 24500
rect 43922 24444 43932 24500
rect 43988 24444 44492 24500
rect 44548 24444 44558 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 15698 24220 15708 24276
rect 15764 24220 16716 24276
rect 16772 24220 16782 24276
rect 32386 24108 32396 24164
rect 32452 24108 36092 24164
rect 36148 24108 36158 24164
rect 10266 23996 10276 24052
rect 10332 23996 10892 24052
rect 10948 23996 10958 24052
rect 14802 23996 14812 24052
rect 14868 23996 15596 24052
rect 15652 23996 15662 24052
rect 18050 23996 18060 24052
rect 18116 23996 18620 24052
rect 18676 23996 18686 24052
rect 24434 23996 24444 24052
rect 24500 23996 25340 24052
rect 25396 23996 25406 24052
rect 28690 23996 28700 24052
rect 28756 23996 29260 24052
rect 29316 23996 30156 24052
rect 30212 23996 30222 24052
rect 31042 23996 31052 24052
rect 31108 23996 33292 24052
rect 33348 23996 33358 24052
rect 33618 23996 33628 24052
rect 33684 23996 35980 24052
rect 36036 23996 36046 24052
rect 38210 23996 38220 24052
rect 38276 23996 41020 24052
rect 41076 23996 41086 24052
rect 14242 23884 14252 23940
rect 14308 23884 15708 23940
rect 15764 23884 15774 23940
rect 16258 23884 16268 23940
rect 16324 23884 17164 23940
rect 17220 23884 18956 23940
rect 19012 23884 19404 23940
rect 19460 23884 19470 23940
rect 19842 23884 19852 23940
rect 19908 23884 21644 23940
rect 21700 23884 21710 23940
rect 35522 23884 35532 23940
rect 35588 23884 36316 23940
rect 36372 23884 36382 23940
rect 39666 23884 39676 23940
rect 39732 23884 40236 23940
rect 40292 23884 40302 23940
rect 27234 23772 27244 23828
rect 27300 23772 27692 23828
rect 27748 23772 27758 23828
rect 26898 23660 26908 23716
rect 26964 23660 29148 23716
rect 29204 23660 29214 23716
rect 22642 23548 22652 23604
rect 22708 23548 25452 23604
rect 25508 23548 25518 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 24210 23436 24220 23492
rect 24276 23436 31388 23492
rect 31444 23436 31454 23492
rect 37538 23436 37548 23492
rect 37604 23436 38108 23492
rect 38164 23436 38174 23492
rect 41906 23436 41916 23492
rect 41972 23436 43372 23492
rect 43428 23436 43438 23492
rect 21858 23324 21868 23380
rect 21924 23324 28812 23380
rect 28868 23324 28878 23380
rect 32722 23324 32732 23380
rect 32788 23324 33572 23380
rect 33628 23324 33638 23380
rect 9874 23212 9884 23268
rect 9940 23212 10556 23268
rect 10612 23212 11676 23268
rect 11732 23212 11742 23268
rect 17938 23212 17948 23268
rect 18004 23212 21084 23268
rect 21140 23212 21308 23268
rect 21364 23212 21374 23268
rect 21634 23212 21644 23268
rect 21700 23212 29932 23268
rect 29988 23212 32172 23268
rect 32228 23212 32238 23268
rect 40450 23212 40460 23268
rect 40516 23212 43036 23268
rect 43092 23212 43820 23268
rect 43876 23212 43886 23268
rect 10882 23100 10892 23156
rect 10948 23100 12796 23156
rect 12852 23100 12862 23156
rect 14466 23100 14476 23156
rect 14532 23100 16156 23156
rect 16212 23100 16222 23156
rect 21186 23100 21196 23156
rect 21252 23100 21756 23156
rect 21812 23100 21822 23156
rect 29362 23100 29372 23156
rect 29428 23100 30808 23156
rect 30864 23100 30874 23156
rect 31490 23100 31500 23156
rect 31556 23100 32060 23156
rect 32116 23100 32126 23156
rect 32498 23100 32508 23156
rect 32564 23100 33292 23156
rect 33348 23100 34860 23156
rect 34916 23100 35532 23156
rect 35588 23100 35598 23156
rect 41346 23100 41356 23156
rect 41412 23100 43484 23156
rect 43540 23100 43550 23156
rect 10770 22988 10780 23044
rect 10836 22988 12572 23044
rect 12628 22988 12638 23044
rect 20850 22988 20860 23044
rect 20916 22988 21532 23044
rect 21588 22988 21598 23044
rect 25890 22988 25900 23044
rect 25956 22988 28308 23044
rect 28364 22988 28374 23044
rect 36978 22988 36988 23044
rect 37044 22988 37100 23044
rect 37156 22988 37166 23044
rect 45200 22932 46000 22960
rect 9762 22876 9772 22932
rect 9828 22876 12684 22932
rect 12740 22876 15148 22932
rect 15204 22876 15214 22932
rect 28802 22876 28812 22932
rect 28868 22876 31500 22932
rect 31556 22876 31566 22932
rect 35970 22876 35980 22932
rect 36036 22876 38556 22932
rect 38612 22876 38622 22932
rect 43036 22876 46000 22932
rect 43036 22820 43092 22876
rect 45200 22848 46000 22876
rect 13682 22764 13692 22820
rect 13748 22764 19628 22820
rect 19684 22764 19694 22820
rect 19861 22764 19871 22820
rect 19927 22764 20356 22820
rect 20412 22764 20422 22820
rect 27458 22764 27468 22820
rect 27524 22764 27692 22820
rect 27748 22764 27758 22820
rect 43026 22764 43036 22820
rect 43092 22764 43102 22820
rect 43558 22764 43596 22820
rect 43652 22764 43662 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 38098 22652 38108 22708
rect 38164 22652 38668 22708
rect 38724 22652 38734 22708
rect 38882 22652 38892 22708
rect 38948 22652 40572 22708
rect 40628 22652 42252 22708
rect 42308 22652 42318 22708
rect 23762 22540 23772 22596
rect 23828 22540 24444 22596
rect 24500 22540 25452 22596
rect 25508 22540 25518 22596
rect 29530 22540 29540 22596
rect 29596 22540 30808 22596
rect 30864 22540 30874 22596
rect 36194 22540 36204 22596
rect 36260 22540 38332 22596
rect 38388 22540 38398 22596
rect 38994 22540 39004 22596
rect 39060 22540 42924 22596
rect 42980 22540 42990 22596
rect 38210 22428 38220 22484
rect 38276 22428 38668 22484
rect 38724 22428 38734 22484
rect 12786 22316 12796 22372
rect 12852 22316 13580 22372
rect 13636 22316 13646 22372
rect 20738 22316 20748 22372
rect 20804 22316 21084 22372
rect 21140 22316 21644 22372
rect 21700 22316 21710 22372
rect 26674 22316 26684 22372
rect 26740 22316 28588 22372
rect 28644 22316 28654 22372
rect 29922 22316 29932 22372
rect 29988 22316 30604 22372
rect 30660 22316 31836 22372
rect 31892 22316 31902 22372
rect 33842 22316 33852 22372
rect 33908 22316 35084 22372
rect 35140 22316 35150 22372
rect 36950 22316 36988 22372
rect 37044 22316 37054 22372
rect 33282 22092 33292 22148
rect 33348 22092 33852 22148
rect 33908 22092 33918 22148
rect 29586 21980 29596 22036
rect 29652 21980 30044 22036
rect 30100 21980 32340 22036
rect 32396 21980 40012 22036
rect 40068 21980 40078 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 26338 21868 26348 21924
rect 26404 21868 26796 21924
rect 26852 21868 28364 21924
rect 28420 21868 29260 21924
rect 29316 21868 29326 21924
rect 15362 21756 15372 21812
rect 15428 21756 15438 21812
rect 15698 21756 15708 21812
rect 15764 21756 18396 21812
rect 18452 21756 19292 21812
rect 19348 21756 19358 21812
rect 19618 21756 19628 21812
rect 19684 21756 24556 21812
rect 24612 21756 24622 21812
rect 29754 21756 29764 21812
rect 29820 21756 31612 21812
rect 31668 21756 32956 21812
rect 33012 21756 33022 21812
rect 35634 21756 35644 21812
rect 35700 21756 35960 21812
rect 36016 21756 36026 21812
rect 37762 21756 37772 21812
rect 37828 21756 38556 21812
rect 38612 21756 39116 21812
rect 39172 21756 39182 21812
rect 15372 21700 15428 21756
rect 15372 21644 15932 21700
rect 15988 21644 15998 21700
rect 28690 21644 28700 21700
rect 28756 21644 32060 21700
rect 32116 21644 32126 21700
rect 42130 21644 42140 21700
rect 42196 21644 43484 21700
rect 43540 21644 43550 21700
rect 8250 21532 8260 21588
rect 8316 21532 9436 21588
rect 9492 21532 9502 21588
rect 16818 21532 16828 21588
rect 16884 21532 21308 21588
rect 21364 21532 21374 21588
rect 24098 21532 24108 21588
rect 24164 21532 24174 21588
rect 24322 21532 24332 21588
rect 24388 21532 26460 21588
rect 26516 21532 26526 21588
rect 29372 21532 30380 21588
rect 30436 21532 32172 21588
rect 32228 21532 34860 21588
rect 34916 21532 34926 21588
rect 39554 21532 39564 21588
rect 39620 21532 41132 21588
rect 41188 21532 41198 21588
rect 24108 21476 24164 21532
rect 29372 21476 29428 21532
rect 9650 21420 9660 21476
rect 9716 21420 12124 21476
rect 12180 21420 12190 21476
rect 14242 21420 14252 21476
rect 14308 21420 17108 21476
rect 24108 21420 25228 21476
rect 25284 21420 25294 21476
rect 29362 21420 29372 21476
rect 29428 21420 29438 21476
rect 17052 21364 17108 21420
rect 8978 21308 8988 21364
rect 9044 21308 16828 21364
rect 16884 21308 16894 21364
rect 17052 21308 19012 21364
rect 19068 21308 19078 21364
rect 30706 21308 30716 21364
rect 30772 21308 40124 21364
rect 40180 21308 40190 21364
rect 14466 21196 14476 21252
rect 14532 21196 21868 21252
rect 21924 21196 22148 21252
rect 22204 21196 22214 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 13438 21084 13448 21140
rect 13504 21084 15148 21140
rect 15698 21084 15708 21140
rect 15764 21084 15932 21140
rect 15988 21084 16940 21140
rect 16996 21084 17948 21140
rect 18004 21084 18014 21140
rect 32050 21084 32060 21140
rect 32116 21084 33740 21140
rect 33796 21084 33806 21140
rect 15092 20804 15148 21084
rect 15586 20972 15596 21028
rect 15652 20972 17612 21028
rect 17668 20972 17678 21028
rect 20197 20972 20207 21028
rect 20263 20972 25396 21028
rect 25452 20972 25462 21028
rect 20850 20860 20860 20916
rect 20916 20860 21402 20916
rect 21458 20860 21468 20916
rect 21634 20860 21644 20916
rect 21700 20860 22820 20916
rect 22876 20860 26684 20916
rect 26740 20860 26750 20916
rect 35186 20860 35196 20916
rect 35252 20860 35756 20916
rect 35812 20860 35822 20916
rect 12002 20748 12012 20804
rect 12068 20748 13580 20804
rect 13636 20748 13646 20804
rect 15092 20748 21756 20804
rect 21812 20748 21822 20804
rect 25106 20748 25116 20804
rect 25172 20748 27356 20804
rect 27412 20748 27692 20804
rect 27748 20748 27758 20804
rect 29698 20748 29708 20804
rect 29764 20748 30380 20804
rect 30436 20748 31724 20804
rect 31780 20748 31790 20804
rect 32498 20748 32508 20804
rect 32564 20748 32956 20804
rect 33012 20748 33516 20804
rect 33572 20748 33582 20804
rect 40114 20748 40124 20804
rect 40180 20748 41300 20804
rect 41356 20748 43148 20804
rect 43204 20748 44268 20804
rect 44324 20748 44492 20804
rect 44548 20748 44558 20804
rect 6290 20636 6300 20692
rect 6356 20636 8092 20692
rect 8148 20636 8158 20692
rect 38770 20636 38780 20692
rect 38836 20636 40796 20692
rect 40852 20636 40862 20692
rect 10210 20524 10220 20580
rect 10276 20524 12236 20580
rect 12292 20524 12302 20580
rect 18498 20524 18508 20580
rect 18564 20524 19292 20580
rect 19348 20524 19684 20580
rect 19740 20524 20916 20580
rect 31322 20524 31332 20580
rect 31444 20524 31454 20580
rect 33898 20524 33908 20580
rect 33964 20524 35644 20580
rect 35700 20524 35710 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 20860 20356 20916 20524
rect 26338 20412 26348 20468
rect 26404 20412 27468 20468
rect 27524 20412 28644 20468
rect 28700 20412 40124 20468
rect 40180 20412 40190 20468
rect 20860 20300 34748 20356
rect 34804 20300 35812 20356
rect 35868 20300 35878 20356
rect 19170 20188 19180 20244
rect 19236 20188 19246 20244
rect 19954 20188 19964 20244
rect 20020 20188 20524 20244
rect 20580 20188 20590 20244
rect 19180 20132 19236 20188
rect 8082 20076 8092 20132
rect 8148 20076 8764 20132
rect 8820 20076 8830 20132
rect 14802 20076 14812 20132
rect 14868 20076 15036 20132
rect 15092 20076 15102 20132
rect 15810 20076 15820 20132
rect 15876 20076 18396 20132
rect 18452 20076 19236 20132
rect 27122 20076 27132 20132
rect 27188 20076 28028 20132
rect 28084 20076 28924 20132
rect 28980 20076 29932 20132
rect 29988 20076 30492 20132
rect 30548 20076 30558 20132
rect 31612 20076 38444 20132
rect 38500 20076 38510 20132
rect 16724 19964 16734 20020
rect 16790 19964 17276 20020
rect 17332 19964 17342 20020
rect 24266 19964 24276 20020
rect 24332 19964 26348 20020
rect 26404 19964 26414 20020
rect 27010 19964 27020 20020
rect 27076 19964 28140 20020
rect 28196 19964 28206 20020
rect 29586 19964 29596 20020
rect 29652 19964 30716 20020
rect 30772 19964 30782 20020
rect 8026 19852 8036 19908
rect 8092 19852 8988 19908
rect 9044 19852 9054 19908
rect 30146 19852 30156 19908
rect 30212 19852 31388 19908
rect 31444 19852 31454 19908
rect 23482 19740 23492 19796
rect 23548 19740 23996 19796
rect 24052 19740 24724 19796
rect 24780 19740 29820 19796
rect 29876 19740 29886 19796
rect 31612 19684 31668 20076
rect 34066 19964 34076 20020
rect 34132 19964 35084 20020
rect 35140 19964 35150 20020
rect 35858 19964 35868 20020
rect 35924 19964 38668 20020
rect 38724 19964 38734 20020
rect 41850 19964 41860 20020
rect 41916 19964 43708 20020
rect 43764 19964 43774 20020
rect 35522 19852 35532 19908
rect 35588 19852 39564 19908
rect 39620 19852 40124 19908
rect 40180 19852 40190 19908
rect 42252 19852 44044 19908
rect 44100 19852 44110 19908
rect 32162 19740 32172 19796
rect 32228 19740 38668 19796
rect 40226 19740 40236 19796
rect 40292 19740 41132 19796
rect 41188 19740 41198 19796
rect 12542 19628 12552 19684
rect 12608 19628 15372 19684
rect 15428 19628 15988 19684
rect 16044 19628 16054 19684
rect 23650 19628 23660 19684
rect 23716 19628 24220 19684
rect 24276 19628 24286 19684
rect 28354 19628 28364 19684
rect 28420 19628 31668 19684
rect 38612 19684 38668 19740
rect 42252 19684 42308 19852
rect 43334 19740 43372 19796
rect 43428 19740 43438 19796
rect 38612 19628 42308 19684
rect 43484 19628 43596 19684
rect 43652 19628 43662 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 8418 19404 8428 19460
rect 8484 19404 9772 19460
rect 9828 19404 11004 19460
rect 11060 19404 11070 19460
rect 26852 19404 28812 19460
rect 28868 19404 28878 19460
rect 39760 19404 39770 19460
rect 39826 19404 40796 19460
rect 40852 19404 40862 19460
rect 26852 19348 26908 19404
rect 8754 19292 8764 19348
rect 8820 19292 11732 19348
rect 13794 19292 13804 19348
rect 13860 19292 15708 19348
rect 15764 19292 15774 19348
rect 21970 19292 21980 19348
rect 22036 19292 22820 19348
rect 22876 19292 24108 19348
rect 24164 19292 26908 19348
rect 35970 19292 35980 19348
rect 36036 19292 37156 19348
rect 37212 19292 37772 19348
rect 37828 19292 37838 19348
rect 38658 19292 38668 19348
rect 38724 19292 39508 19348
rect 40506 19292 40516 19348
rect 40572 19292 41804 19348
rect 41860 19292 43148 19348
rect 43204 19292 43214 19348
rect 11676 19236 11732 19292
rect 39452 19236 39508 19292
rect 8362 19180 8372 19236
rect 8428 19180 9436 19236
rect 9492 19180 9502 19236
rect 11666 19180 11676 19236
rect 11732 19180 11742 19236
rect 12674 19180 12684 19236
rect 12740 19180 13468 19236
rect 13524 19180 13534 19236
rect 21466 19180 21476 19236
rect 21532 19180 21756 19236
rect 21812 19180 21822 19236
rect 26898 19180 26908 19236
rect 26964 19180 30156 19236
rect 30212 19180 30222 19236
rect 36978 19180 36988 19236
rect 37044 19180 38780 19236
rect 38836 19180 38846 19236
rect 39442 19180 39452 19236
rect 39508 19180 40908 19236
rect 40964 19180 40974 19236
rect 43484 19124 43540 19628
rect 45200 19572 46000 19600
rect 43698 19516 43708 19572
rect 43764 19516 44380 19572
rect 44436 19516 46000 19572
rect 45200 19488 46000 19516
rect 12786 19068 12796 19124
rect 12852 19068 13804 19124
rect 13860 19068 13870 19124
rect 21298 19068 21308 19124
rect 21364 19068 22204 19124
rect 22260 19068 22270 19124
rect 40674 19068 40684 19124
rect 40740 19068 43148 19124
rect 43204 19068 43540 19124
rect 15922 18956 15932 19012
rect 15988 18956 16492 19012
rect 16548 18956 17108 19012
rect 17164 18956 33404 19012
rect 33460 18956 33740 19012
rect 33796 18956 34020 19012
rect 34076 18956 34086 19012
rect 28130 18844 28140 18900
rect 28196 18844 28700 18900
rect 28756 18844 28766 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 29250 18620 29260 18676
rect 29316 18620 30828 18676
rect 30884 18620 32060 18676
rect 32116 18620 32126 18676
rect 37650 18620 37660 18676
rect 37716 18620 37828 18676
rect 42690 18620 42700 18676
rect 42756 18620 43260 18676
rect 43316 18620 43484 18676
rect 43540 18620 43550 18676
rect 8306 18508 8316 18564
rect 8372 18508 10892 18564
rect 10948 18508 10958 18564
rect 19842 18508 19852 18564
rect 19908 18508 22540 18564
rect 22596 18508 22606 18564
rect 28242 18508 28252 18564
rect 28308 18508 28318 18564
rect 30706 18508 30716 18564
rect 30772 18508 31388 18564
rect 31444 18508 31454 18564
rect 31714 18508 31724 18564
rect 31780 18508 35868 18564
rect 35924 18508 36988 18564
rect 37044 18508 37054 18564
rect 28252 18452 28308 18508
rect 10210 18396 10220 18452
rect 10276 18396 12012 18452
rect 12068 18396 12348 18452
rect 12404 18396 12414 18452
rect 22866 18396 22876 18452
rect 22932 18396 23996 18452
rect 24052 18396 24062 18452
rect 24770 18396 24780 18452
rect 24836 18396 25452 18452
rect 25508 18396 25518 18452
rect 26562 18396 26572 18452
rect 26628 18396 27356 18452
rect 27412 18396 27422 18452
rect 27804 18396 28812 18452
rect 28868 18396 28878 18452
rect 36194 18396 36204 18452
rect 36260 18396 37548 18452
rect 37604 18396 37614 18452
rect 27804 18340 27860 18396
rect 37772 18340 37828 18620
rect 39330 18396 39340 18452
rect 39396 18396 39788 18452
rect 39844 18396 40796 18452
rect 40852 18396 40862 18452
rect 43026 18396 43036 18452
rect 43092 18396 43596 18452
rect 43652 18396 44212 18452
rect 44268 18396 44278 18452
rect 10434 18284 10444 18340
rect 10500 18284 11452 18340
rect 11508 18284 11518 18340
rect 23744 18284 23754 18340
rect 23810 18284 25116 18340
rect 25172 18284 25182 18340
rect 25778 18284 25788 18340
rect 25844 18284 26796 18340
rect 26852 18284 26862 18340
rect 27020 18284 27804 18340
rect 27860 18284 27870 18340
rect 28242 18284 28252 18340
rect 28308 18284 28700 18340
rect 28756 18284 29484 18340
rect 29540 18284 29550 18340
rect 35746 18284 35756 18340
rect 35812 18284 42812 18340
rect 42868 18284 42878 18340
rect 43586 18284 43596 18340
rect 43652 18284 43820 18340
rect 43876 18284 43886 18340
rect 27020 18228 27076 18284
rect 24490 18172 24500 18228
rect 24556 18172 26460 18228
rect 26516 18172 27076 18228
rect 27234 18172 27244 18228
rect 27300 18172 28140 18228
rect 28196 18172 28206 18228
rect 32386 18172 32396 18228
rect 32452 18172 38668 18228
rect 27244 18116 27300 18172
rect 38612 18116 38668 18172
rect 7970 18060 7980 18116
rect 8036 18060 9100 18116
rect 9156 18060 10108 18116
rect 10164 18060 10174 18116
rect 17714 18060 17724 18116
rect 17780 18060 18900 18116
rect 18956 18060 19628 18116
rect 19684 18060 24724 18116
rect 26562 18060 26572 18116
rect 26628 18060 27300 18116
rect 27570 18060 27580 18116
rect 27636 18060 29148 18116
rect 29204 18060 29214 18116
rect 35578 18060 35588 18116
rect 35644 18060 36764 18116
rect 36820 18060 36830 18116
rect 38612 18060 40684 18116
rect 40740 18060 40750 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 24668 18004 24724 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 22194 17948 22204 18004
rect 22260 17948 24444 18004
rect 24500 17948 24510 18004
rect 24668 17948 26908 18004
rect 27122 17948 27132 18004
rect 27188 17948 27916 18004
rect 27972 17948 31724 18004
rect 31780 17948 31790 18004
rect 26852 17892 26908 17948
rect 14130 17836 14140 17892
rect 14196 17836 15372 17892
rect 15428 17836 15438 17892
rect 24322 17836 24332 17892
rect 24388 17836 25452 17892
rect 25508 17836 26012 17892
rect 26068 17836 26078 17892
rect 26852 17836 34300 17892
rect 34356 17836 34366 17892
rect 34794 17836 34804 17892
rect 34860 17836 36316 17892
rect 36372 17836 36382 17892
rect 37202 17836 37212 17892
rect 37268 17836 38668 17892
rect 38724 17836 38734 17892
rect 8530 17724 8540 17780
rect 8596 17724 10220 17780
rect 10276 17724 11228 17780
rect 11284 17724 11620 17780
rect 21522 17724 21532 17780
rect 21588 17724 23660 17780
rect 23716 17724 23726 17780
rect 24546 17724 24556 17780
rect 24612 17724 25788 17780
rect 25844 17724 25854 17780
rect 31826 17724 31836 17780
rect 31892 17724 33852 17780
rect 33908 17724 34972 17780
rect 35028 17724 35038 17780
rect 42802 17724 42812 17780
rect 42868 17724 43932 17780
rect 43988 17724 43998 17780
rect 11564 17668 11620 17724
rect 11554 17612 11564 17668
rect 11620 17612 11630 17668
rect 14334 17612 14344 17668
rect 14400 17612 18172 17668
rect 18228 17612 18508 17668
rect 18564 17612 18574 17668
rect 19394 17612 19404 17668
rect 19460 17612 19470 17668
rect 20850 17612 20860 17668
rect 20916 17612 23118 17668
rect 23174 17612 23184 17668
rect 24098 17612 24108 17668
rect 24164 17612 26124 17668
rect 26180 17612 26190 17668
rect 29586 17612 29596 17668
rect 29652 17612 30380 17668
rect 30436 17612 30446 17668
rect 30538 17612 30548 17668
rect 30604 17612 32844 17668
rect 32900 17612 32910 17668
rect 35410 17612 35420 17668
rect 35476 17612 35868 17668
rect 35924 17612 35934 17668
rect 36082 17612 36092 17668
rect 36148 17612 40012 17668
rect 40068 17612 40078 17668
rect 19404 17556 19460 17612
rect 36092 17556 36148 17612
rect 19404 17500 22204 17556
rect 22260 17500 27020 17556
rect 27076 17500 27086 17556
rect 31714 17500 31724 17556
rect 31780 17500 32172 17556
rect 32228 17500 32238 17556
rect 34066 17500 34076 17556
rect 34132 17500 36148 17556
rect 12430 17388 12440 17444
rect 12496 17388 22428 17444
rect 22484 17388 22494 17444
rect 32274 17388 32284 17444
rect 32340 17388 33180 17444
rect 33236 17388 33246 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 28578 17164 28588 17220
rect 28644 17164 29372 17220
rect 29428 17164 29438 17220
rect 39778 17164 39788 17220
rect 39844 17164 41076 17220
rect 41132 17164 43820 17220
rect 43876 17164 43886 17220
rect 12786 17052 12796 17108
rect 12852 17052 14476 17108
rect 14532 17052 14542 17108
rect 19842 17052 19852 17108
rect 19908 17052 21532 17108
rect 21588 17052 21598 17108
rect 24490 17052 24500 17108
rect 24556 17052 25452 17108
rect 25508 17052 27244 17108
rect 27300 17052 27310 17108
rect 27906 17052 27916 17108
rect 27972 17052 28476 17108
rect 28532 17052 30156 17108
rect 30212 17052 31164 17108
rect 31220 17052 31230 17108
rect 34290 17052 34300 17108
rect 34356 17052 34804 17108
rect 34860 17052 35980 17108
rect 36036 17052 36046 17108
rect 41682 17052 41692 17108
rect 41748 17052 42924 17108
rect 42980 17052 42990 17108
rect 9090 16940 9100 16996
rect 9156 16940 10444 16996
rect 10500 16940 13244 16996
rect 13300 16940 13310 16996
rect 27455 16940 27465 16996
rect 27521 16940 28028 16996
rect 28084 16940 29820 16996
rect 29876 16940 31948 16996
rect 32004 16940 32014 16996
rect 42354 16940 42364 16996
rect 42420 16940 43148 16996
rect 43204 16940 43214 16996
rect 8754 16828 8764 16884
rect 8820 16828 12124 16884
rect 12180 16828 12908 16884
rect 12964 16828 13468 16884
rect 13524 16828 13534 16884
rect 17714 16828 17724 16884
rect 17780 16828 18956 16884
rect 19012 16828 19022 16884
rect 19170 16828 19180 16884
rect 19236 16828 19740 16884
rect 19796 16828 19806 16884
rect 23986 16828 23996 16884
rect 24052 16828 25340 16884
rect 25396 16828 25406 16884
rect 26002 16828 26012 16884
rect 26068 16828 26908 16884
rect 26964 16828 30492 16884
rect 30548 16828 30558 16884
rect 30818 16828 30828 16884
rect 30884 16828 31388 16884
rect 31444 16828 31454 16884
rect 31602 16828 31612 16884
rect 31668 16828 32060 16884
rect 32116 16828 34188 16884
rect 34244 16828 34254 16884
rect 34962 16828 34972 16884
rect 35028 16828 35644 16884
rect 35700 16828 39116 16884
rect 39172 16828 41692 16884
rect 41748 16828 42812 16884
rect 42868 16828 42878 16884
rect 24210 16716 24220 16772
rect 24276 16716 27692 16772
rect 27748 16716 27758 16772
rect 29698 16716 29708 16772
rect 29764 16716 31948 16772
rect 32004 16716 32014 16772
rect 26002 16604 26012 16660
rect 26068 16604 26236 16660
rect 26292 16604 26302 16660
rect 26898 16604 26908 16660
rect 26964 16604 27468 16660
rect 27524 16604 27534 16660
rect 31490 16604 31500 16660
rect 31556 16604 31836 16660
rect 31892 16604 31902 16660
rect 8876 16492 13580 16548
rect 13636 16492 13646 16548
rect 24658 16492 24668 16548
rect 24724 16492 27580 16548
rect 27636 16492 27804 16548
rect 27860 16492 27870 16548
rect 31910 16492 31948 16548
rect 32004 16492 32014 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 8876 16436 8932 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 8866 16380 8876 16436
rect 8932 16380 8942 16436
rect 23874 16268 23884 16324
rect 23940 16268 24892 16324
rect 24948 16268 29932 16324
rect 29988 16268 31052 16324
rect 31108 16268 32508 16324
rect 32564 16268 32574 16324
rect 43530 16268 43540 16324
rect 43596 16268 44380 16324
rect 44436 16268 44446 16324
rect 45200 16212 46000 16240
rect 23090 16156 23100 16212
rect 23156 16156 23660 16212
rect 23716 16156 23726 16212
rect 27458 16156 27468 16212
rect 27524 16156 29596 16212
rect 29652 16156 29662 16212
rect 38434 16156 38444 16212
rect 38500 16156 39340 16212
rect 39396 16156 39900 16212
rect 39956 16156 40292 16212
rect 40348 16156 40358 16212
rect 44202 16156 44212 16212
rect 44268 16156 46000 16212
rect 45200 16128 46000 16156
rect 14334 16044 14344 16100
rect 14400 16044 18060 16100
rect 18116 16044 18126 16100
rect 22866 16044 22876 16100
rect 22932 16044 23324 16100
rect 23380 16044 23390 16100
rect 26786 16044 26796 16100
rect 26852 16044 26908 16100
rect 26964 16044 26974 16100
rect 27794 16044 27804 16100
rect 27860 16044 28364 16100
rect 28420 16044 29148 16100
rect 29204 16044 29214 16100
rect 29474 15932 29484 15988
rect 29540 15932 30604 15988
rect 30660 15932 30670 15988
rect 34514 15932 34524 15988
rect 34580 15932 39116 15988
rect 39172 15932 41468 15988
rect 41524 15932 41534 15988
rect 8978 15820 8988 15876
rect 9044 15820 10220 15876
rect 10276 15820 10286 15876
rect 10546 15820 10556 15876
rect 10612 15820 13468 15876
rect 13524 15820 13534 15876
rect 26114 15820 26124 15876
rect 26180 15820 28028 15876
rect 28084 15820 28094 15876
rect 35298 15820 35308 15876
rect 35364 15820 36540 15876
rect 36596 15820 36606 15876
rect 10556 15764 10612 15820
rect 7970 15708 7980 15764
rect 8036 15708 10612 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 12542 15596 12552 15652
rect 12608 15596 15148 15652
rect 15092 15540 15148 15596
rect 11554 15484 11564 15540
rect 11620 15484 12012 15540
rect 12068 15484 12684 15540
rect 12740 15484 12750 15540
rect 15092 15484 18228 15540
rect 18284 15484 18732 15540
rect 18788 15484 18798 15540
rect 23762 15484 23772 15540
rect 23828 15484 24276 15540
rect 24332 15484 25900 15540
rect 25956 15484 25966 15540
rect 28130 15484 28140 15540
rect 28196 15484 29036 15540
rect 29092 15484 36372 15540
rect 36428 15484 36438 15540
rect 43362 15484 43372 15540
rect 43428 15484 43652 15540
rect 43708 15484 43718 15540
rect 19506 15372 19516 15428
rect 19572 15372 19582 15428
rect 27458 15372 27468 15428
rect 27524 15372 29820 15428
rect 29876 15372 29886 15428
rect 30482 15372 30492 15428
rect 30548 15372 32004 15428
rect 32060 15372 32396 15428
rect 32452 15372 32462 15428
rect 19516 15316 19572 15372
rect 14802 15260 14812 15316
rect 14868 15260 16492 15316
rect 16548 15260 18396 15316
rect 18452 15260 19852 15316
rect 19908 15260 19918 15316
rect 21746 15260 21756 15316
rect 21812 15260 25788 15316
rect 25844 15260 26124 15316
rect 26180 15260 26190 15316
rect 28690 15260 28700 15316
rect 28756 15260 31052 15316
rect 31108 15260 31118 15316
rect 31490 15260 31500 15316
rect 31556 15260 32956 15316
rect 33012 15260 33022 15316
rect 36754 15260 36764 15316
rect 36820 15260 37212 15316
rect 37268 15260 40796 15316
rect 40852 15260 40862 15316
rect 8082 15148 8092 15204
rect 8148 15148 9100 15204
rect 9156 15148 11452 15204
rect 11508 15148 11518 15204
rect 18050 15148 18060 15204
rect 18116 15148 18844 15204
rect 18900 15148 18910 15204
rect 19282 15148 19292 15204
rect 19348 15148 19358 15204
rect 23090 15148 23100 15204
rect 23156 15148 24444 15204
rect 24500 15148 26012 15204
rect 26068 15148 26078 15204
rect 27570 15148 27580 15204
rect 27636 15148 31388 15204
rect 31444 15148 31454 15204
rect 36362 15148 36372 15204
rect 36428 15148 37660 15204
rect 37716 15148 37726 15204
rect 41580 15148 43036 15204
rect 43092 15148 43102 15204
rect 19292 15092 19348 15148
rect 41580 15092 41636 15148
rect 16146 15036 16156 15092
rect 16212 15036 18172 15092
rect 18228 15036 19348 15092
rect 30604 15036 30828 15092
rect 30884 15036 30894 15092
rect 35522 15036 35532 15092
rect 35588 15036 36876 15092
rect 36932 15036 36942 15092
rect 41570 15036 41580 15092
rect 41636 15036 41646 15092
rect 42372 15036 42382 15092
rect 42438 15036 43372 15092
rect 43428 15036 43438 15092
rect 30604 14980 30660 15036
rect 13682 14924 13692 14980
rect 13748 14924 14588 14980
rect 14644 14924 14654 14980
rect 18946 14924 18956 14980
rect 19012 14924 19516 14980
rect 19572 14924 22988 14980
rect 23044 14924 23054 14980
rect 28102 14924 28140 14980
rect 28196 14924 28206 14980
rect 30594 14924 30604 14980
rect 30660 14924 30670 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 13458 14812 13468 14868
rect 13524 14812 13534 14868
rect 42130 14812 42140 14868
rect 42196 14812 43596 14868
rect 43652 14812 43662 14868
rect 7522 14700 7532 14756
rect 7588 14700 8428 14756
rect 8484 14700 8494 14756
rect 8754 14588 8764 14644
rect 8820 14588 11564 14644
rect 11620 14588 11630 14644
rect 13468 14532 13524 14812
rect 37090 14700 37100 14756
rect 37156 14700 37772 14756
rect 37828 14700 37838 14756
rect 37986 14700 37996 14756
rect 38052 14700 38780 14756
rect 38836 14700 38846 14756
rect 42140 14644 42196 14812
rect 15922 14588 15932 14644
rect 15988 14588 21196 14644
rect 21252 14588 21420 14644
rect 21476 14588 21486 14644
rect 28914 14588 28924 14644
rect 28980 14588 29484 14644
rect 29540 14588 31332 14644
rect 31388 14588 42196 14644
rect 13458 14476 13468 14532
rect 13524 14476 13534 14532
rect 15586 14476 15596 14532
rect 15652 14476 16044 14532
rect 16100 14476 16110 14532
rect 26450 14476 26460 14532
rect 26516 14476 27244 14532
rect 27300 14476 28588 14532
rect 28644 14476 28654 14532
rect 35186 14476 35196 14532
rect 35252 14476 35980 14532
rect 36036 14476 36372 14532
rect 36428 14476 36438 14532
rect 7746 14364 7756 14420
rect 7812 14364 12124 14420
rect 12180 14364 12190 14420
rect 14334 14364 14344 14420
rect 14400 14364 19628 14420
rect 19684 14364 20020 14420
rect 20076 14364 20086 14420
rect 30594 14364 30604 14420
rect 30660 14364 31164 14420
rect 31220 14364 31230 14420
rect 35858 14364 35868 14420
rect 35924 14364 36988 14420
rect 37044 14364 37054 14420
rect 37892 14364 37902 14420
rect 37958 14364 39116 14420
rect 39172 14364 39182 14420
rect 15698 14252 15708 14308
rect 15764 14252 17164 14308
rect 17220 14252 17230 14308
rect 20290 14252 20300 14308
rect 20356 14252 22652 14308
rect 22708 14252 22718 14308
rect 26506 14252 26516 14308
rect 26572 14252 28140 14308
rect 28196 14252 28206 14308
rect 35690 14252 35700 14308
rect 35756 14252 35980 14308
rect 36036 14252 36046 14308
rect 42130 14252 42140 14308
rect 42196 14252 44100 14308
rect 44156 14252 44166 14308
rect 41626 14140 41636 14196
rect 41692 14140 43484 14196
rect 43540 14140 43550 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 8418 13916 8428 13972
rect 8484 13916 9716 13972
rect 21298 13916 21308 13972
rect 21364 13916 23100 13972
rect 23156 13916 24948 13972
rect 25004 13916 25014 13972
rect 36082 13916 36092 13972
rect 36148 13916 37324 13972
rect 37380 13916 37390 13972
rect 37650 13916 37660 13972
rect 37716 13916 41188 13972
rect 41244 13916 43148 13972
rect 43204 13916 43214 13972
rect 9660 13860 9716 13916
rect 7634 13804 7644 13860
rect 7700 13804 8540 13860
rect 8596 13804 8606 13860
rect 9650 13804 9660 13860
rect 9716 13804 13132 13860
rect 13188 13804 13198 13860
rect 41458 13804 41468 13860
rect 41524 13804 43484 13860
rect 43540 13804 43550 13860
rect 8082 13692 8092 13748
rect 8148 13692 8652 13748
rect 8708 13692 11340 13748
rect 11396 13692 11406 13748
rect 13234 13692 13244 13748
rect 13300 13692 13804 13748
rect 13860 13692 13870 13748
rect 16034 13692 16044 13748
rect 16100 13692 17052 13748
rect 17108 13692 17276 13748
rect 17332 13692 17342 13748
rect 21858 13692 21868 13748
rect 21924 13692 23996 13748
rect 24052 13692 26908 13748
rect 26964 13692 27692 13748
rect 27748 13692 27758 13748
rect 40450 13692 40460 13748
rect 40516 13692 42906 13748
rect 42962 13692 42972 13748
rect 8530 13580 8540 13636
rect 8596 13580 11676 13636
rect 11732 13580 11742 13636
rect 23202 13580 23212 13636
rect 23268 13580 24444 13636
rect 24500 13580 24510 13636
rect 35970 13580 35980 13636
rect 36036 13580 38780 13636
rect 38836 13580 38846 13636
rect 13468 13468 16660 13524
rect 16716 13468 16726 13524
rect 30594 13468 30604 13524
rect 30660 13468 31724 13524
rect 31780 13468 31790 13524
rect 32946 13468 32956 13524
rect 33012 13468 33292 13524
rect 33348 13468 34076 13524
rect 34132 13468 35868 13524
rect 35924 13468 35934 13524
rect 41794 13468 41804 13524
rect 41860 13468 43484 13524
rect 43540 13468 43550 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 13468 13300 13524 13468
rect 14476 13412 14532 13468
rect 14466 13356 14476 13412
rect 14532 13356 14542 13412
rect 31042 13356 31052 13412
rect 31108 13356 33628 13412
rect 33684 13356 33694 13412
rect 43250 13356 43260 13412
rect 43316 13356 43652 13412
rect 43708 13356 43718 13412
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 13458 13244 13468 13300
rect 13524 13244 13534 13300
rect 30930 13244 30940 13300
rect 30996 13244 31724 13300
rect 31780 13244 31790 13300
rect 28466 13132 28476 13188
rect 28532 13132 29372 13188
rect 29428 13132 29438 13188
rect 30594 13132 30604 13188
rect 30660 13132 31556 13188
rect 31500 13076 31556 13132
rect 8082 13020 8092 13076
rect 8148 13020 8988 13076
rect 9044 13020 9054 13076
rect 31490 13020 31500 13076
rect 31556 13020 36092 13076
rect 36148 13020 36158 13076
rect 40114 13020 40124 13076
rect 40180 13020 41356 13076
rect 41412 13020 41422 13076
rect 7354 12908 7364 12964
rect 7420 12908 9436 12964
rect 9492 12908 9502 12964
rect 32274 12908 32284 12964
rect 32340 12908 33460 12964
rect 33516 12908 33526 12964
rect 34346 12908 34356 12964
rect 34412 12908 35420 12964
rect 35476 12908 35486 12964
rect 35746 12908 35756 12964
rect 35812 12908 35980 12964
rect 36036 12908 36046 12964
rect 39778 12908 39788 12964
rect 39844 12908 40572 12964
rect 40628 12908 40638 12964
rect 45200 12852 46000 12880
rect 27346 12796 27356 12852
rect 27412 12796 33740 12852
rect 33796 12796 33806 12852
rect 37090 12796 37100 12852
rect 37156 12796 38892 12852
rect 38948 12796 38958 12852
rect 44370 12796 44380 12852
rect 44436 12796 46000 12852
rect 45200 12768 46000 12796
rect 25330 12684 25340 12740
rect 25396 12684 28252 12740
rect 28308 12684 28318 12740
rect 29698 12684 29708 12740
rect 29764 12684 31164 12740
rect 31220 12684 33068 12740
rect 33124 12684 33134 12740
rect 34962 12684 34972 12740
rect 35028 12684 36148 12740
rect 36204 12684 36214 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 35092 12460 35102 12516
rect 35158 12460 36092 12516
rect 36148 12460 36158 12516
rect 20738 12348 20748 12404
rect 20804 12348 28868 12404
rect 28924 12348 28934 12404
rect 33842 12348 33852 12404
rect 33908 12348 36428 12404
rect 36484 12348 36494 12404
rect 25218 12236 25228 12292
rect 25284 12236 26572 12292
rect 26628 12236 26638 12292
rect 35410 12236 35420 12292
rect 35476 12236 35644 12292
rect 35700 12236 35710 12292
rect 8194 12124 8204 12180
rect 8260 12124 10220 12180
rect 10276 12124 10286 12180
rect 16146 12124 16156 12180
rect 16212 12124 17612 12180
rect 17668 12124 17678 12180
rect 31826 12124 31836 12180
rect 31892 12124 35084 12180
rect 35140 12124 37324 12180
rect 37380 12124 37390 12180
rect 37762 12124 37772 12180
rect 37828 12124 40908 12180
rect 40964 12124 40974 12180
rect 41682 12124 41692 12180
rect 41748 12124 43932 12180
rect 43988 12124 43998 12180
rect 27234 12012 27244 12068
rect 27300 12012 33964 12068
rect 34020 12012 34030 12068
rect 24770 11900 24780 11956
rect 24836 11900 26142 11956
rect 26198 11900 26208 11956
rect 23650 11788 23660 11844
rect 23716 11788 24556 11844
rect 24612 11788 25396 11844
rect 25452 11788 25462 11844
rect 41701 11788 41711 11844
rect 41767 11788 43260 11844
rect 43316 11788 43326 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 26002 11676 26012 11732
rect 26068 11676 27020 11732
rect 27076 11676 27086 11732
rect 18610 11564 18620 11620
rect 18676 11564 19852 11620
rect 19908 11564 22316 11620
rect 22372 11564 22382 11620
rect 25330 11564 25340 11620
rect 25396 11564 26740 11620
rect 26796 11564 26806 11620
rect 31714 11564 31724 11620
rect 31780 11564 43932 11620
rect 43988 11564 43998 11620
rect 18386 11452 18396 11508
rect 18452 11452 20636 11508
rect 20692 11452 22428 11508
rect 22484 11452 22494 11508
rect 34290 11452 34300 11508
rect 34356 11452 35868 11508
rect 35924 11452 35934 11508
rect 31714 11340 31724 11396
rect 31780 11340 32508 11396
rect 32564 11340 33068 11396
rect 33124 11340 33134 11396
rect 34850 11340 34860 11396
rect 34916 11340 35980 11396
rect 36036 11340 36046 11396
rect 36194 11340 36204 11396
rect 36260 11340 36298 11396
rect 43530 11340 43540 11396
rect 43596 11340 44268 11396
rect 44324 11340 44334 11396
rect 32274 11228 32284 11284
rect 32340 11228 37212 11284
rect 37268 11228 39788 11284
rect 39844 11228 39854 11284
rect 41430 11228 41468 11284
rect 41524 11228 41534 11284
rect 14018 11116 14028 11172
rect 14084 11116 17108 11172
rect 17164 11116 18060 11172
rect 18116 11116 18126 11172
rect 32386 11116 32396 11172
rect 32452 11116 33944 11172
rect 34000 11116 34010 11172
rect 42970 11116 42980 11172
rect 43036 11116 44380 11172
rect 44436 11116 44446 11172
rect 29810 11004 29820 11060
rect 29876 11004 32508 11060
rect 32564 11004 32574 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 22642 10780 22652 10836
rect 22708 10780 24444 10836
rect 24500 10780 24510 10836
rect 36614 10780 36652 10836
rect 36708 10780 36718 10836
rect 32610 10668 32620 10724
rect 32676 10668 34412 10724
rect 34468 10668 34636 10724
rect 34692 10668 34702 10724
rect 39442 10668 39452 10724
rect 39508 10668 40012 10724
rect 40068 10668 41020 10724
rect 41076 10668 41086 10724
rect 16706 10556 16716 10612
rect 16772 10556 17836 10612
rect 17892 10556 17902 10612
rect 34178 10556 34188 10612
rect 34244 10556 38780 10612
rect 38836 10556 38846 10612
rect 39666 10556 39676 10612
rect 39732 10556 41244 10612
rect 41300 10556 41310 10612
rect 43894 10556 43932 10612
rect 43988 10556 43998 10612
rect 14802 10444 14812 10500
rect 14868 10444 17388 10500
rect 17444 10444 17454 10500
rect 27234 10444 27244 10500
rect 27300 10444 28476 10500
rect 28532 10444 28542 10500
rect 35606 10444 35644 10500
rect 35700 10444 35710 10500
rect 32610 10332 32620 10388
rect 32676 10332 35084 10388
rect 35140 10332 35150 10388
rect 24546 10220 24556 10276
rect 24612 10220 24622 10276
rect 26002 10220 26012 10276
rect 26068 10220 27112 10276
rect 27168 10220 27178 10276
rect 36316 10220 39340 10276
rect 39396 10220 39406 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 17938 9996 17948 10052
rect 18004 9996 18732 10052
rect 18788 9996 22316 10052
rect 22372 9996 22382 10052
rect 24556 9940 24612 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 24770 10108 24780 10164
rect 24836 10108 24846 10164
rect 30258 10108 30268 10164
rect 30324 10108 31612 10164
rect 31668 10108 31678 10164
rect 24780 10052 24836 10108
rect 36316 10052 36372 10220
rect 43810 10108 43820 10164
rect 43876 10108 43932 10164
rect 43988 10108 43998 10164
rect 24780 9996 25452 10052
rect 25508 9996 25518 10052
rect 35196 9996 36092 10052
rect 36148 9996 36158 10052
rect 36306 9996 36316 10052
rect 36372 9996 36382 10052
rect 36530 9996 36540 10052
rect 36596 9996 36652 10052
rect 36708 9996 36718 10052
rect 19730 9884 19740 9940
rect 19796 9884 21644 9940
rect 21700 9884 21710 9940
rect 23426 9884 23436 9940
rect 23492 9884 24612 9940
rect 35196 9828 35252 9996
rect 18610 9772 18620 9828
rect 18676 9772 21308 9828
rect 21364 9772 21374 9828
rect 35186 9772 35196 9828
rect 35252 9772 35262 9828
rect 39890 9772 39900 9828
rect 39956 9772 40180 9828
rect 40236 9772 40246 9828
rect 19282 9660 19292 9716
rect 19348 9660 24108 9716
rect 24164 9660 24174 9716
rect 30594 9660 30604 9716
rect 30660 9660 39452 9716
rect 39508 9660 39518 9716
rect 40450 9660 40460 9716
rect 40516 9660 42588 9716
rect 42644 9660 42924 9716
rect 42980 9660 42990 9716
rect 16930 9548 16940 9604
rect 16996 9548 17836 9604
rect 17892 9548 26236 9604
rect 26292 9548 26302 9604
rect 38612 9548 43932 9604
rect 43988 9548 43998 9604
rect 35522 9436 35532 9492
rect 35588 9436 35644 9492
rect 35700 9436 35710 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 38612 9380 38668 9548
rect 45200 9492 46000 9520
rect 44258 9436 44268 9492
rect 44324 9436 46000 9492
rect 45200 9408 46000 9436
rect 32162 9324 32172 9380
rect 32228 9324 38668 9380
rect 18946 9212 18956 9268
rect 19012 9212 23324 9268
rect 23380 9212 23390 9268
rect 35858 9212 35868 9268
rect 35924 9212 37996 9268
rect 38052 9212 40348 9268
rect 40404 9212 40414 9268
rect 17938 9100 17948 9156
rect 18004 9100 19292 9156
rect 19348 9100 19796 9156
rect 16314 8988 16324 9044
rect 16380 8988 18844 9044
rect 18900 8988 18910 9044
rect 19740 8932 19796 9100
rect 30930 8988 30940 9044
rect 30996 8988 31948 9044
rect 32004 8988 32014 9044
rect 37314 8988 37324 9044
rect 37380 8988 39452 9044
rect 39508 8988 39518 9044
rect 43082 8988 43092 9044
rect 43148 8988 43708 9044
rect 43764 8988 43774 9044
rect 16482 8876 16492 8932
rect 16548 8876 18620 8932
rect 18676 8876 18686 8932
rect 19730 8876 19740 8932
rect 19796 8876 19806 8932
rect 29138 8876 29148 8932
rect 29204 8876 29708 8932
rect 29764 8876 32956 8932
rect 33012 8876 33022 8932
rect 36166 8876 36204 8932
rect 36260 8876 36270 8932
rect 41010 8876 41020 8932
rect 41076 8876 43820 8932
rect 43876 8876 43886 8932
rect 17770 8764 17780 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 17836 8372 17892 8820
rect 34066 8764 34076 8820
rect 34132 8764 36652 8820
rect 36708 8764 36718 8820
rect 18610 8652 18620 8708
rect 18676 8652 19180 8708
rect 19236 8652 19246 8708
rect 20066 8652 20076 8708
rect 20132 8652 21196 8708
rect 21252 8652 21262 8708
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 24332 8540 25564 8596
rect 25620 8540 25630 8596
rect 24332 8484 24388 8540
rect 24220 8428 24388 8484
rect 24770 8428 24780 8484
rect 24836 8428 25228 8484
rect 25284 8428 25294 8484
rect 39890 8428 39900 8484
rect 39956 8428 40684 8484
rect 40740 8428 40750 8484
rect 17836 8316 19068 8372
rect 19124 8316 19134 8372
rect 24220 8260 24276 8428
rect 25666 8316 25676 8372
rect 25732 8316 26684 8372
rect 26740 8316 26750 8372
rect 29810 8316 29820 8372
rect 29876 8316 31164 8372
rect 31220 8316 31230 8372
rect 36530 8316 36540 8372
rect 36596 8316 37212 8372
rect 37268 8316 37884 8372
rect 37940 8316 37950 8372
rect 18844 8204 21532 8260
rect 21588 8204 23996 8260
rect 24052 8204 24062 8260
rect 24210 8204 24220 8260
rect 24276 8204 24286 8260
rect 24974 8204 24984 8260
rect 25040 8204 29260 8260
rect 29316 8204 29932 8260
rect 29988 8204 29998 8260
rect 32274 8204 32284 8260
rect 32340 8204 37548 8260
rect 37604 8204 37614 8260
rect 39218 8204 39228 8260
rect 39284 8204 39788 8260
rect 39844 8204 40908 8260
rect 40964 8204 40974 8260
rect 18844 7924 18900 8204
rect 23314 8092 23324 8148
rect 23380 8092 25770 8148
rect 25826 8092 25836 8148
rect 26002 8092 26012 8148
rect 26068 8092 27188 8148
rect 27244 8092 27254 8148
rect 28802 8092 28812 8148
rect 28868 8092 31948 8148
rect 32004 8092 32014 8148
rect 34402 8092 34412 8148
rect 34468 8092 39004 8148
rect 39060 8092 39070 8148
rect 26674 7980 26684 8036
rect 26740 7980 27636 8036
rect 27692 7980 28644 8036
rect 28700 7980 28710 8036
rect 36082 7980 36092 8036
rect 36148 7980 37212 8036
rect 37268 7980 41692 8036
rect 41748 7980 41758 8036
rect 18834 7868 18844 7924
rect 18900 7868 18910 7924
rect 25890 7868 25900 7924
rect 25956 7868 27020 7924
rect 27076 7868 27086 7924
rect 27178 7868 27188 7924
rect 27244 7868 30156 7924
rect 30212 7868 30222 7924
rect 37986 7868 37996 7924
rect 38052 7868 39564 7924
rect 39620 7868 39630 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 36978 7756 36988 7812
rect 37044 7756 41468 7812
rect 41524 7756 41534 7812
rect 37090 7644 37100 7700
rect 37156 7644 37324 7700
rect 37380 7644 37390 7700
rect 37548 7644 37772 7700
rect 37828 7644 37838 7700
rect 37548 7588 37604 7644
rect 26226 7532 26236 7588
rect 26292 7532 26908 7588
rect 29474 7532 29484 7588
rect 29540 7532 30044 7588
rect 30100 7532 31052 7588
rect 31108 7532 31118 7588
rect 36866 7532 36876 7588
rect 36932 7532 37604 7588
rect 37986 7532 37996 7588
rect 38052 7532 42812 7588
rect 42868 7532 42878 7588
rect 26852 7476 26908 7532
rect 16930 7420 16940 7476
rect 16996 7420 17724 7476
rect 17780 7420 17790 7476
rect 22306 7420 22316 7476
rect 22372 7420 22382 7476
rect 26852 7420 29372 7476
rect 29428 7420 34188 7476
rect 34244 7420 34254 7476
rect 35746 7420 35756 7476
rect 35812 7420 42252 7476
rect 42308 7420 43820 7476
rect 43876 7420 43886 7476
rect 22316 7364 22372 7420
rect 18946 7308 18956 7364
rect 19012 7308 21756 7364
rect 21812 7308 22372 7364
rect 37874 7308 37884 7364
rect 37940 7308 38444 7364
rect 38500 7308 38510 7364
rect 42914 7308 42924 7364
rect 42980 7308 43708 7364
rect 43764 7308 43774 7364
rect 37650 7196 37660 7252
rect 37716 7196 40124 7252
rect 40180 7196 40190 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 25890 6972 25900 7028
rect 25956 6972 26908 7028
rect 26964 6972 26974 7028
rect 27234 6972 27244 7028
rect 27300 6972 28364 7028
rect 28420 6972 28430 7028
rect 18498 6860 18508 6916
rect 18564 6860 22316 6916
rect 22372 6860 22382 6916
rect 37538 6860 37548 6916
rect 37604 6860 38892 6916
rect 38948 6860 38958 6916
rect 18610 6748 18620 6804
rect 18676 6748 22092 6804
rect 22148 6748 22158 6804
rect 28242 6748 28252 6804
rect 28308 6748 28644 6804
rect 28700 6748 28710 6804
rect 37314 6748 37324 6804
rect 37380 6748 37390 6804
rect 37324 6692 37380 6748
rect 19058 6636 19068 6692
rect 19124 6636 19134 6692
rect 20626 6636 20636 6692
rect 20692 6636 24444 6692
rect 24500 6636 24510 6692
rect 28110 6636 28120 6692
rect 28176 6636 29372 6692
rect 29428 6636 29652 6692
rect 29708 6636 29718 6692
rect 35410 6636 35420 6692
rect 35476 6636 36988 6692
rect 37044 6636 37054 6692
rect 37324 6636 39228 6692
rect 39284 6636 39294 6692
rect 19068 6468 19124 6636
rect 20382 6524 20392 6580
rect 20448 6524 23660 6580
rect 23716 6524 23726 6580
rect 24098 6524 24108 6580
rect 24164 6524 25788 6580
rect 25844 6524 25854 6580
rect 35634 6524 35644 6580
rect 35700 6524 37660 6580
rect 37716 6524 37726 6580
rect 41346 6524 41356 6580
rect 41412 6524 43036 6580
rect 43092 6524 43102 6580
rect 19068 6412 20244 6468
rect 24434 6412 24444 6468
rect 24500 6412 26031 6468
rect 26087 6412 26097 6468
rect 30146 6412 30156 6468
rect 30212 6412 31668 6468
rect 31724 6412 35756 6468
rect 35812 6412 35822 6468
rect 40114 6412 40124 6468
rect 40180 6412 43148 6468
rect 43204 6412 43214 6468
rect 20188 6356 20244 6412
rect 20188 6300 27244 6356
rect 27300 6300 27310 6356
rect 33740 6300 34748 6356
rect 34804 6300 34814 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 18610 6188 18620 6244
rect 18676 6188 19292 6244
rect 19348 6188 19358 6244
rect 33740 6132 33796 6300
rect 35242 6188 35252 6244
rect 35308 6188 39564 6244
rect 39620 6188 39630 6244
rect 45200 6132 46000 6160
rect 17714 6076 17724 6132
rect 17780 6076 18396 6132
rect 18452 6076 27692 6132
rect 27748 6076 27758 6132
rect 32162 6076 32172 6132
rect 32228 6076 33740 6132
rect 33796 6076 33806 6132
rect 36530 6076 36540 6132
rect 36596 6076 39676 6132
rect 39732 6076 40908 6132
rect 40964 6076 40974 6132
rect 44258 6076 44268 6132
rect 44324 6076 46000 6132
rect 45200 6048 46000 6076
rect 16930 5964 16940 6020
rect 16996 5964 17612 6020
rect 17668 5964 20636 6020
rect 20692 5964 25340 6020
rect 25396 5964 25406 6020
rect 35522 5964 35532 6020
rect 35588 5964 41692 6020
rect 41748 5964 41758 6020
rect 15138 5852 15148 5908
rect 15204 5852 16492 5908
rect 16548 5852 17836 5908
rect 17892 5852 19516 5908
rect 19572 5852 19582 5908
rect 22306 5852 22316 5908
rect 22372 5852 23436 5908
rect 23492 5852 23502 5908
rect 24994 5852 25004 5908
rect 25060 5852 25452 5908
rect 25508 5852 26216 5908
rect 26272 5852 26282 5908
rect 28558 5852 28568 5908
rect 28624 5852 29596 5908
rect 29652 5852 29662 5908
rect 33898 5852 33908 5908
rect 33964 5852 35663 5908
rect 35719 5852 35729 5908
rect 38882 5852 38892 5908
rect 38948 5852 39340 5908
rect 39396 5852 41244 5908
rect 41300 5852 41310 5908
rect 16594 5740 16604 5796
rect 16660 5740 17388 5796
rect 17444 5740 17454 5796
rect 18610 5740 18620 5796
rect 18676 5740 20412 5796
rect 20468 5740 20478 5796
rect 38770 5740 38780 5796
rect 38836 5740 40236 5796
rect 40292 5740 42700 5796
rect 42756 5740 42766 5796
rect 16762 5628 16772 5684
rect 16828 5628 17836 5684
rect 17892 5628 17902 5684
rect 34644 5628 34654 5684
rect 34710 5628 35924 5684
rect 35868 5572 35924 5628
rect 35858 5516 35868 5572
rect 35924 5516 35934 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 38546 5404 38556 5460
rect 38612 5404 44268 5460
rect 44324 5404 44334 5460
rect 31378 5292 31388 5348
rect 31444 5292 43932 5348
rect 43988 5292 43998 5348
rect 18274 5180 18284 5236
rect 18340 5180 22316 5236
rect 22372 5180 22382 5236
rect 25788 5180 27468 5236
rect 27524 5180 27534 5236
rect 38612 5180 39900 5236
rect 39956 5180 39966 5236
rect 21532 5124 21588 5180
rect 25788 5124 25844 5180
rect 38612 5124 38668 5180
rect 18050 5068 18060 5124
rect 18116 5068 18732 5124
rect 18788 5068 18798 5124
rect 21522 5068 21532 5124
rect 21588 5068 21598 5124
rect 21746 5068 21756 5124
rect 21812 5068 25788 5124
rect 25844 5068 25854 5124
rect 26786 5068 26796 5124
rect 26852 5068 28028 5124
rect 28084 5068 28094 5124
rect 33730 5068 33740 5124
rect 33796 5068 36316 5124
rect 36372 5068 36382 5124
rect 36642 5068 36652 5124
rect 36708 5068 37660 5124
rect 37716 5068 37726 5124
rect 38556 5068 38668 5124
rect 38770 5068 38780 5124
rect 38836 5068 40684 5124
rect 40740 5068 40750 5124
rect 17490 4956 17500 5012
rect 17556 4956 18284 5012
rect 18340 4956 20188 5012
rect 20244 4956 20254 5012
rect 21354 4844 21364 4900
rect 21420 4844 22204 4900
rect 22260 4844 22270 4900
rect 38490 4844 38500 4900
rect 38556 4844 38612 5068
rect 40338 4956 40348 5012
rect 40404 4956 42140 5012
rect 42196 4956 42588 5012
rect 42644 4956 42654 5012
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 22866 4508 22876 4564
rect 22932 4508 27244 4564
rect 27300 4508 27310 4564
rect 34850 4508 34860 4564
rect 34916 4508 36092 4564
rect 36148 4508 37231 4564
rect 37287 4508 37297 4564
rect 24322 4396 24332 4452
rect 24388 4396 28700 4452
rect 28756 4396 28766 4452
rect 17938 4284 17948 4340
rect 18004 4284 22540 4340
rect 22596 4284 22606 4340
rect 29026 4284 29036 4340
rect 29092 4284 30268 4340
rect 30324 4284 33628 4340
rect 33684 4284 33694 4340
rect 38518 4284 38556 4340
rect 38612 4284 38622 4340
rect 39106 4284 39116 4340
rect 39172 4284 40348 4340
rect 40404 4284 40414 4340
rect 21410 4172 21420 4228
rect 21476 4172 22428 4228
rect 22484 4172 22494 4228
rect 38322 4172 38332 4228
rect 38388 4172 41356 4228
rect 41412 4172 43932 4228
rect 43988 4172 43998 4228
rect 19506 4060 19516 4116
rect 19572 4060 22876 4116
rect 22932 4060 22942 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 22530 3724 22540 3780
rect 22596 3724 25564 3780
rect 25620 3724 25630 3780
rect 28354 3724 28364 3780
rect 28420 3724 29278 3780
rect 29334 3724 29344 3780
rect 17490 3500 17500 3556
rect 17556 3500 19516 3556
rect 19572 3500 19582 3556
rect 22978 3500 22988 3556
rect 23044 3500 24108 3556
rect 24164 3500 24556 3556
rect 24612 3500 24622 3556
rect 42130 3388 42140 3444
rect 42196 3388 42700 3444
rect 42756 3388 42766 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 45200 2772 46000 2800
rect 36866 2716 36876 2772
rect 36932 2716 46000 2772
rect 45200 2688 46000 2716
<< via3 >>
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 34412 37548 34468 37604
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 34524 37212 34580 37268
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 34524 36540 34580 36596
rect 34412 36204 34468 36260
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 24780 33740 24836 33796
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 24780 32956 24836 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 35644 32396 35700 32452
rect 30492 32284 30548 32340
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 35644 31724 35700 31780
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 30492 31052 30548 31108
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 36988 22988 37044 23044
rect 43596 22764 43652 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 36988 22316 37044 22372
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 16828 21532 16884 21588
rect 16828 21308 16884 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 31388 20524 31444 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 43372 19740 43428 19796
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 43596 18284 43652 18340
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 31948 16940 32004 16996
rect 31948 16492 32004 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 28140 15484 28196 15540
rect 43372 15484 43428 15540
rect 28140 14924 28196 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 36204 11340 36260 11396
rect 41468 11228 41524 11284
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 36652 10780 36708 10836
rect 43932 10556 43988 10612
rect 35644 10444 35700 10500
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 43932 10108 43988 10164
rect 36092 9996 36148 10052
rect 36652 9996 36708 10052
rect 35644 9436 35700 9492
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 36204 8876 36260 8932
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 41468 7756 41524 7812
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 38556 5404 38612 5460
rect 31388 5292 31444 5348
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 38556 4284 38612 4340
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 42396
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 42364 20128 42396
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 35168 41580 35488 42396
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 19808 36092 20128 37604
rect 34412 37604 34468 37614
rect 34412 36260 34468 37548
rect 34524 37268 34580 37278
rect 34524 36596 34580 37212
rect 34524 36530 34580 36540
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 34412 36194 34468 36204
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 24780 33796 24836 33806
rect 24780 33012 24836 33740
rect 24780 32946 24836 32956
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 30492 32340 30548 32350
rect 30492 31108 30548 32284
rect 30492 31042 30548 31052
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 16828 21588 16884 21598
rect 16828 21364 16884 21532
rect 16828 21298 16884 21308
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 20412 20128 21924
rect 35168 30604 35488 32116
rect 35644 32452 35700 32462
rect 35644 31780 35700 32396
rect 35644 31714 35700 31724
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 36988 23044 37044 23054
rect 36988 22372 37044 22988
rect 36988 22306 37044 22316
rect 43596 22820 43652 22830
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 31388 20580 31444 20590
rect 28140 15540 28196 15550
rect 28140 14980 28196 15484
rect 28140 14914 28196 14924
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 31388 5348 31444 20524
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 31948 16996 32004 17006
rect 31948 16548 32004 16940
rect 31948 16482 32004 16492
rect 35168 16492 35488 18004
rect 31388 5282 31444 5292
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 43372 19796 43428 19806
rect 43372 15540 43428 19740
rect 43596 18340 43652 22764
rect 43596 18274 43652 18284
rect 43372 15474 43428 15484
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 36204 11396 36260 11406
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35644 10500 35700 10510
rect 35644 9492 35700 10444
rect 36092 10052 36148 10062
rect 36204 10052 36260 11340
rect 41468 11284 41524 11294
rect 36148 9996 36260 10052
rect 36092 9986 36148 9996
rect 35644 9426 35700 9436
rect 36204 8932 36260 9996
rect 36652 10836 36708 10846
rect 36652 10052 36708 10780
rect 36652 9986 36708 9996
rect 36204 8866 36260 8876
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 41468 7812 41524 11228
rect 43932 10612 43988 10622
rect 43932 10164 43988 10556
rect 43932 10098 43988 10108
rect 41468 7746 41524 7756
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 3948 35488 5460
rect 38556 5460 38612 5470
rect 38556 4340 38612 5404
rect 38556 4274 38612 4284
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0529_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751534193
transform -1 0 22736 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0530_
timestamp 1751534193
transform -1 0 21840 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0531_
timestamp 1751534193
transform -1 0 19152 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0532_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751740063
transform 1 0 17696 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0533_
timestamp 1751740063
transform -1 0 12096 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0534_
timestamp 1751740063
transform 1 0 9968 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0535_
timestamp 1751740063
transform -1 0 12880 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0536_
timestamp 1751534193
transform -1 0 19824 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0537_
timestamp 1751740063
transform -1 0 16240 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0538_
timestamp 1751740063
transform -1 0 19264 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0539_
timestamp 1751740063
transform -1 0 16240 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0540_
timestamp 1751740063
transform -1 0 17472 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _0541_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751905124
transform -1 0 31248 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0542_
timestamp 1751534193
transform 1 0 31808 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0543_
timestamp 1751534193
transform -1 0 31024 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0544_
timestamp 1751534193
transform -1 0 32368 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0545_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752345181
transform -1 0 30352 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0546_
timestamp 1752345181
transform -1 0 31024 0 -1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0547_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889408
transform 1 0 30128 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0548_
timestamp 1752345181
transform -1 0 28112 0 1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0549_
timestamp 1752345181
transform -1 0 28672 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0550_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751531619
transform 1 0 29008 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _0551_
timestamp 1751905124
transform 1 0 20720 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0552_
timestamp 1751534193
transform 1 0 22288 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0553_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753277515
transform -1 0 43232 0 -1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0554_
timestamp 1753277515
transform -1 0 44016 0 1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0555_
timestamp 1753277515
transform 1 0 38416 0 -1 26656
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0556_
timestamp 1753277515
transform 1 0 33488 0 -1 26656
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0557_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753172561
transform -1 0 41552 0 1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0558_
timestamp 1753277515
transform 1 0 34720 0 -1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0559_
timestamp 1753277515
transform -1 0 39984 0 1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0560_
timestamp 1753277515
transform 1 0 38976 0 -1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0561_
timestamp 1752345181
transform 1 0 38416 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0562_
timestamp 1753277515
transform 1 0 36288 0 -1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0563_
timestamp 1753277515
transform 1 0 34944 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0564_
timestamp 1753277515
transform 1 0 36848 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0565_
timestamp 1753277515
transform -1 0 44240 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0566_
timestamp 1753172561
transform 1 0 37856 0 -1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0567_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753182340
transform -1 0 38416 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0568_
timestamp 1751534193
transform -1 0 31024 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0569_
timestamp 1751889408
transform 1 0 29120 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0570_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753960525
transform -1 0 30128 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0571_
timestamp 1753277515
transform 1 0 29792 0 -1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0572_
timestamp 1751534193
transform -1 0 36624 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0573_
timestamp 1751534193
transform 1 0 38528 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0574_
timestamp 1751740063
transform 1 0 40880 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0575_
timestamp 1751740063
transform -1 0 44016 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0576_
timestamp 1751740063
transform -1 0 44352 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0577_
timestamp 1751740063
transform 1 0 40768 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0578_
timestamp 1751534193
transform 1 0 32032 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0579_
timestamp 1751740063
transform -1 0 37632 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0580_
timestamp 1751740063
transform -1 0 34272 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0581_
timestamp 1751740063
transform -1 0 36624 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0582_
timestamp 1751740063
transform 1 0 32816 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0583_
timestamp 1751740063
transform 1 0 35280 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0584_
timestamp 1751740063
transform 1 0 36960 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0585_
timestamp 1751740063
transform 1 0 29008 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0586_
timestamp 1751534193
transform -1 0 27328 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0587_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform 1 0 27440 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0588_
timestamp 1751534193
transform -1 0 28784 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0589_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889808
transform -1 0 27552 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0590_
timestamp 1753277515
transform 1 0 23968 0 1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0591_
timestamp 1753277515
transform 1 0 22176 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0592_
timestamp 1753277515
transform 1 0 22624 0 -1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0593_
timestamp 1752345181
transform -1 0 25200 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0594_
timestamp 1753277515
transform -1 0 27104 0 1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0595_
timestamp 1753277515
transform 1 0 19376 0 1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0596_
timestamp 1753277515
transform 1 0 23296 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0597_
timestamp 1753277515
transform 1 0 23968 0 1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0598_
timestamp 1753172561
transform 1 0 23968 0 1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0599_
timestamp 1753277515
transform 1 0 25200 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0600_
timestamp 1753277515
transform 1 0 27104 0 1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0601_
timestamp 1753277515
transform 1 0 26096 0 1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0602_
timestamp 1753277515
transform 1 0 27552 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0603_
timestamp 1753172561
transform 1 0 26768 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0604_
timestamp 1753182340
transform 1 0 25088 0 -1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0605_
timestamp 1751534193
transform -1 0 25760 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0606_
timestamp 1751889408
transform -1 0 24416 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0607_
timestamp 1753960525
transform 1 0 24528 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0608_
timestamp 1753277515
transform -1 0 21280 0 -1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0609_
timestamp 1751534193
transform -1 0 19040 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0610_
timestamp 1751534193
transform 1 0 20272 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0611_
timestamp 1751740063
transform 1 0 17472 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0612_
timestamp 1751740063
transform -1 0 23072 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0613_
timestamp 1751740063
transform 1 0 18032 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0614_
timestamp 1751740063
transform 1 0 18816 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0615_
timestamp 1751534193
transform -1 0 20384 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0616_
timestamp 1751740063
transform 1 0 19488 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0617_
timestamp 1751740063
transform 1 0 18256 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0618_
timestamp 1751740063
transform -1 0 19040 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0619_
timestamp 1751740063
transform -1 0 18816 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0620_
timestamp 1751740063
transform -1 0 18032 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0621_
timestamp 1751740063
transform -1 0 18032 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0622_
timestamp 1753277515
transform 1 0 13328 0 1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0623_
timestamp 1753277515
transform 1 0 13440 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0624_
timestamp 1753277515
transform 1 0 13440 0 1 20384
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0625_
timestamp 1752345181
transform 1 0 14448 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0626_
timestamp 1753277515
transform 1 0 12432 0 -1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0627_
timestamp 1753277515
transform 1 0 13328 0 1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0628_
timestamp 1753277515
transform 1 0 13328 0 1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0629_
timestamp 1753277515
transform 1 0 12992 0 -1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0630_
timestamp 1753172561
transform 1 0 13104 0 -1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0631_
timestamp 1753277515
transform 1 0 11424 0 1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0632_
timestamp 1753277515
transform 1 0 11536 0 1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0633_
timestamp 1753277515
transform 1 0 12432 0 -1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0634_
timestamp 1753277515
transform 1 0 11536 0 1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0635_
timestamp 1753172561
transform 1 0 13328 0 1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0636_
timestamp 1753182340
transform 1 0 14896 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0637_
timestamp 1751534193
transform 1 0 17584 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0638_
timestamp 1751740063
transform 1 0 27552 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0639_
timestamp 1751531619
transform -1 0 27664 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0640_
timestamp 1751740063
transform -1 0 30576 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_4  _0641_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751882821
transform 1 0 25984 0 -1 18816
box -86 -86 1542 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0642_
timestamp 1751531619
transform -1 0 25088 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0643_
timestamp 1751889408
transform -1 0 26880 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0644_
timestamp 1751531619
transform -1 0 24304 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0645_
timestamp 1752345181
transform -1 0 22400 0 1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0646_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753868718
transform -1 0 21392 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0647_
timestamp 1753277515
transform -1 0 20944 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0648_
timestamp 1751534193
transform 1 0 8512 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0649_
timestamp 1751534193
transform -1 0 11536 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0650_
timestamp 1751740063
transform 1 0 8400 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0651_
timestamp 1751740063
transform 1 0 7616 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0652_
timestamp 1751740063
transform 1 0 8176 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0653_
timestamp 1751740063
transform 1 0 8400 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0654_
timestamp 1751534193
transform -1 0 14560 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0655_
timestamp 1751740063
transform -1 0 10752 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0656_
timestamp 1751740063
transform 1 0 9408 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0657_
timestamp 1751740063
transform -1 0 11088 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0658_
timestamp 1751740063
transform -1 0 12880 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0659_
timestamp 1751740063
transform -1 0 11536 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0660_
timestamp 1751740063
transform 1 0 7616 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0661_
timestamp 1753277515
transform -1 0 36736 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0662_
timestamp 1753277515
transform -1 0 38304 0 -1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0663_
timestamp 1753277515
transform 1 0 34496 0 1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0664_
timestamp 1752345181
transform 1 0 36848 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0665_
timestamp 1753277515
transform -1 0 42560 0 -1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0666_
timestamp 1753277515
transform 1 0 35056 0 1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0667_
timestamp 1753277515
transform -1 0 41216 0 1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0668_
timestamp 1753277515
transform 1 0 32928 0 -1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0669_
timestamp 1753172561
transform -1 0 39984 0 -1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0670_
timestamp 1753277515
transform -1 0 44128 0 -1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0671_
timestamp 1753277515
transform -1 0 39760 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0672_
timestamp 1753277515
transform -1 0 40544 0 -1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0673_
timestamp 1753277515
transform -1 0 42784 0 1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0674_
timestamp 1753172561
transform -1 0 38192 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0675_
timestamp 1753182340
transform 1 0 39312 0 -1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0676_
timestamp 1751534193
transform -1 0 30688 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0677_
timestamp 1751532043
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0678_
timestamp 1751889808
transform 1 0 29344 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0679_
timestamp 1751889808
transform 1 0 30016 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0680_
timestamp 1751534193
transform 1 0 32816 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0681_
timestamp 1751740063
transform 1 0 28672 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0682_
timestamp 1751531619
transform 1 0 30912 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0683_
timestamp 1751531619
transform 1 0 32032 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0684_
timestamp 1752345181
transform -1 0 32480 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0685_
timestamp 1753868718
transform 1 0 28560 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0686_
timestamp 1753277515
transform 1 0 29792 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0687_
timestamp 1751534193
transform 1 0 31920 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0688_
timestamp 1751534193
transform -1 0 35840 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0689_
timestamp 1751740063
transform 1 0 42896 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0690_
timestamp 1751740063
transform -1 0 44240 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0691_
timestamp 1751740063
transform -1 0 39424 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0692_
timestamp 1751740063
transform 1 0 40768 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0693_
timestamp 1751534193
transform -1 0 34496 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0694_
timestamp 1751740063
transform 1 0 34496 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0695_
timestamp 1751740063
transform -1 0 36512 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0696_
timestamp 1751740063
transform -1 0 36624 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0697_
timestamp 1751740063
transform -1 0 37632 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0698_
timestamp 1751740063
transform -1 0 40544 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0699_
timestamp 1751740063
transform -1 0 44352 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0700__1
timestamp 1751532043
transform -1 0 20944 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0701_
timestamp 1751532043
transform -1 0 20160 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0702_
timestamp 1751532043
transform -1 0 23184 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0703_
timestamp 1751532043
transform 1 0 29456 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0704_
timestamp 1751532043
transform -1 0 29120 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0705_
timestamp 1751532043
transform -1 0 25536 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0706_
timestamp 1751532043
transform 1 0 28112 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0707_
timestamp 1751532043
transform -1 0 29904 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0708_
timestamp 1751532043
transform -1 0 12544 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0709_
timestamp 1753277515
transform 1 0 9408 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0710_
timestamp 1753277515
transform -1 0 10976 0 -1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0711_
timestamp 1753277515
transform -1 0 12768 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0712_
timestamp 1751534193
transform -1 0 37520 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0713_
timestamp 1751534193
transform -1 0 32032 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0714_
timestamp 1751531619
transform 1 0 34048 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0715_
timestamp 1751531619
transform 1 0 33712 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0716_
timestamp 1751740063
transform -1 0 37184 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0717_
timestamp 1751534193
transform 1 0 37856 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0718_
timestamp 1751534193
transform 1 0 39200 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0719_
timestamp 1751534193
transform -1 0 35392 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0720_
timestamp 1751740063
transform 1 0 36848 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0721_
timestamp 1751889408
transform 1 0 38080 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0722_
timestamp 1753182340
transform 1 0 36848 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0723_
timestamp 1751534193
transform 1 0 37632 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0724_
timestamp 1751740063
transform -1 0 36624 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0725_
timestamp 1751889408
transform -1 0 37184 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0726_
timestamp 1753182340
transform -1 0 36624 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0727_
timestamp 1751534193
transform -1 0 35840 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0728_
timestamp 1753277515
transform -1 0 34496 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0729_
timestamp 1751740063
transform -1 0 31808 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0730_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753371985
transform 1 0 32032 0 -1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0731_
timestamp 1751740063
transform -1 0 33936 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0732_
timestamp 1751532043
transform -1 0 36624 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0733_
timestamp 1751740063
transform 1 0 35616 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0734_
timestamp 1751534193
transform 1 0 37184 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0735_
timestamp 1751534193
transform 1 0 39872 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0736_
timestamp 1753868718
transform 1 0 39312 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0737_
timestamp 1751534193
transform -1 0 40544 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0738_
timestamp 1753868718
transform -1 0 41552 0 1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0739_
timestamp 1751534193
transform -1 0 39872 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0740_
timestamp 1753868718
transform 1 0 39312 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0741_
timestamp 1751534193
transform 1 0 43344 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0742_
timestamp 1753868718
transform 1 0 41440 0 1 37632
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0743_
timestamp 1751534193
transform 1 0 42672 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0744_
timestamp 1751534193
transform -1 0 31920 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0745_
timestamp 1751534193
transform 1 0 34496 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0746_
timestamp 1751531619
transform -1 0 33712 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0747_
timestamp 1751889408
transform -1 0 32256 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0748_
timestamp 1753868718
transform -1 0 41552 0 1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0749_
timestamp 1751534193
transform -1 0 39872 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0750_
timestamp 1751889408
transform -1 0 34048 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0751_
timestamp 1751889408
transform 1 0 32928 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0752_
timestamp 1751534193
transform 1 0 35280 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0753_
timestamp 1751532043
transform 1 0 38640 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0754_
timestamp 1751534193
transform -1 0 39760 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0755_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751914308
transform 1 0 22064 0 -1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0756_
timestamp 1751534193
transform -1 0 20944 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0757_
timestamp 1751534193
transform 1 0 43680 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0758_
timestamp 1751914308
transform 1 0 21168 0 1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0759_
timestamp 1751534193
transform 1 0 22176 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0760_
timestamp 1751534193
transform 1 0 43008 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0761_
timestamp 1751914308
transform -1 0 22512 0 1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0762_
timestamp 1751534193
transform -1 0 20944 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0763_
timestamp 1751534193
transform -1 0 32256 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0764_
timestamp 1751534193
transform 1 0 24080 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0765_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752061876
transform -1 0 25872 0 1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0766_
timestamp 1751889408
transform 1 0 29008 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0767_
timestamp 1751534193
transform -1 0 31136 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0768_
timestamp 1751889808
transform -1 0 27552 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0769_
timestamp 1751531619
transform 1 0 25984 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0770_
timestamp 1751740063
transform -1 0 27104 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0771_
timestamp 1751889808
transform 1 0 28112 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0772_
timestamp 1752345181
transform 1 0 27104 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0773_
timestamp 1751889408
transform 1 0 24080 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0774_
timestamp 1751889408
transform -1 0 26320 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0775_
timestamp 1751534193
transform -1 0 24864 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0776_
timestamp 1751532043
transform 1 0 23744 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0777_
timestamp 1751740063
transform -1 0 23632 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _0778_
timestamp 1751905124
transform 1 0 22512 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0779_
timestamp 1753371985
transform -1 0 23856 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0780_
timestamp 1751889408
transform 1 0 23296 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0781_
timestamp 1751889808
transform -1 0 22848 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0782_
timestamp 1751531619
transform -1 0 22512 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0783_
timestamp 1751740063
transform -1 0 20944 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0784_
timestamp 1751889408
transform -1 0 23296 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0785_
timestamp 1751889808
transform 1 0 23408 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0786_
timestamp 1751531619
transform -1 0 22512 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0787_
timestamp 1751740063
transform -1 0 20944 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0788_
timestamp 1751531619
transform 1 0 21168 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0789_
timestamp 1751889808
transform 1 0 22624 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0790_
timestamp 1751889408
transform -1 0 22736 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0791_
timestamp 1751889408
transform 1 0 22736 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0792_
timestamp 1751534193
transform -1 0 21840 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0793_
timestamp 1753277515
transform 1 0 21168 0 1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0794_
timestamp 1751889408
transform -1 0 23184 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0795_
timestamp 1751534193
transform -1 0 20944 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0796_
timestamp 1751889808
transform -1 0 31808 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0797_
timestamp 1751889408
transform -1 0 31136 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0798_
timestamp 1751534193
transform -1 0 30352 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0799_
timestamp 1751531619
transform -1 0 34832 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0800_
timestamp 1751889808
transform -1 0 33712 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0801_
timestamp 1751889808
transform 1 0 31808 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0802_
timestamp 1751889408
transform 1 0 30800 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0803_
timestamp 1751889408
transform -1 0 32032 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0804_
timestamp 1751534193
transform 1 0 32032 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0805_
timestamp 1751534193
transform 1 0 25536 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0806_
timestamp 1751534193
transform 1 0 29232 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0807_
timestamp 1751534193
transform 1 0 26320 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0808_
timestamp 1753868718
transform -1 0 25760 0 1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0809_
timestamp 1753172561
transform -1 0 26656 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0810_
timestamp 1752061876
transform 1 0 32816 0 1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0811_
timestamp 1753960525
transform -1 0 35056 0 1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0812_
timestamp 1753960525
transform -1 0 27776 0 -1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0813_
timestamp 1751889408
transform 1 0 26096 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0814_
timestamp 1751534193
transform 1 0 29008 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0815_
timestamp 1751531619
transform 1 0 24080 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0816_
timestamp 1751889408
transform -1 0 24864 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0817_
timestamp 1753277515
transform 1 0 26432 0 1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0818_
timestamp 1753277515
transform 1 0 26768 0 1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0819_
timestamp 1753868718
transform -1 0 38080 0 -1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0820_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753441877
transform 1 0 35504 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0821_
timestamp 1751534193
transform 1 0 37968 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0822_
timestamp 1751531619
transform 1 0 28000 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _0823_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753272495
transform 1 0 29008 0 1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0824_
timestamp 1751889408
transform 1 0 24976 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0825_
timestamp 1751889408
transform 1 0 28448 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0826_
timestamp 1753277515
transform 1 0 30128 0 1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0827_
timestamp 1751531619
transform 1 0 31808 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0828_
timestamp 1751740063
transform 1 0 31024 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0829_
timestamp 1751532043
transform 1 0 33376 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0830_
timestamp 1753868718
transform -1 0 37520 0 -1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0831_
timestamp 1753960525
transform -1 0 35504 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0832_
timestamp 1751534193
transform 1 0 34832 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0833_
timestamp 1753172561
transform 1 0 26656 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0834_
timestamp 1753868718
transform 1 0 27104 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0835_
timestamp 1751889408
transform 1 0 30576 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0836_
timestamp 1753441877
transform 1 0 31584 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0837_
timestamp 1751531619
transform 1 0 34048 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0838_
timestamp 1751889808
transform 1 0 35504 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0839_
timestamp 1753868718
transform -1 0 38080 0 1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0840_
timestamp 1753960525
transform -1 0 34944 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0841_
timestamp 1751534193
transform 1 0 35504 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0842_
timestamp 1751532043
transform 1 0 30128 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0843_
timestamp 1753441877
transform 1 0 30464 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _0844_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753579406
transform -1 0 33264 0 1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0845_
timestamp 1751889408
transform 1 0 31360 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0846_
timestamp 1751889408
transform 1 0 28112 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0847_
timestamp 1753277515
transform 1 0 31472 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0848_
timestamp 1753868718
transform 1 0 31472 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0849_
timestamp 1751531619
transform 1 0 30576 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0850_
timestamp 1753277515
transform 1 0 31136 0 -1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0851_
timestamp 1753441877
transform 1 0 33040 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0852_
timestamp 1753441877
transform 1 0 33264 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0853_
timestamp 1751531619
transform -1 0 35280 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0854_
timestamp 1751889808
transform 1 0 34944 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0855_
timestamp 1751531619
transform 1 0 31920 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _0856_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753891287
transform -1 0 34496 0 -1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0857_
timestamp 1753441877
transform 1 0 32928 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0858_
timestamp 1753960525
transform 1 0 33824 0 -1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0859_
timestamp 1753868718
transform -1 0 40544 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0860_
timestamp 1751534193
transform 1 0 39872 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_4  _0861_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752051650
transform 1 0 27328 0 -1 17248
box -86 -86 1881 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0862_
timestamp 1751914308
transform -1 0 24864 0 -1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0863_
timestamp 1751534193
transform 1 0 25088 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0864_
timestamp 1751914308
transform -1 0 24864 0 -1 17248
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0865_
timestamp 1751534193
transform -1 0 23520 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0866_
timestamp 1751914308
transform -1 0 30352 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0867_
timestamp 1751534193
transform 1 0 29008 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0868_
timestamp 1751534193
transform -1 0 27552 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0869_
timestamp 1751914308
transform 1 0 27328 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0870_
timestamp 1751534193
transform 1 0 31024 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0871_
timestamp 1752061876
transform -1 0 28784 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0872_
timestamp 1751534193
transform -1 0 19040 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0873_
timestamp 1751889808
transform 1 0 16128 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0874_
timestamp 1751534193
transform -1 0 15232 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0875_
timestamp 1751534193
transform -1 0 19936 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0876_
timestamp 1751889408
transform 1 0 16240 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0877_
timestamp 1751534193
transform 1 0 18256 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0878_
timestamp 1751889808
transform 1 0 17024 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0879_
timestamp 1751534193
transform 1 0 17248 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0880_
timestamp 1751889408
transform -1 0 18032 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0881_
timestamp 1751534193
transform -1 0 15120 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0882_
timestamp 1751889808
transform -1 0 15904 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0883_
timestamp 1751534193
transform -1 0 14000 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0884_
timestamp 1751889408
transform 1 0 16240 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0885_
timestamp 1751534193
transform -1 0 16912 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0886_
timestamp 1751889808
transform -1 0 18032 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0887_
timestamp 1751534193
transform -1 0 16912 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0888_
timestamp 1751889808
transform 1 0 17584 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0889_
timestamp 1751534193
transform 1 0 18032 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0890_
timestamp 1751534193
transform 1 0 34160 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0891_
timestamp 1751914308
transform -1 0 39312 0 1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0892_
timestamp 1751534193
transform 1 0 38416 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0893_
timestamp 1751914308
transform 1 0 41328 0 -1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0894_
timestamp 1751534193
transform 1 0 42672 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0895_
timestamp 1751914308
transform 1 0 41328 0 -1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0896_
timestamp 1751534193
transform 1 0 43568 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0897_
timestamp 1751914308
transform -1 0 44016 0 -1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0898_
timestamp 1751534193
transform -1 0 40544 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0899_
timestamp 1751534193
transform 1 0 39760 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0900_
timestamp 1751534193
transform -1 0 34160 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0901_
timestamp 1751534193
transform 1 0 32928 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0902_
timestamp 1751914308
transform -1 0 33152 0 1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0903_
timestamp 1751534193
transform -1 0 32144 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0904_
timestamp 1751534193
transform -1 0 44352 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0905_
timestamp 1751534193
transform -1 0 35616 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0906_
timestamp 1751914308
transform 1 0 34048 0 1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0907_
timestamp 1751534193
transform 1 0 36064 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0908_
timestamp 1751534193
transform -1 0 43008 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0909_
timestamp 1751534193
transform 1 0 35616 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0910_
timestamp 1751914308
transform -1 0 36064 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0911_
timestamp 1751534193
transform 1 0 35168 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0912_
timestamp 1751914308
transform 1 0 36848 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0913_
timestamp 1751534193
transform 1 0 39088 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0914_
timestamp 1751532043
transform 1 0 42896 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0915_
timestamp 1751532043
transform 1 0 39984 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0916_
timestamp 1751532043
transform -1 0 37296 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0917_
timestamp 1751532043
transform -1 0 35840 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0918_
timestamp 1751532043
transform -1 0 32704 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0919_
timestamp 1751532043
transform -1 0 31696 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0920_
timestamp 1751740063
transform -1 0 32816 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0921_
timestamp 1751532043
transform 1 0 42672 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0922_
timestamp 1751532043
transform 1 0 38304 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0923_
timestamp 1751532043
transform 1 0 42784 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0924_
timestamp 1751532043
transform 1 0 43792 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0925_
timestamp 1751889408
transform -1 0 19712 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0926_
timestamp 1751534193
transform 1 0 19712 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0927_
timestamp 1751531619
transform 1 0 31248 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0928_
timestamp 1751914308
transform -1 0 34272 0 -1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0929_
timestamp 1751534193
transform -1 0 32480 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0930_
timestamp 1751914308
transform -1 0 35616 0 -1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0931_
timestamp 1751534193
transform -1 0 34272 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0932_
timestamp 1751914308
transform -1 0 35168 0 1 17248
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0933_
timestamp 1751534193
transform 1 0 34160 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0934_
timestamp 1751532043
transform -1 0 7616 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0935_
timestamp 1751532043
transform -1 0 8512 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0936_
timestamp 1751532043
transform -1 0 8624 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0937_
timestamp 1751532043
transform -1 0 10864 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0938_
timestamp 1751740063
transform -1 0 8960 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0939_
timestamp 1751532043
transform 1 0 8064 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0940_
timestamp 1751532043
transform -1 0 9968 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0941_
timestamp 1751532043
transform -1 0 9184 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0942_
timestamp 1751532043
transform -1 0 12992 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0943_
timestamp 1751532043
transform -1 0 7616 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0944_
timestamp 1751532043
transform 1 0 29008 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0945_
timestamp 1751532043
transform 1 0 25200 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0946_
timestamp 1751532043
transform 1 0 22960 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0947_
timestamp 1751532043
transform 1 0 7728 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0948_
timestamp 1751534193
transform -1 0 19488 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0949_
timestamp 1751914308
transform 1 0 15680 0 -1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0950_
timestamp 1751534193
transform 1 0 17248 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0951_
timestamp 1751914308
transform -1 0 19376 0 1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0952_
timestamp 1751534193
transform -1 0 16912 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0953_
timestamp 1751914308
transform -1 0 18592 0 -1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0954_
timestamp 1751534193
transform -1 0 17024 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0955_
timestamp 1751534193
transform -1 0 26432 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0956_
timestamp 1751914308
transform -1 0 18592 0 -1 17248
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0957_
timestamp 1751534193
transform -1 0 17024 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0958_
timestamp 1751534193
transform -1 0 19936 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0959_
timestamp 1751914308
transform 1 0 14672 0 -1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0960_
timestamp 1751534193
transform 1 0 17248 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0961_
timestamp 1751914308
transform -1 0 17024 0 -1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0962_
timestamp 1751534193
transform -1 0 15680 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0963_
timestamp 1751914308
transform -1 0 18592 0 -1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0964_
timestamp 1751534193
transform -1 0 17024 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0965_
timestamp 1751914308
transform -1 0 20384 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0966_
timestamp 1751534193
transform -1 0 19264 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0967_
timestamp 1751534193
transform -1 0 34272 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0968_
timestamp 1751914308
transform -1 0 34944 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0969_
timestamp 1751534193
transform 1 0 34272 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0970_
timestamp 1751534193
transform -1 0 35728 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0971_
timestamp 1751914308
transform 1 0 34944 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0972_
timestamp 1751534193
transform 1 0 36400 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0973_
timestamp 1751534193
transform -1 0 34944 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0974_
timestamp 1751914308
transform 1 0 33600 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0975_
timestamp 1751534193
transform 1 0 35952 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0976_
timestamp 1751532043
transform -1 0 17024 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0977_
timestamp 1751532043
transform -1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0978_
timestamp 1751532043
transform -1 0 17024 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0979_
timestamp 1751532043
transform -1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0980_
timestamp 1751740063
transform -1 0 18032 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0981_
timestamp 1751532043
transform -1 0 17024 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0982_
timestamp 1751532043
transform -1 0 22512 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0983_
timestamp 1751532043
transform -1 0 18032 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0984_
timestamp 1751532043
transform 1 0 18928 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0985_
timestamp 1751532043
transform -1 0 21616 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0986_
timestamp 1751532043
transform -1 0 17584 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_4  _0987_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751830969
transform -1 0 26544 0 1 17248
box -86 -86 1545 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0988_
timestamp 1751914308
transform 1 0 26544 0 1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0989_
timestamp 1751534193
transform 1 0 27776 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0990_
timestamp 1751914308
transform 1 0 25088 0 -1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0991_
timestamp 1751534193
transform -1 0 24864 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0992_
timestamp 1751914308
transform 1 0 26432 0 -1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0993_
timestamp 1751534193
transform 1 0 28112 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0994_
timestamp 1751914308
transform -1 0 25312 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0995_
timestamp 1751534193
transform 1 0 24080 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_4  _0996_
timestamp 1751830969
transform -1 0 26656 0 -1 17248
box -86 -86 1545 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0997_
timestamp 1751914308
transform 1 0 28224 0 1 3136
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0998_
timestamp 1751534193
transform -1 0 28448 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0999_
timestamp 1751914308
transform -1 0 26880 0 1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1000_
timestamp 1751534193
transform -1 0 23296 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1001_
timestamp 1751914308
transform 1 0 25424 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1002_
timestamp 1751534193
transform 1 0 26768 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1003_
timestamp 1751914308
transform -1 0 23968 0 -1 15680
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1004_
timestamp 1751534193
transform -1 0 22624 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1005_
timestamp 1751531619
transform 1 0 30352 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1006_
timestamp 1751914308
transform 1 0 29456 0 -1 4704
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1007_
timestamp 1751534193
transform 1 0 30240 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1008_
timestamp 1751914308
transform 1 0 29344 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1009_
timestamp 1751534193
transform 1 0 30688 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1010_
timestamp 1751914308
transform -1 0 30240 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1011_
timestamp 1751534193
transform 1 0 29456 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1012_
timestamp 1751532043
transform -1 0 40432 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1013_
timestamp 1751532043
transform -1 0 36400 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1014_
timestamp 1751532043
transform -1 0 33824 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1015_
timestamp 1751532043
transform -1 0 33376 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1016_
timestamp 1751740063
transform -1 0 32704 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1017_
timestamp 1751532043
transform 1 0 33040 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1018_
timestamp 1751532043
transform -1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1019_
timestamp 1751532043
transform -1 0 36960 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1020_
timestamp 1751532043
transform 1 0 40656 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1021_
timestamp 1751532043
transform -1 0 41552 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1022_
timestamp 1751532043
transform -1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_4  _1023_
timestamp 1751830969
transform 1 0 30576 0 -1 20384
box -86 -86 1545 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1024_
timestamp 1751914308
transform 1 0 35280 0 1 17248
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1025_
timestamp 1751534193
transform 1 0 36848 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1026_
timestamp 1751914308
transform 1 0 36848 0 1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1027_
timestamp 1751534193
transform 1 0 38192 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1028_
timestamp 1751914308
transform 1 0 38304 0 1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1029_
timestamp 1751534193
transform 1 0 39424 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1030_
timestamp 1751914308
transform -1 0 40992 0 1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1031_
timestamp 1751534193
transform 1 0 39872 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_4  _1032_
timestamp 1751830969
transform 1 0 31248 0 -1 18816
box -86 -86 1545 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1033_
timestamp 1751914308
transform -1 0 40880 0 1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1034_
timestamp 1751534193
transform 1 0 40768 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1035_
timestamp 1751914308
transform -1 0 43680 0 1 17248
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1036_
timestamp 1751534193
transform 1 0 42560 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1037_
timestamp 1751914308
transform -1 0 42560 0 -1 17248
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1038_
timestamp 1751534193
transform 1 0 41664 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1039_
timestamp 1751914308
transform -1 0 44016 0 1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1040_
timestamp 1751534193
transform -1 0 42672 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1041_
timestamp 1751534193
transform -1 0 30352 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1042_
timestamp 1753182340
transform 1 0 28112 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1043_
timestamp 1751534193
transform 1 0 37744 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1044_
timestamp 1752061876
transform 1 0 29792 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1045_
timestamp 1751532043
transform -1 0 14336 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1046_
timestamp 1751532043
transform -1 0 13888 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1047_
timestamp 1751740063
transform 1 0 19936 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1048_
timestamp 1751532043
transform 1 0 16576 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1049_
timestamp 1751532043
transform 1 0 13328 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1050_
timestamp 1751532043
transform -1 0 11872 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1051_
timestamp 1751532043
transform -1 0 9968 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1052_
timestamp 1751532043
transform 1 0 10864 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1053_
timestamp 1751532043
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1054_
timestamp 1751534193
transform 1 0 25088 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1055_
timestamp 1751889808
transform -1 0 27440 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1056_
timestamp 1751740063
transform -1 0 29792 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1057_
timestamp 1751740063
transform 1 0 27552 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1058_
timestamp 1751740063
transform -1 0 29344 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1059_
timestamp 1753182340
transform 1 0 26544 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1060_
timestamp 1751534193
transform 1 0 27776 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1061_
timestamp 1751740063
transform -1 0 28336 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1062_
timestamp 1751740063
transform -1 0 28896 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1063_
timestamp 1753182340
transform 1 0 25312 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1064_
timestamp 1751534193
transform -1 0 24864 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1065_
timestamp 1751740063
transform -1 0 26880 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1066_
timestamp 1751740063
transform 1 0 27104 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1067_
timestamp 1753182340
transform 1 0 25760 0 -1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1068_
timestamp 1751534193
transform -1 0 26320 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1069_
timestamp 1751740063
transform -1 0 27552 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1070_
timestamp 1751740063
transform 1 0 26320 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1071_
timestamp 1753182340
transform 1 0 26432 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1072_
timestamp 1751534193
transform -1 0 25648 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1073_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751632746
transform -1 0 41440 0 1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1074_
timestamp 1751632746
transform 1 0 35392 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1075_
timestamp 1751632746
transform 1 0 35056 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1076_
timestamp 1751632746
transform 1 0 29680 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1077_
timestamp 1751632746
transform 1 0 30128 0 1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1078_
timestamp 1751632746
transform 1 0 40768 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1079_
timestamp 1751632746
transform 1 0 40768 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1080_
timestamp 1751632746
transform 1 0 40544 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1081_
timestamp 1751632746
transform -1 0 43792 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1082_
timestamp 1751632746
transform 1 0 40880 0 -1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1083_
timestamp 1751632746
transform 1 0 40768 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1084_
timestamp 1751632746
transform 1 0 39424 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1085_
timestamp 1751632746
transform 1 0 19712 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1086_
timestamp 1751632746
transform 1 0 19040 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1087_
timestamp 1751632746
transform 1 0 19152 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1088_
timestamp 1751632746
transform 1 0 24080 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1089_
timestamp 1751632746
transform 1 0 25088 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1090_
timestamp 1751632746
transform 1 0 25088 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1091_
timestamp 1751632746
transform 1 0 20720 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1092_
timestamp 1751632746
transform 1 0 19712 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1093_
timestamp 1751632746
transform 1 0 19600 0 -1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1094_
timestamp 1751632746
transform -1 0 22960 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1095_
timestamp 1751632746
transform 1 0 21392 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1096_
timestamp 1751632746
transform 1 0 28000 0 -1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1097_
timestamp 1751632746
transform 1 0 30240 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1098_
timestamp 1751632746
transform 1 0 26880 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1099_
timestamp 1751632746
transform -1 0 39872 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1100_
timestamp 1751632746
transform 1 0 34944 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1101_
timestamp 1751632746
transform 1 0 34944 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1102_
timestamp 1751632746
transform -1 0 35168 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1103_
timestamp 1751632746
transform 1 0 39872 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1104_
timestamp 1751632746
transform -1 0 9184 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1105_
timestamp 1751632746
transform 1 0 20832 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1106_
timestamp 1751632746
transform 1 0 21168 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1107_
timestamp 1751632746
transform 1 0 21168 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1108_
timestamp 1751632746
transform 1 0 20160 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1109_
timestamp 1751632746
transform 1 0 6048 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1110_
timestamp 1751632746
transform 1 0 9072 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1111_
timestamp 1751632746
transform 1 0 9520 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1112_
timestamp 1751632746
transform -1 0 13104 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1113_
timestamp 1751632746
transform 1 0 10976 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1114_
timestamp 1751632746
transform 1 0 13104 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1115_
timestamp 1751632746
transform 1 0 23744 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1116_
timestamp 1751632746
transform 1 0 22848 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1117_
timestamp 1751632746
transform 1 0 27664 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1118_
timestamp 1751632746
transform 1 0 26768 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1119_
timestamp 1751632746
transform 1 0 14000 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1120_
timestamp 1751632746
transform -1 0 18256 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1121_
timestamp 1751632746
transform 1 0 17248 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1122_
timestamp 1751632746
transform 1 0 12656 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1123_
timestamp 1751632746
transform 1 0 13440 0 -1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1124_
timestamp 1751632746
transform 1 0 14000 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1125_
timestamp 1751632746
transform 1 0 15120 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1126_
timestamp 1751632746
transform 1 0 17024 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1127_
timestamp 1751632746
transform 1 0 37184 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1128_
timestamp 1751632746
transform 1 0 40768 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1129_
timestamp 1751632746
transform 1 0 40880 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1130_
timestamp 1751632746
transform 1 0 40544 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1131_
timestamp 1751632746
transform 1 0 29680 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1132_
timestamp 1751632746
transform 1 0 33040 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1133_
timestamp 1751632746
transform 1 0 36064 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1134_
timestamp 1751632746
transform -1 0 39872 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1135_
timestamp 1751632746
transform -1 0 43792 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1136_
timestamp 1751632746
transform -1 0 22512 0 -1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1137_
timestamp 1751632746
transform 1 0 39872 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1138_
timestamp 1751632746
transform 1 0 36848 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1139_
timestamp 1751632746
transform 1 0 35392 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1140_
timestamp 1751632746
transform 1 0 33488 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1141_
timestamp 1751632746
transform 1 0 31696 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1142_
timestamp 1751632746
transform 1 0 29008 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1143_
timestamp 1751632746
transform -1 0 42672 0 1 3136
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1144_
timestamp 1751632746
transform 1 0 39872 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1145_
timestamp 1751632746
transform -1 0 44128 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1146_
timestamp 1751632746
transform -1 0 44128 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1147_
timestamp 1751632746
transform -1 0 20944 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1148_
timestamp 1751632746
transform 1 0 32928 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1149_
timestamp 1751632746
transform 1 0 32480 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1150_
timestamp 1751632746
transform 1 0 33488 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1151_
timestamp 1751632746
transform 1 0 7840 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1152_
timestamp 1751632746
transform 1 0 7504 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1153_
timestamp 1751632746
transform 1 0 9408 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1154_
timestamp 1751632746
transform 1 0 10080 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1155_
timestamp 1751632746
transform -1 0 9072 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1156_
timestamp 1751632746
transform 1 0 9408 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1157_
timestamp 1751632746
transform 1 0 9072 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1158_
timestamp 1751632746
transform 1 0 9408 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1159_
timestamp 1751632746
transform -1 0 12432 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1160_
timestamp 1751632746
transform 1 0 9408 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1161_
timestamp 1751632746
transform 1 0 21168 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1162_
timestamp 1751632746
transform -1 0 28784 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1163_
timestamp 1751632746
transform 1 0 25648 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1164_
timestamp 1751632746
transform 1 0 23408 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1165_
timestamp 1751632746
transform 1 0 8960 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1166_
timestamp 1751632746
transform -1 0 18032 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1167_
timestamp 1751632746
transform -1 0 17024 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1168_
timestamp 1751632746
transform 1 0 15344 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1169_
timestamp 1751632746
transform 1 0 15792 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1170_
timestamp 1751632746
transform -1 0 17024 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1171_
timestamp 1751632746
transform -1 0 17248 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1172_
timestamp 1751632746
transform 1 0 16016 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1173_
timestamp 1751632746
transform 1 0 17248 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1174_
timestamp 1751632746
transform 1 0 33376 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1175_
timestamp 1751632746
transform 1 0 36848 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1176_
timestamp 1751632746
transform 1 0 32928 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1177_
timestamp 1751632746
transform -1 0 17920 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1178_
timestamp 1751632746
transform 1 0 15792 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1179_
timestamp 1751632746
transform 1 0 16464 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1180_
timestamp 1751632746
transform 1 0 18816 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1181_
timestamp 1751632746
transform 1 0 14000 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1182_
timestamp 1751632746
transform 1 0 17920 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1183_
timestamp 1751632746
transform -1 0 22064 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1184_
timestamp 1751632746
transform 1 0 19040 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1185_
timestamp 1751632746
transform 1 0 19600 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1186_
timestamp 1751632746
transform -1 0 22288 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1187_
timestamp 1751632746
transform 1 0 25088 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1188_
timestamp 1751632746
transform 1 0 17920 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1189_
timestamp 1751632746
transform -1 0 28784 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1190_
timestamp 1751632746
transform 1 0 21840 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1191_
timestamp 1751632746
transform -1 0 28112 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1192_
timestamp 1751632746
transform -1 0 24080 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1193_
timestamp 1751632746
transform 1 0 25984 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1194_
timestamp 1751632746
transform 1 0 21728 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1195_
timestamp 1751632746
transform -1 0 27776 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1196_
timestamp 1751632746
transform 1 0 21168 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1197_
timestamp 1751632746
transform -1 0 32368 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1198_
timestamp 1751632746
transform -1 0 32144 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1199_
timestamp 1751632746
transform -1 0 32032 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1200_
timestamp 1751632746
transform -1 0 40544 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1201_
timestamp 1751632746
transform -1 0 37296 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1202_
timestamp 1751632746
transform 1 0 32928 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1203_
timestamp 1751632746
transform 1 0 32816 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1204_
timestamp 1751632746
transform 1 0 29904 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1205_
timestamp 1751632746
transform 1 0 33600 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1206_
timestamp 1751632746
transform 1 0 35056 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1207_
timestamp 1751632746
transform 1 0 37856 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1208_
timestamp 1751632746
transform 1 0 40880 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1209_
timestamp 1751632746
transform 1 0 41104 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1210_
timestamp 1751632746
transform 1 0 29456 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1211_
timestamp 1751632746
transform 1 0 41104 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1212_
timestamp 1751632746
transform -1 0 39536 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1213_
timestamp 1751632746
transform -1 0 38752 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1214_
timestamp 1751632746
transform -1 0 40544 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1215_
timestamp 1751632746
transform 1 0 39648 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1216_
timestamp 1751632746
transform 1 0 39312 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1217_
timestamp 1751632746
transform 1 0 40880 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1218_
timestamp 1751632746
transform 1 0 40768 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1219_
timestamp 1751632746
transform 1 0 41104 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1220_
timestamp 1751632746
transform 1 0 39536 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1221_
timestamp 1751632746
transform 1 0 39648 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1222_
timestamp 1751632746
transform 1 0 14336 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1223_
timestamp 1751632746
transform 1 0 14000 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1224_
timestamp 1751632746
transform 1 0 21168 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1225_
timestamp 1751632746
transform 1 0 17248 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1226_
timestamp 1751632746
transform 1 0 13776 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1227_
timestamp 1751632746
transform 1 0 10752 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1228_
timestamp 1751632746
transform 1 0 10080 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1229_
timestamp 1751632746
transform -1 0 13104 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1230_
timestamp 1751632746
transform 1 0 17360 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1231_
timestamp 1751632746
transform 1 0 26992 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1232_
timestamp 1751632746
transform 1 0 24528 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1233_
timestamp 1751632746
transform 1 0 25536 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1234_
timestamp 1751632746
transform -1 0 26432 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1235_
timestamp 1751534193
transform 1 0 42336 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1236_
timestamp 1751534193
transform -1 0 43792 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1237_
timestamp 1751534193
transform -1 0 43568 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1238_
timestamp 1751534193
transform 1 0 42448 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1239_
timestamp 1751534193
transform 1 0 43568 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0532__B dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform -1 0 18704 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0541__A
timestamp 1751532392
transform 1 0 31248 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0544__A
timestamp 1751532392
transform 1 0 32592 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0546__B
timestamp 1751532392
transform 1 0 31920 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0551__B
timestamp 1751532392
transform 1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0685__B
timestamp 1751532392
transform 1 0 31472 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0713__A
timestamp 1751532392
transform 1 0 31136 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0754__A
timestamp 1751532392
transform -1 0 39984 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0755__A
timestamp 1751532392
transform 1 0 23408 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0757__A
timestamp 1751532392
transform -1 0 42000 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0758__A
timestamp 1751532392
transform 1 0 22736 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0760__A
timestamp 1751532392
transform -1 0 43680 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0761__A
timestamp 1751532392
transform 1 0 22736 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0862__A
timestamp 1751532392
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0864__A
timestamp 1751532392
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0866__A
timestamp 1751532392
transform -1 0 31472 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0868__A
timestamp 1751532392
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0869__A
timestamp 1751532392
transform -1 0 26656 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0891__A
timestamp 1751532392
transform 1 0 40208 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0893__A
timestamp 1751532392
transform 1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0895__A
timestamp 1751532392
transform 1 0 43568 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0897__A
timestamp 1751532392
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0899__A
timestamp 1751532392
transform 1 0 40992 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0902__A
timestamp 1751532392
transform -1 0 33600 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0904__A
timestamp 1751532392
transform -1 0 43680 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0906__A
timestamp 1751532392
transform 1 0 36064 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0908__A
timestamp 1751532392
transform 1 0 44128 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0910__A
timestamp 1751532392
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0912__A
timestamp 1751532392
transform 1 0 36288 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0928__A
timestamp 1751532392
transform 1 0 33936 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0930__A
timestamp 1751532392
transform 1 0 35728 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0932__A
timestamp 1751532392
transform 1 0 34720 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0949__A
timestamp 1751532392
transform 1 0 17024 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0951__A
timestamp 1751532392
transform 1 0 19600 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0953__A
timestamp 1751532392
transform -1 0 19040 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0955__A
timestamp 1751532392
transform -1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0959__A
timestamp 1751532392
transform 1 0 16016 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0961__A
timestamp 1751532392
transform -1 0 18368 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0963__A
timestamp 1751532392
transform 1 0 19488 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0971__A
timestamp 1751532392
transform 1 0 36288 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0990__A
timestamp 1751532392
transform 1 0 26320 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0997__S
timestamp 1751532392
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0999__A
timestamp 1751532392
transform 1 0 27104 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0999__S
timestamp 1751532392
transform 1 0 27552 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1001__S
timestamp 1751532392
transform 1 0 28560 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1003__S
timestamp 1751532392
transform 1 0 24192 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1008__A
timestamp 1751532392
transform -1 0 31808 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1030__A
timestamp 1751532392
transform 1 0 41216 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1039__A
timestamp 1751532392
transform 1 0 44128 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1043__A
timestamp 1751532392
transform 1 0 37520 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1052__A
timestamp 1751532392
transform -1 0 10416 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1056__A
timestamp 1751532392
transform 1 0 32256 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1062__A
timestamp 1751532392
transform -1 0 32144 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1065__A
timestamp 1751532392
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1069__A
timestamp 1751532392
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1089__CLK
timestamp 1751532392
transform 1 0 28560 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1090__CLK
timestamp 1751532392
transform 1 0 29120 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1094__CLK
timestamp 1751532392
transform 1 0 23184 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1095__CLK
timestamp 1751532392
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1098__CLK
timestamp 1751532392
transform 1 0 25872 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1136__CLK
timestamp 1751532392
transform -1 0 22960 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1142__CLK
timestamp 1751532392
transform 1 0 28784 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1155__CLK
timestamp 1751532392
transform 1 0 7952 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1181__CLK
timestamp 1751532392
transform 1 0 17024 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1204__CLK
timestamp 1751532392
transform 1 0 29680 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1220__D
timestamp 1751532392
transform 1 0 42784 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1221__CLK
timestamp 1751532392
transform 1 0 39424 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1221__D
timestamp 1751532392
transform 1 0 42896 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1751532392
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload0_A
timestamp 1751532392
transform 1 0 27888 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_fanout20_A
timestamp 1751532392
transform 1 0 19376 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input1_A
timestamp 1751532392
transform -1 0 44352 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input2_A
timestamp 1751532392
transform -1 0 43680 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input3_A
timestamp 1751532392
transform -1 0 44352 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input4_A
timestamp 1751532392
transform -1 0 44352 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input5_A
timestamp 1751532392
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0209_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751661108
transform 1 0 23296 0 1 21952
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0210_
timestamp 1751661108
transform 1 0 25312 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0228_
timestamp 1751661108
transform 1 0 33152 0 1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0229_
timestamp 1751661108
transform 1 0 36848 0 1 26656
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0230_
timestamp 1751661108
transform 1 0 40880 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0231_
timestamp 1751661108
transform 1 0 35952 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0254_
timestamp 1751661108
transform 1 0 19040 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0255_
timestamp 1751661108
transform 1 0 21168 0 1 9408
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0256_
timestamp 1751661108
transform 1 0 20608 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0257_
timestamp 1751661108
transform -1 0 20944 0 1 9408
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0282_
timestamp 1751661108
transform -1 0 13888 0 -1 23520
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0283_
timestamp 1751661108
transform -1 0 9184 0 -1 18816
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0284_
timestamp 1751661108
transform 1 0 9744 0 -1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0285_
timestamp 1751661108
transform -1 0 15232 0 -1 20384
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0310_
timestamp 1751661108
transform 1 0 33264 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0311_
timestamp 1751661108
transform 1 0 37408 0 1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0312_
timestamp 1751661108
transform 1 0 41552 0 -1 6272
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0__0313_
timestamp 1751661108
transform 1 0 36512 0 -1 9408
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0_clk
timestamp 1751661108
transform -1 0 34608 0 1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0209_
timestamp 1751661108
transform -1 0 24080 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0210_
timestamp 1751661108
transform -1 0 24192 0 -1 23520
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0228_
timestamp 1751661108
transform -1 0 32704 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0229_
timestamp 1751661108
transform -1 0 32704 0 -1 28224
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0230_
timestamp 1751661108
transform -1 0 40544 0 -1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0231_
timestamp 1751661108
transform -1 0 35280 0 1 28224
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0254_
timestamp 1751661108
transform 1 0 21840 0 -1 9408
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0255_
timestamp 1751661108
transform -1 0 20384 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0256_
timestamp 1751661108
transform 1 0 24416 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0257_
timestamp 1751661108
transform 1 0 21168 0 1 6272
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0282_
timestamp 1751661108
transform -1 0 9968 0 1 21952
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0283_
timestamp 1751661108
transform 1 0 9968 0 1 14112
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0284_
timestamp 1751661108
transform -1 0 12544 0 1 10976
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0285_
timestamp 1751661108
transform -1 0 14448 0 -1 18816
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0310_
timestamp 1751661108
transform -1 0 32144 0 -1 10976
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0311_
timestamp 1751661108
transform -1 0 39648 0 1 10976
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0312_
timestamp 1751661108
transform -1 0 40544 0 -1 6272
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_0__f__0313_
timestamp 1751661108
transform -1 0 35728 0 1 10976
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0209_
timestamp 1751661108
transform 1 0 25312 0 -1 21952
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0210_
timestamp 1751661108
transform 1 0 29008 0 1 23520
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0228_
timestamp 1751661108
transform 1 0 36848 0 1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0229_
timestamp 1751661108
transform 1 0 40768 0 -1 26656
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0230_
timestamp 1751661108
transform 1 0 41552 0 1 23520
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0231_
timestamp 1751661108
transform 1 0 39648 0 1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0254_
timestamp 1751661108
transform 1 0 21168 0 1 14112
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0255_
timestamp 1751661108
transform -1 0 18144 0 1 9408
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0256_
timestamp 1751661108
transform -1 0 23968 0 1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0257_
timestamp 1751661108
transform 1 0 21168 0 1 10976
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0282_
timestamp 1751661108
transform 1 0 15008 0 1 21952
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0283_
timestamp 1751661108
transform 1 0 8624 0 1 18816
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0284_
timestamp 1751661108
transform 1 0 12432 0 -1 17248
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0285_
timestamp 1751661108
transform -1 0 13216 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0310_
timestamp 1751661108
transform 1 0 37184 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0311_
timestamp 1751661108
transform 1 0 40768 0 -1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0312_
timestamp 1751661108
transform 1 0 38304 0 1 6272
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_1_1__f__0313_
timestamp 1751661108
transform 1 0 40208 0 1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_0__f_clk
timestamp 1751661108
transform -1 0 28448 0 -1 34496
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_1__f_clk
timestamp 1751661108
transform -1 0 30912 0 -1 39200
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_2__f_clk
timestamp 1751661108
transform 1 0 37744 0 -1 34496
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_3__f_clk
timestamp 1751661108
transform 1 0 36848 0 1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_8  clkload0 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752063729
transform 1 0 25648 0 1 34496
box -86 -86 2102 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751558652
transform 1 0 27552 0 1 37632
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751633659
transform 1 0 38080 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload3
timestamp 1751558652
transform -1 0 26656 0 1 20384
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload4
timestamp 1751558652
transform 1 0 18256 0 -1 4704
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload5
timestamp 1751558652
transform -1 0 28784 0 1 23520
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload6
timestamp 1751558652
transform -1 0 44016 0 1 7840
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload7
timestamp 1751558652
transform 1 0 8960 0 1 14112
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload8
timestamp 1751558652
transform 1 0 39648 0 1 26656
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout11
timestamp 1751534193
transform 1 0 20272 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout12
timestamp 1751534193
transform -1 0 9184 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout13
timestamp 1751534193
transform 1 0 13328 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout14
timestamp 1751534193
transform -1 0 12208 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout15
timestamp 1751534193
transform -1 0 17808 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout16
timestamp 1751534193
transform -1 0 18480 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout17
timestamp 1751534193
transform -1 0 16240 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout18
timestamp 1751534193
transform 1 0 18480 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout19
timestamp 1751534193
transform -1 0 14560 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout20
timestamp 1751534193
transform -1 0 20944 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout21
timestamp 1751534193
transform -1 0 20272 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout22
timestamp 1751534193
transform -1 0 16016 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout23
timestamp 1751534193
transform -1 0 21840 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout24
timestamp 1751534193
transform -1 0 27328 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout25
timestamp 1751534193
transform -1 0 25760 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout26
timestamp 1751534193
transform 1 0 26096 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout27
timestamp 1751534193
transform 1 0 27664 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout28
timestamp 1751534193
transform -1 0 15792 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout29
timestamp 1751534193
transform 1 0 18368 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout30
timestamp 1751534193
transform -1 0 19712 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout31
timestamp 1751534193
transform -1 0 24192 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout32
timestamp 1751534193
transform 1 0 24192 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout33
timestamp 1751534193
transform -1 0 24304 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout34
timestamp 1751534193
transform -1 0 23632 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout35
timestamp 1751534193
transform -1 0 29232 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout36
timestamp 1751534193
transform -1 0 31584 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout37
timestamp 1751534193
transform -1 0 37184 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout38
timestamp 1751534193
transform 1 0 37296 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout39
timestamp 1751534193
transform 1 0 30240 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout40
timestamp 1751534193
transform -1 0 32032 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout41
timestamp 1751534193
transform 1 0 35504 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout42
timestamp 1751534193
transform -1 0 40208 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout43
timestamp 1751534193
transform 1 0 34832 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout44
timestamp 1751534193
transform -1 0 29792 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout45
timestamp 1751534193
transform 1 0 31360 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout46
timestamp 1751534193
transform 1 0 24192 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532351
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_18
timestamp 1751532351
transform 1 0 3360 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_36
timestamp 1751532351
transform 1 0 5376 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_52
timestamp 1751532351
transform 1 0 7168 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_70
timestamp 1751532351
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_86
timestamp 1751532351
transform 1 0 10976 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_104
timestamp 1751532351
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_120
timestamp 1751532351
transform 1 0 14784 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532440
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_140 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532423
transform 1 0 17024 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_197 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_201
timestamp 1751532440
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_203
timestamp 1751532423
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_231
timestamp 1751532246
transform 1 0 27216 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_235
timestamp 1751532423
transform 1 0 27664 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_252
timestamp 1751532351
transform 1 0 29568 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_268
timestamp 1751532246
transform 1 0 31360 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_274
timestamp 1751532351
transform 1 0 32032 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_290
timestamp 1751532246
transform 1 0 33824 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_300
timestamp 1751532246
transform 1 0 34944 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_304
timestamp 1751532440
transform 1 0 35392 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_308
timestamp 1751532246
transform 1 0 35840 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_312
timestamp 1751532423
transform 1 0 36288 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_319 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532312
transform 1 0 37072 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_327
timestamp 1751532246
transform 1 0 37968 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_373
timestamp 1751532423
transform 1 0 43120 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_383
timestamp 1751532423
transform 1 0 44240 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_2
timestamp 1751532351
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_18
timestamp 1751532351
transform 1 0 3360 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_34
timestamp 1751532351
transform 1 0 5152 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_50
timestamp 1751532351
transform 1 0 6944 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_66
timestamp 1751532246
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_72
timestamp 1751532351
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_88
timestamp 1751532351
transform 1 0 11200 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_104
timestamp 1751532351
transform 1 0 12992 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_120
timestamp 1751532351
transform 1 0 14784 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_136
timestamp 1751532246
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_142
timestamp 1751532440
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_194
timestamp 1751532351
transform 1 0 23072 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_212
timestamp 1751532312
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_247
timestamp 1751532246
transform 1 0 29008 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_263
timestamp 1751532351
transform 1 0 30800 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_279
timestamp 1751532423
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_282
timestamp 1751532246
transform 1 0 32928 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_313
timestamp 1751532440
transform 1 0 36400 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_315
timestamp 1751532423
transform 1 0 36624 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_334
timestamp 1751532440
transform 1 0 38752 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_352
timestamp 1751532440
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_354
timestamp 1751532423
transform 1 0 40992 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_382
timestamp 1751532440
transform 1 0 44128 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_2
timestamp 1751532351
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_18
timestamp 1751532351
transform 1 0 3360 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_34
timestamp 1751532423
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_37
timestamp 1751532351
transform 1 0 5488 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_53
timestamp 1751532351
transform 1 0 7280 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_69
timestamp 1751532351
transform 1 0 9072 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_85
timestamp 1751532351
transform 1 0 10864 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_101
timestamp 1751532246
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_107
timestamp 1751532312
transform 1 0 13328 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_115
timestamp 1751532246
transform 1 0 14224 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_119
timestamp 1751532440
transform 1 0 14672 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_181
timestamp 1751532423
transform 1 0 21616 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_242
timestamp 1751532440
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_244
timestamp 1751532423
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_247
timestamp 1751532440
transform 1 0 29008 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_249
timestamp 1751532423
transform 1 0 29232 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_277
timestamp 1751532246
transform 1 0 32368 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_281
timestamp 1751532423
transform 1 0 32816 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_2
timestamp 1751532351
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_18
timestamp 1751532351
transform 1 0 3360 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_34
timestamp 1751532351
transform 1 0 5152 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_50
timestamp 1751532351
transform 1 0 6944 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_66
timestamp 1751532246
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_72
timestamp 1751532351
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_88
timestamp 1751532351
transform 1 0 11200 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_104
timestamp 1751532351
transform 1 0 12992 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_120
timestamp 1751532312
transform 1 0 14784 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_128
timestamp 1751532246
transform 1 0 15680 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_212
timestamp 1751532423
transform 1 0 25088 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_233
timestamp 1751532423
transform 1 0 27440 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_275
timestamp 1751532246
transform 1 0 32144 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_279
timestamp 1751532423
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_282
timestamp 1751532246
transform 1 0 32928 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_286
timestamp 1751532440
transform 1 0 33376 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_300
timestamp 1751532440
transform 1 0 34944 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_316
timestamp 1751532423
transform 1 0 36736 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_324
timestamp 1751532423
transform 1 0 37632 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_2
timestamp 1751532351
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_18
timestamp 1751532351
transform 1 0 3360 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_34
timestamp 1751532423
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_37
timestamp 1751532351
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_53
timestamp 1751532351
transform 1 0 7280 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_69
timestamp 1751532351
transform 1 0 9072 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_85
timestamp 1751532351
transform 1 0 10864 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_101
timestamp 1751532246
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_107
timestamp 1751532351
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_123
timestamp 1751532246
transform 1 0 15120 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_127
timestamp 1751532440
transform 1 0 15568 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_156
timestamp 1751532423
transform 1 0 18816 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_244
timestamp 1751532423
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_247
timestamp 1751532440
transform 1 0 29008 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_249
timestamp 1751532423
transform 1 0 29232 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_268
timestamp 1751532440
transform 1 0 31360 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_272
timestamp 1751532351
transform 1 0 31808 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_312
timestamp 1751532440
transform 1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_314
timestamp 1751532423
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_328
timestamp 1751532440
transform 1 0 38080 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_382
timestamp 1751532440
transform 1 0 44128 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_2
timestamp 1751532351
transform 1 0 1568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_18
timestamp 1751532351
transform 1 0 3360 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_34
timestamp 1751532351
transform 1 0 5152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_50
timestamp 1751532351
transform 1 0 6944 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_66
timestamp 1751532246
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_72
timestamp 1751532351
transform 1 0 9408 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_88
timestamp 1751532351
transform 1 0 11200 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_104
timestamp 1751532351
transform 1 0 12992 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_120
timestamp 1751532351
transform 1 0 14784 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_149
timestamp 1751532440
transform 1 0 18032 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_185
timestamp 1751532423
transform 1 0 22064 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_200
timestamp 1751532312
transform 1 0 23744 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_208
timestamp 1751532440
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_212
timestamp 1751532440
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_214
timestamp 1751532423
transform 1 0 25312 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_241
timestamp 1751532440
transform 1 0 28336 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_245
timestamp 1751532423
transform 1 0 28784 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_264
timestamp 1751532351
transform 1 0 30912 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_282
timestamp 1751532351
transform 1 0 32928 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_298
timestamp 1751532246
transform 1 0 34720 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_2
timestamp 1751532351
transform 1 0 1568 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_18
timestamp 1751532351
transform 1 0 3360 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_34
timestamp 1751532423
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_37
timestamp 1751532351
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_53
timestamp 1751532351
transform 1 0 7280 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_69
timestamp 1751532351
transform 1 0 9072 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_85
timestamp 1751532351
transform 1 0 10864 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_101
timestamp 1751532246
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_107
timestamp 1751532351
transform 1 0 13328 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_123
timestamp 1751532312
transform 1 0 15120 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_131
timestamp 1751532246
transform 1 0 16016 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_228
timestamp 1751532440
transform 1 0 26880 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_232
timestamp 1751532440
transform 1 0 27328 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_236
timestamp 1751532312
transform 1 0 27776 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_244
timestamp 1751532423
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_274
timestamp 1751532351
transform 1 0 32032 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_310
timestamp 1751532440
transform 1 0 36064 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_314
timestamp 1751532423
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_321
timestamp 1751532423
transform 1 0 37296 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_381
timestamp 1751532440
transform 1 0 44016 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_383
timestamp 1751532423
transform 1 0 44240 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_2
timestamp 1751532351
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_18
timestamp 1751532351
transform 1 0 3360 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_34
timestamp 1751532351
transform 1 0 5152 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_50
timestamp 1751532351
transform 1 0 6944 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_66
timestamp 1751532246
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_72
timestamp 1751532351
transform 1 0 9408 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_88
timestamp 1751532351
transform 1 0 11200 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_104
timestamp 1751532351
transform 1 0 12992 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_120
timestamp 1751532312
transform 1 0 14784 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_128
timestamp 1751532246
transform 1 0 15680 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_142
timestamp 1751532440
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_144
timestamp 1751532423
transform 1 0 17472 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_208
timestamp 1751532440
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_223
timestamp 1751532351
transform 1 0 26320 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_239
timestamp 1751532246
transform 1 0 28112 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_249
timestamp 1751532440
transform 1 0 29232 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_257
timestamp 1751532351
transform 1 0 30128 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_279
timestamp 1751532423
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_282
timestamp 1751532246
transform 1 0 32928 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_286
timestamp 1751532423
transform 1 0 33376 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_383
timestamp 1751532423
transform 1 0 44240 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_2
timestamp 1751532351
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_18
timestamp 1751532351
transform 1 0 3360 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_34
timestamp 1751532423
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_37
timestamp 1751532351
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_53
timestamp 1751532351
transform 1 0 7280 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_69
timestamp 1751532351
transform 1 0 9072 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_85
timestamp 1751532351
transform 1 0 10864 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_101
timestamp 1751532246
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_107
timestamp 1751532351
transform 1 0 13328 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_123
timestamp 1751532440
transform 1 0 15120 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_216
timestamp 1751532246
transform 1 0 25536 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_220
timestamp 1751532423
transform 1 0 25984 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_235
timestamp 1751532312
transform 1 0 27664 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_243
timestamp 1751532440
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_247
timestamp 1751532312
transform 1 0 29008 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_255
timestamp 1751532423
transform 1 0 29904 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_262
timestamp 1751532246
transform 1 0 30688 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_266
timestamp 1751532423
transform 1 0 31136 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_298
timestamp 1751532440
transform 1 0 34720 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_300
timestamp 1751532423
transform 1 0 34944 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_375
timestamp 1751532440
transform 1 0 43344 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_377
timestamp 1751532423
transform 1 0 43568 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_2
timestamp 1751532351
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_18
timestamp 1751532351
transform 1 0 3360 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_34
timestamp 1751532351
transform 1 0 5152 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_50
timestamp 1751532351
transform 1 0 6944 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_66
timestamp 1751532246
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_72
timestamp 1751532351
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_88
timestamp 1751532351
transform 1 0 11200 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_104
timestamp 1751532312
transform 1 0 12992 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_112
timestamp 1751532423
transform 1 0 13888 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_149
timestamp 1751532440
transform 1 0 18032 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_151
timestamp 1751532423
transform 1 0 18256 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_189
timestamp 1751532423
transform 1 0 22512 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_245
timestamp 1751532246
transform 1 0 28784 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_249
timestamp 1751532423
transform 1 0 29232 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_275
timestamp 1751532423
transform 1 0 32144 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_303
timestamp 1751532423
transform 1 0 35280 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_349
timestamp 1751532423
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_352
timestamp 1751532440
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_382
timestamp 1751532440
transform 1 0 44128 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_2
timestamp 1751532351
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_18
timestamp 1751532351
transform 1 0 3360 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_34
timestamp 1751532423
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_37
timestamp 1751532351
transform 1 0 5488 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_53
timestamp 1751532351
transform 1 0 7280 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_69
timestamp 1751532246
transform 1 0 9072 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_73
timestamp 1751532440
transform 1 0 9520 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_100
timestamp 1751532246
transform 1 0 12544 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_104
timestamp 1751532423
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_107
timestamp 1751532351
transform 1 0 13328 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_123
timestamp 1751532351
transform 1 0 15120 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_139
timestamp 1751532423
transform 1 0 16912 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_142
timestamp 1751532246
transform 1 0 17248 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_146
timestamp 1751532440
transform 1 0 17696 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_213
timestamp 1751532246
transform 1 0 25200 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_217
timestamp 1751532423
transform 1 0 25648 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_281
timestamp 1751532423
transform 1 0 32816 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_314
timestamp 1751532423
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_374
timestamp 1751532440
transform 1 0 43232 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_2
timestamp 1751532351
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_18
timestamp 1751532351
transform 1 0 3360 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_34
timestamp 1751532351
transform 1 0 5152 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_50
timestamp 1751532351
transform 1 0 6944 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_66
timestamp 1751532246
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_142
timestamp 1751532312
transform 1 0 17248 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_150
timestamp 1751532423
transform 1 0 18144 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_242
timestamp 1751532440
transform 1 0 28448 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_244
timestamp 1751532423
transform 1 0 28672 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_247
timestamp 1751532246
transform 1 0 29008 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_251
timestamp 1751532440
transform 1 0 29456 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_282
timestamp 1751532440
transform 1 0 32928 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_284
timestamp 1751532423
transform 1 0 33152 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_316
timestamp 1751532246
transform 1 0 36736 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_345
timestamp 1751532246
transform 1 0 39984 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_349
timestamp 1751532423
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_352
timestamp 1751532423
transform 1 0 40768 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_380
timestamp 1751532440
transform 1 0 43904 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_2
timestamp 1751532351
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_18
timestamp 1751532351
transform 1 0 3360 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_34
timestamp 1751532423
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_37
timestamp 1751532351
transform 1 0 5488 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_53
timestamp 1751532312
transform 1 0 7280 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_61
timestamp 1751532246
transform 1 0 8176 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_65
timestamp 1751532440
transform 1 0 8624 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_67
timestamp 1751532423
transform 1 0 8848 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_95
timestamp 1751532312
transform 1 0 11984 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_103
timestamp 1751532440
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_107
timestamp 1751532312
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_148
timestamp 1751532440
transform 1 0 17920 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_152
timestamp 1751532312
transform 1 0 18368 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_160
timestamp 1751532246
transform 1 0 19264 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_170
timestamp 1751532246
transform 1 0 20384 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_174
timestamp 1751532423
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_204
timestamp 1751532312
transform 1 0 24192 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_218
timestamp 1751532246
transform 1 0 25760 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_222
timestamp 1751532423
transform 1 0 26208 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_237
timestamp 1751532312
transform 1 0 27888 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_253
timestamp 1751532246
transform 1 0 29680 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_257
timestamp 1751532423
transform 1 0 30128 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_270
timestamp 1751532440
transform 1 0 31584 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_284
timestamp 1751532440
transform 1 0 33152 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_288
timestamp 1751532246
transform 1 0 33600 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_308
timestamp 1751532440
transform 1 0 35840 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_312
timestamp 1751532440
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_314
timestamp 1751532423
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_344
timestamp 1751532246
transform 1 0 39872 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_348
timestamp 1751532440
transform 1 0 40320 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_383
timestamp 1751532423
transform 1 0 44240 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_2
timestamp 1751532351
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_18
timestamp 1751532351
transform 1 0 3360 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_34
timestamp 1751532351
transform 1 0 5152 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_50
timestamp 1751532440
transform 1 0 6944 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_99
timestamp 1751532246
transform 1 0 12432 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_103
timestamp 1751532423
transform 1 0 12880 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_118
timestamp 1751532246
transform 1 0 14560 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_169
timestamp 1751532246
transform 1 0 20272 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_173
timestamp 1751532440
transform 1 0 20720 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_175
timestamp 1751532423
transform 1 0 20944 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_209
timestamp 1751532423
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_212
timestamp 1751532351
transform 1 0 25088 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_228
timestamp 1751532246
transform 1 0 26880 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_232
timestamp 1751532440
transform 1 0 27328 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_234
timestamp 1751532423
transform 1 0 27552 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_262
timestamp 1751532246
transform 1 0 30688 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_266
timestamp 1751532440
transform 1 0 31136 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_268
timestamp 1751532423
transform 1 0 31360 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_275
timestamp 1751532246
transform 1 0 32144 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_279
timestamp 1751532423
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_282
timestamp 1751532423
transform 1 0 32928 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_343
timestamp 1751532423
transform 1 0 39760 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_352
timestamp 1751532440
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_354
timestamp 1751532423
transform 1 0 40992 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_381
timestamp 1751532440
transform 1 0 44016 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_383
timestamp 1751532423
transform 1 0 44240 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_2
timestamp 1751532351
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_18
timestamp 1751532351
transform 1 0 3360 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_34
timestamp 1751532423
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_37
timestamp 1751532351
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_53
timestamp 1751532246
transform 1 0 7280 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_102
timestamp 1751532440
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_104
timestamp 1751532423
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_121
timestamp 1751532246
transform 1 0 14896 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_170
timestamp 1751532246
transform 1 0 20384 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_174
timestamp 1751532423
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_214
timestamp 1751532312
transform 1 0 25312 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_222
timestamp 1751532440
transform 1 0 26208 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_244
timestamp 1751532423
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_265
timestamp 1751532440
transform 1 0 31024 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_269
timestamp 1751532351
transform 1 0 31472 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_285
timestamp 1751532440
transform 1 0 33264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_287
timestamp 1751532423
transform 1 0 33488 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_294
timestamp 1751532246
transform 1 0 34272 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_310
timestamp 1751532440
transform 1 0 36064 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_314
timestamp 1751532423
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_329
timestamp 1751532440
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_337
timestamp 1751532312
transform 1 0 39088 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_345
timestamp 1751532246
transform 1 0 39984 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_349
timestamp 1751532440
transform 1 0 40432 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_351
timestamp 1751532423
transform 1 0 40656 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_379
timestamp 1751532440
transform 1 0 43792 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_383
timestamp 1751532423
transform 1 0 44240 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_2
timestamp 1751532351
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_18
timestamp 1751532351
transform 1 0 3360 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_34
timestamp 1751532351
transform 1 0 5152 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_50
timestamp 1751532440
transform 1 0 6944 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_72
timestamp 1751532440
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_74
timestamp 1751532423
transform 1 0 9632 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_104
timestamp 1751532423
transform 1 0 12992 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_131
timestamp 1751532440
transform 1 0 16016 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_133
timestamp 1751532423
transform 1 0 16240 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_160
timestamp 1751532440
transform 1 0 19264 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_164
timestamp 1751532312
transform 1 0 19712 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_172
timestamp 1751532246
transform 1 0 20608 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_176
timestamp 1751532423
transform 1 0 21056 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_183
timestamp 1751532423
transform 1 0 21840 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_202
timestamp 1751532440
transform 1 0 23968 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_206
timestamp 1751532246
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_212
timestamp 1751532440
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_216
timestamp 1751532246
transform 1 0 25536 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_220
timestamp 1751532423
transform 1 0 25984 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_271
timestamp 1751532440
transform 1 0 31696 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_275
timestamp 1751532246
transform 1 0 32144 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_279
timestamp 1751532423
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_288
timestamp 1751532246
transform 1 0 33600 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_292
timestamp 1751532440
transform 1 0 34048 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_300
timestamp 1751532440
transform 1 0 34944 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_308
timestamp 1751532246
transform 1 0 35840 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_347
timestamp 1751532440
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_349
timestamp 1751532423
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_352
timestamp 1751532246
transform 1 0 40768 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_356
timestamp 1751532423
transform 1 0 41216 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_375
timestamp 1751532440
transform 1 0 43344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_379
timestamp 1751532246
transform 1 0 43792 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_383
timestamp 1751532423
transform 1 0 44240 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_2
timestamp 1751532351
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_18
timestamp 1751532351
transform 1 0 3360 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_34
timestamp 1751532423
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_37
timestamp 1751532351
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_53
timestamp 1751532246
transform 1 0 7280 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_57
timestamp 1751532423
transform 1 0 7728 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_121
timestamp 1751532246
transform 1 0 14896 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_152
timestamp 1751532312
transform 1 0 18368 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_166
timestamp 1751532312
transform 1 0 19936 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_174
timestamp 1751532423
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_177
timestamp 1751532312
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_185
timestamp 1751532246
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_189
timestamp 1751532440
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_191
timestamp 1751532423
transform 1 0 22736 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_219
timestamp 1751532440
transform 1 0 25872 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_261
timestamp 1751532440
transform 1 0 30576 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_263
timestamp 1751532423
transform 1 0 30800 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_277
timestamp 1751532440
transform 1 0 32368 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_281
timestamp 1751532246
transform 1 0 32816 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_285
timestamp 1751532440
transform 1 0 33264 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_299
timestamp 1751532440
transform 1 0 34832 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_307
timestamp 1751532312
transform 1 0 35728 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_317
timestamp 1751532246
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_339
timestamp 1751532246
transform 1 0 39312 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_345
timestamp 1751532440
transform 1 0 39984 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_349
timestamp 1751532351
transform 1 0 40432 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_365
timestamp 1751532312
transform 1 0 42224 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_373
timestamp 1751532440
transform 1 0 43120 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_375
timestamp 1751532423
transform 1 0 43344 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_378
timestamp 1751532246
transform 1 0 43680 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_2
timestamp 1751532351
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_18
timestamp 1751532351
transform 1 0 3360 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_34
timestamp 1751532351
transform 1 0 5152 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_50
timestamp 1751532312
transform 1 0 6944 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_58
timestamp 1751532440
transform 1 0 7840 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_64
timestamp 1751532440
transform 1 0 8512 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_124
timestamp 1751532246
transform 1 0 15232 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_128
timestamp 1751532440
transform 1 0 15680 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_130
timestamp 1751532423
transform 1 0 15904 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_133
timestamp 1751532423
transform 1 0 16240 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_154
timestamp 1751532312
transform 1 0 18592 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_162
timestamp 1751532440
transform 1 0 19488 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_191
timestamp 1751532423
transform 1 0 22736 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_212
timestamp 1751532423
transform 1 0 25088 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_266
timestamp 1751532423
transform 1 0 31136 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_278
timestamp 1751532440
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_282
timestamp 1751532351
transform 1 0 32928 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_312
timestamp 1751532351
transform 1 0 36288 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_328
timestamp 1751532312
transform 1 0 38080 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_336
timestamp 1751532423
transform 1 0 38976 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_349
timestamp 1751532423
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_352
timestamp 1751532440
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_374
timestamp 1751532440
transform 1 0 43232 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_2
timestamp 1751532351
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_18
timestamp 1751532351
transform 1 0 3360 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_34
timestamp 1751532423
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_37
timestamp 1751532351
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_53
timestamp 1751532440
transform 1 0 7280 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_82
timestamp 1751532312
transform 1 0 10528 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_104
timestamp 1751532423
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_121
timestamp 1751532312
transform 1 0 14896 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_162
timestamp 1751532246
transform 1 0 19488 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_166
timestamp 1751532440
transform 1 0 19936 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_168
timestamp 1751532423
transform 1 0 20160 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_188
timestamp 1751532312
transform 1 0 22400 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_196
timestamp 1751532440
transform 1 0 23296 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_225
timestamp 1751532440
transform 1 0 26544 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_227
timestamp 1751532423
transform 1 0 26768 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_247
timestamp 1751532440
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_249
timestamp 1751532423
transform 1 0 29232 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_264
timestamp 1751532440
transform 1 0 30912 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_266
timestamp 1751532423
transform 1 0 31136 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_287
timestamp 1751532440
transform 1 0 33488 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_289
timestamp 1751532423
transform 1 0 33712 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_302
timestamp 1751532423
transform 1 0 35168 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_323
timestamp 1751532351
transform 1 0 37520 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_2
timestamp 1751532351
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_18
timestamp 1751532351
transform 1 0 3360 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_34
timestamp 1751532312
transform 1 0 5152 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_42
timestamp 1751532440
transform 1 0 6048 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_44
timestamp 1751532423
transform 1 0 6272 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_72
timestamp 1751532423
transform 1 0 9408 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_91
timestamp 1751532423
transform 1 0 11536 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_128
timestamp 1751532246
transform 1 0 15680 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_132
timestamp 1751532440
transform 1 0 16128 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_154
timestamp 1751532440
transform 1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_197
timestamp 1751532423
transform 1 0 23408 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_218
timestamp 1751532440
transform 1 0 25760 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_251
timestamp 1751532246
transform 1 0 29456 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_255
timestamp 1751532423
transform 1 0 29904 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_263
timestamp 1751532246
transform 1 0 30800 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_282
timestamp 1751532246
transform 1 0 32928 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_286
timestamp 1751532423
transform 1 0 33376 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_347
timestamp 1751532440
transform 1 0 40208 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_349
timestamp 1751532423
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_379
timestamp 1751532440
transform 1 0 43792 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_381
timestamp 1751532423
transform 1 0 44016 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_2
timestamp 1751532351
transform 1 0 1568 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_18
timestamp 1751532351
transform 1 0 3360 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_34
timestamp 1751532423
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_37
timestamp 1751532351
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_53
timestamp 1751532312
transform 1 0 7280 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_90
timestamp 1751532423
transform 1 0 11424 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_132
timestamp 1751532312
transform 1 0 16128 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_142
timestamp 1751532351
transform 1 0 17248 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_158
timestamp 1751532351
transform 1 0 19040 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_174
timestamp 1751532423
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_189
timestamp 1751532440
transform 1 0 22512 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_193
timestamp 1751532246
transform 1 0 22960 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_199
timestamp 1751532423
transform 1 0 23632 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_241
timestamp 1751532440
transform 1 0 28336 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_254
timestamp 1751532351
transform 1 0 29792 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_270
timestamp 1751532351
transform 1 0 31584 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_286
timestamp 1751532246
transform 1 0 33376 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_290
timestamp 1751532423
transform 1 0 33824 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_311
timestamp 1751532246
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_335
timestamp 1751532246
transform 1 0 38864 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_339
timestamp 1751532440
transform 1 0 39312 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_380
timestamp 1751532440
transform 1 0 43904 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_2
timestamp 1751532351
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_18
timestamp 1751532351
transform 1 0 3360 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_34
timestamp 1751532351
transform 1 0 5152 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_50
timestamp 1751532312
transform 1 0 6944 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_58
timestamp 1751532423
transform 1 0 7840 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_68
timestamp 1751532440
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_124
timestamp 1751532246
transform 1 0 15232 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_148
timestamp 1751532312
transform 1 0 17920 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_156
timestamp 1751532440
transform 1 0 18816 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_158
timestamp 1751532423
transform 1 0 19040 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_192
timestamp 1751532312
transform 1 0 22848 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_200
timestamp 1751532246
transform 1 0 23744 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_206
timestamp 1751532440
transform 1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_224
timestamp 1751532440
transform 1 0 26432 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_237
timestamp 1751532440
transform 1 0 27888 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_250
timestamp 1751532440
transform 1 0 29344 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_252
timestamp 1751532423
transform 1 0 29568 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_259
timestamp 1751532440
transform 1 0 30352 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_274
timestamp 1751532246
transform 1 0 32032 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_278
timestamp 1751532440
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_306
timestamp 1751532423
transform 1 0 35616 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_334
timestamp 1751532312
transform 1 0 38752 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_342
timestamp 1751532440
transform 1 0 39648 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_358
timestamp 1751532440
transform 1 0 41440 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_2
timestamp 1751532351
transform 1 0 1568 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_18
timestamp 1751532351
transform 1 0 3360 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_34
timestamp 1751532423
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_37
timestamp 1751532246
transform 1 0 5488 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_41
timestamp 1751532423
transform 1 0 5936 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_103
timestamp 1751532440
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_107
timestamp 1751532423
transform 1 0 13328 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_161
timestamp 1751532440
transform 1 0 19376 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_165
timestamp 1751532246
transform 1 0 19824 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_189
timestamp 1751532440
transform 1 0 22512 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_193
timestamp 1751532312
transform 1 0 22960 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_201
timestamp 1751532246
transform 1 0 23856 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_205
timestamp 1751532440
transform 1 0 24304 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_226
timestamp 1751532423
transform 1 0 26656 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_241
timestamp 1751532440
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_247
timestamp 1751532423
transform 1 0 29008 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_264
timestamp 1751532440
transform 1 0 30912 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_266
timestamp 1751532423
transform 1 0 31136 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_269
timestamp 1751532440
transform 1 0 31472 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_271
timestamp 1751532423
transform 1 0 31696 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_305
timestamp 1751532440
transform 1 0 35504 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_309
timestamp 1751532246
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_313
timestamp 1751532440
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_317
timestamp 1751532312
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_325
timestamp 1751532246
transform 1 0 37744 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_329
timestamp 1751532423
transform 1 0 38192 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_354
timestamp 1751532440
transform 1 0 40992 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_358
timestamp 1751532440
transform 1 0 41440 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_360
timestamp 1751532423
transform 1 0 41664 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_381
timestamp 1751532440
transform 1 0 44016 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_383
timestamp 1751532423
transform 1 0 44240 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_2
timestamp 1751532351
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_18
timestamp 1751532351
transform 1 0 3360 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_34
timestamp 1751532351
transform 1 0 5152 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_50
timestamp 1751532312
transform 1 0 6944 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_58
timestamp 1751532440
transform 1 0 7840 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_142
timestamp 1751532440
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_144
timestamp 1751532423
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_151
timestamp 1751532423
transform 1 0 18256 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_178
timestamp 1751532351
transform 1 0 21280 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_194
timestamp 1751532246
transform 1 0 23072 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_198
timestamp 1751532423
transform 1 0 23520 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_206
timestamp 1751532246
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_212
timestamp 1751532440
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_246
timestamp 1751532423
transform 1 0 28896 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_267
timestamp 1751532440
transform 1 0 31248 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_271
timestamp 1751532440
transform 1 0 31696 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_275
timestamp 1751532246
transform 1 0 32144 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_279
timestamp 1751532423
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_309
timestamp 1751532312
transform 1 0 35952 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_317
timestamp 1751532246
transform 1 0 36848 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_321
timestamp 1751532440
transform 1 0 37296 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_352
timestamp 1751532440
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_354
timestamp 1751532423
transform 1 0 40992 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_382
timestamp 1751532440
transform 1 0 44128 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_2
timestamp 1751532351
transform 1 0 1568 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_18
timestamp 1751532351
transform 1 0 3360 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_34
timestamp 1751532423
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_37
timestamp 1751532312
transform 1 0 5488 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_45
timestamp 1751532246
transform 1 0 6384 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_49
timestamp 1751532440
transform 1 0 6832 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_51
timestamp 1751532423
transform 1 0 7056 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_77
timestamp 1751532423
transform 1 0 9968 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_107
timestamp 1751532423
transform 1 0 13328 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_147
timestamp 1751532312
transform 1 0 17808 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_155
timestamp 1751532246
transform 1 0 18704 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_159
timestamp 1751532440
transform 1 0 19152 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_177
timestamp 1751532312
transform 1 0 21168 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_185
timestamp 1751532440
transform 1 0 22064 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_193
timestamp 1751532440
transform 1 0 22960 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_195
timestamp 1751532423
transform 1 0 23184 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_241
timestamp 1751532440
transform 1 0 28336 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_274
timestamp 1751532440
transform 1 0 32032 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_278
timestamp 1751532312
transform 1 0 32480 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_286
timestamp 1751532440
transform 1 0 33376 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_294
timestamp 1751532246
transform 1 0 34272 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_298
timestamp 1751532440
transform 1 0 34720 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_314
timestamp 1751532423
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_383
timestamp 1751532423
transform 1 0 44240 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_2
timestamp 1751532351
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_18
timestamp 1751532351
transform 1 0 3360 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_34
timestamp 1751532351
transform 1 0 5152 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_50
timestamp 1751532351
transform 1 0 6944 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_66
timestamp 1751532246
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_79
timestamp 1751532423
transform 1 0 10192 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_118
timestamp 1751532246
transform 1 0 14560 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_122
timestamp 1751532423
transform 1 0 15008 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_129
timestamp 1751532246
transform 1 0 15792 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_139
timestamp 1751532423
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_142
timestamp 1751532351
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_158
timestamp 1751532312
transform 1 0 19040 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_166
timestamp 1751532440
transform 1 0 19936 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_204
timestamp 1751532246
transform 1 0 24192 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_208
timestamp 1751532440
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_290
timestamp 1751532312
transform 1 0 33824 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_352
timestamp 1751532423
transform 1 0 40768 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_381
timestamp 1751532440
transform 1 0 44016 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_383
timestamp 1751532423
transform 1 0 44240 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_2
timestamp 1751532351
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_18
timestamp 1751532351
transform 1 0 3360 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_34
timestamp 1751532423
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_37
timestamp 1751532351
transform 1 0 5488 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_53
timestamp 1751532351
transform 1 0 7280 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_69
timestamp 1751532312
transform 1 0 9072 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_77
timestamp 1751532440
transform 1 0 9968 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_103
timestamp 1751532440
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_107
timestamp 1751532351
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_123
timestamp 1751532440
transform 1 0 15120 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_125
timestamp 1751532423
transform 1 0 15344 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_133
timestamp 1751532246
transform 1 0 16240 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_144
timestamp 1751532312
transform 1 0 17472 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_152
timestamp 1751532423
transform 1 0 18368 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_166
timestamp 1751532312
transform 1 0 19936 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_174
timestamp 1751532423
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_204
timestamp 1751532440
transform 1 0 24192 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_206
timestamp 1751532423
transform 1 0 24416 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_234
timestamp 1751532440
transform 1 0 27552 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_278
timestamp 1751532440
transform 1 0 32480 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_280
timestamp 1751532423
transform 1 0 32704 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_317
timestamp 1751532440
transform 1 0 36848 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_319
timestamp 1751532423
transform 1 0 37072 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_2
timestamp 1751532351
transform 1 0 1568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_18
timestamp 1751532351
transform 1 0 3360 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_34
timestamp 1751532351
transform 1 0 5152 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_50
timestamp 1751532351
transform 1 0 6944 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_66
timestamp 1751532246
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_72
timestamp 1751532312
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_80
timestamp 1751532423
transform 1 0 10304 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_106
timestamp 1751532423
transform 1 0 13216 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_111
timestamp 1751532440
transform 1 0 13776 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_169
timestamp 1751532312
transform 1 0 20272 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_177
timestamp 1751532423
transform 1 0 21168 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_203
timestamp 1751532423
transform 1 0 24080 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_212
timestamp 1751532440
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_246
timestamp 1751532440
transform 1 0 28896 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_334
timestamp 1751532440
transform 1 0 38752 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_352
timestamp 1751532423
transform 1 0 40768 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_2
timestamp 1751532351
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_18
timestamp 1751532351
transform 1 0 3360 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_34
timestamp 1751532423
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_37
timestamp 1751532351
transform 1 0 5488 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_53
timestamp 1751532351
transform 1 0 7280 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_28_69
timestamp 1751532312
transform 1 0 9072 0 1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_77
timestamp 1751532423
transform 1 0 9968 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_107
timestamp 1751532423
transform 1 0 13328 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_170
timestamp 1751532423
transform 1 0 20384 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_28_204
timestamp 1751532312
transform 1 0 24192 0 1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_212
timestamp 1751532440
transform 1 0 25088 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_242
timestamp 1751532440
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_244
timestamp 1751532423
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_247
timestamp 1751532246
transform 1 0 29008 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_251
timestamp 1751532440
transform 1 0 29456 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_282
timestamp 1751532440
transform 1 0 32928 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_381
timestamp 1751532440
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_383
timestamp 1751532423
transform 1 0 44240 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_2
timestamp 1751532351
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_18
timestamp 1751532351
transform 1 0 3360 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_34
timestamp 1751532351
transform 1 0 5152 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_50
timestamp 1751532351
transform 1 0 6944 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_66
timestamp 1751532246
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_72
timestamp 1751532423
transform 1 0 9408 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_138
timestamp 1751532440
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_165
timestamp 1751532423
transform 1 0 19824 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_183
timestamp 1751532440
transform 1 0 21840 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_195
timestamp 1751532312
transform 1 0 23184 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_203
timestamp 1751532246
transform 1 0 24080 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_207
timestamp 1751532440
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_209
timestamp 1751532423
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_256
timestamp 1751532440
transform 1 0 30016 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_258
timestamp 1751532423
transform 1 0 30240 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_265
timestamp 1751532312
transform 1 0 31024 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_282
timestamp 1751532423
transform 1 0 32928 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_328
timestamp 1751532440
transform 1 0 38080 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_330
timestamp 1751532423
transform 1 0 38304 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_349
timestamp 1751532423
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_2
timestamp 1751532351
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_18
timestamp 1751532351
transform 1 0 3360 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_34
timestamp 1751532423
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_37
timestamp 1751532351
transform 1 0 5488 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_53
timestamp 1751532351
transform 1 0 7280 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_69
timestamp 1751532312
transform 1 0 9072 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_77
timestamp 1751532423
transform 1 0 9968 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_107
timestamp 1751532246
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_111
timestamp 1751532423
transform 1 0 13776 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_118
timestamp 1751532312
transform 1 0 14560 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_133
timestamp 1751532440
transform 1 0 16240 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_135
timestamp 1751532423
transform 1 0 16464 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_140
timestamp 1751532312
transform 1 0 17024 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_148
timestamp 1751532246
transform 1 0 17920 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_152
timestamp 1751532423
transform 1 0 18368 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_155
timestamp 1751532246
transform 1 0 18704 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_159
timestamp 1751532440
transform 1 0 19152 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_183
timestamp 1751532440
transform 1 0 21840 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_187
timestamp 1751532423
transform 1 0 22288 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_195
timestamp 1751532440
transform 1 0 23184 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_247
timestamp 1751532246
transform 1 0 29008 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_278
timestamp 1751532440
transform 1 0 32480 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_280
timestamp 1751532423
transform 1 0 32704 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_382
timestamp 1751532440
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_2
timestamp 1751532351
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_18
timestamp 1751532351
transform 1 0 3360 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_34
timestamp 1751532351
transform 1 0 5152 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_50
timestamp 1751532351
transform 1 0 6944 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_66
timestamp 1751532246
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_72
timestamp 1751532351
transform 1 0 9408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_88
timestamp 1751532440
transform 1 0 11200 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_94
timestamp 1751532351
transform 1 0 11872 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_110
timestamp 1751532351
transform 1 0 13664 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_126
timestamp 1751532246
transform 1 0 15456 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_130
timestamp 1751532440
transform 1 0 15904 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_132
timestamp 1751532423
transform 1 0 16128 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_139
timestamp 1751532423
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_142
timestamp 1751532351
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_158
timestamp 1751532351
transform 1 0 19040 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_174
timestamp 1751532246
transform 1 0 20832 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_178
timestamp 1751532423
transform 1 0 21280 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_206
timestamp 1751532440
transform 1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_212
timestamp 1751532246
transform 1 0 25088 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_250
timestamp 1751532423
transform 1 0 29344 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_282
timestamp 1751532246
transform 1 0 32928 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_286
timestamp 1751532423
transform 1 0 33376 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_321
timestamp 1751532440
transform 1 0 37296 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_352
timestamp 1751532440
transform 1 0 40768 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_354
timestamp 1751532423
transform 1 0 40992 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_382
timestamp 1751532440
transform 1 0 44128 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_2
timestamp 1751532351
transform 1 0 1568 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_18
timestamp 1751532351
transform 1 0 3360 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_34
timestamp 1751532423
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_37
timestamp 1751532351
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_53
timestamp 1751532351
transform 1 0 7280 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_69
timestamp 1751532351
transform 1 0 9072 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_85
timestamp 1751532351
transform 1 0 10864 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_101
timestamp 1751532246
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_107
timestamp 1751532351
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_150
timestamp 1751532351
transform 1 0 18144 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_166
timestamp 1751532440
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_168
timestamp 1751532423
transform 1 0 20160 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_191
timestamp 1751532246
transform 1 0 22736 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_195
timestamp 1751532440
transform 1 0 23184 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_197
timestamp 1751532423
transform 1 0 23408 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_210
timestamp 1751532423
transform 1 0 24864 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_237
timestamp 1751532312
transform 1 0 27888 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_247
timestamp 1751532312
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_255
timestamp 1751532246
transform 1 0 29904 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_259
timestamp 1751532440
transform 1 0 30352 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_275
timestamp 1751532440
transform 1 0 32144 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_277
timestamp 1751532423
transform 1 0 32368 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_314
timestamp 1751532423
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_324
timestamp 1751532440
transform 1 0 37632 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_380
timestamp 1751532440
transform 1 0 43904 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_2
timestamp 1751532351
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_18
timestamp 1751532351
transform 1 0 3360 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_34
timestamp 1751532351
transform 1 0 5152 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_50
timestamp 1751532351
transform 1 0 6944 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_66
timestamp 1751532246
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_72
timestamp 1751532351
transform 1 0 9408 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_88
timestamp 1751532351
transform 1 0 11200 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_104
timestamp 1751532246
transform 1 0 12992 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_135
timestamp 1751532246
transform 1 0 16464 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_139
timestamp 1751532423
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_142
timestamp 1751532440
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_144
timestamp 1751532423
transform 1 0 17472 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_158
timestamp 1751532246
transform 1 0 19040 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_189
timestamp 1751532440
transform 1 0 22512 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_205
timestamp 1751532246
transform 1 0 24304 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_209
timestamp 1751532423
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_212
timestamp 1751532246
transform 1 0 25088 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_222
timestamp 1751532351
transform 1 0 26208 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_238
timestamp 1751532351
transform 1 0 28000 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_254
timestamp 1751532312
transform 1 0 29792 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_262
timestamp 1751532246
transform 1 0 30688 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_282
timestamp 1751532351
transform 1 0 32928 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_298
timestamp 1751532312
transform 1 0 34720 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_306
timestamp 1751532440
transform 1 0 35616 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_308
timestamp 1751532423
transform 1 0 35840 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_313
timestamp 1751532423
transform 1 0 36400 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_2
timestamp 1751532351
transform 1 0 1568 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_18
timestamp 1751532351
transform 1 0 3360 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_34
timestamp 1751532423
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_37
timestamp 1751532351
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_53
timestamp 1751532351
transform 1 0 7280 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_69
timestamp 1751532351
transform 1 0 9072 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_85
timestamp 1751532351
transform 1 0 10864 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_101
timestamp 1751532246
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_167
timestamp 1751532440
transform 1 0 20048 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_210
timestamp 1751532423
transform 1 0 24864 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_218
timestamp 1751532246
transform 1 0 25760 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_222
timestamp 1751532423
transform 1 0 26208 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_229
timestamp 1751532423
transform 1 0 26992 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_241
timestamp 1751532246
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_247
timestamp 1751532351
transform 1 0 29008 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_263
timestamp 1751532246
transform 1 0 30800 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_267
timestamp 1751532440
transform 1 0 31248 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_293
timestamp 1751532351
transform 1 0 34160 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_309
timestamp 1751532246
transform 1 0 35952 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_313
timestamp 1751532440
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_317
timestamp 1751532246
transform 1 0 36848 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_321
timestamp 1751532440
transform 1 0 37296 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_331
timestamp 1751532423
transform 1 0 38416 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_338
timestamp 1751532440
transform 1 0 39200 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_369
timestamp 1751532440
transform 1 0 42672 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_34_373
timestamp 1751532312
transform 1 0 43120 0 1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_381
timestamp 1751532440
transform 1 0 44016 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_383
timestamp 1751532423
transform 1 0 44240 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_2
timestamp 1751532351
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_18
timestamp 1751532351
transform 1 0 3360 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_34
timestamp 1751532351
transform 1 0 5152 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_50
timestamp 1751532351
transform 1 0 6944 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_66
timestamp 1751532246
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_72
timestamp 1751532351
transform 1 0 9408 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_88
timestamp 1751532312
transform 1 0 11200 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_96
timestamp 1751532246
transform 1 0 12096 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_100
timestamp 1751532423
transform 1 0 12544 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_128
timestamp 1751532246
transform 1 0 15680 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_132
timestamp 1751532423
transform 1 0 16128 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_155
timestamp 1751532312
transform 1 0 18704 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_163
timestamp 1751532423
transform 1 0 19600 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_195
timestamp 1751532312
transform 1 0 23184 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_203
timestamp 1751532246
transform 1 0 24080 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_207
timestamp 1751532440
transform 1 0 24528 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_209
timestamp 1751532423
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_240
timestamp 1751532440
transform 1 0 28224 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_255
timestamp 1751532440
transform 1 0 29904 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_268
timestamp 1751532423
transform 1 0 31360 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_299
timestamp 1751532423
transform 1 0 34832 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_327
timestamp 1751532351
transform 1 0 37968 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_343
timestamp 1751532246
transform 1 0 39760 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_347
timestamp 1751532440
transform 1 0 40208 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_349
timestamp 1751532423
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_352
timestamp 1751532440
transform 1 0 40768 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_354
timestamp 1751532423
transform 1 0 40992 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_359
timestamp 1751532246
transform 1 0 41552 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_363
timestamp 1751532440
transform 1 0 42000 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_365
timestamp 1751532423
transform 1 0 42224 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_372
timestamp 1751532312
transform 1 0 43008 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_380
timestamp 1751532246
transform 1 0 43904 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_2
timestamp 1751532351
transform 1 0 1568 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_18
timestamp 1751532351
transform 1 0 3360 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_34
timestamp 1751532423
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_37
timestamp 1751532351
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_53
timestamp 1751532351
transform 1 0 7280 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_69
timestamp 1751532351
transform 1 0 9072 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_85
timestamp 1751532351
transform 1 0 10864 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_101
timestamp 1751532246
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_107
timestamp 1751532312
transform 1 0 13328 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_115
timestamp 1751532440
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_130
timestamp 1751532440
transform 1 0 15904 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_132
timestamp 1751532423
transform 1 0 16128 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_139
timestamp 1751532440
transform 1 0 16912 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_159
timestamp 1751532351
transform 1 0 19152 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_204
timestamp 1751532440
transform 1 0 24192 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_206
timestamp 1751532423
transform 1 0 24416 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_255
timestamp 1751532440
transform 1 0 29904 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_312
timestamp 1751532440
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_314
timestamp 1751532423
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_317
timestamp 1751532351
transform 1 0 36848 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_333
timestamp 1751532312
transform 1 0 38640 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_368
timestamp 1751532440
transform 1 0 42560 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_372
timestamp 1751532312
transform 1 0 43008 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_380
timestamp 1751532246
transform 1 0 43904 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_2
timestamp 1751532351
transform 1 0 1568 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_18
timestamp 1751532351
transform 1 0 3360 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_37_34
timestamp 1751532312
transform 1 0 5152 0 -1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_42
timestamp 1751532423
transform 1 0 6048 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_72
timestamp 1751532423
transform 1 0 9408 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_100
timestamp 1751532351
transform 1 0 12544 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_116
timestamp 1751532351
transform 1 0 14336 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_37_132
timestamp 1751532312
transform 1 0 16128 0 -1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_37_149
timestamp 1751532312
transform 1 0 18032 0 -1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_170
timestamp 1751532246
transform 1 0 20384 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_201
timestamp 1751532440
transform 1 0 23856 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_212
timestamp 1751532423
transform 1 0 25088 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_37_248
timestamp 1751532312
transform 1 0 29120 0 -1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_256
timestamp 1751532246
transform 1 0 30016 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_282
timestamp 1751532246
transform 1 0 32928 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_337
timestamp 1751532440
transform 1 0 39088 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_352
timestamp 1751532246
transform 1 0 40768 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_356
timestamp 1751532440
transform 1 0 41216 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_358
timestamp 1751532423
transform 1 0 41440 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_2
timestamp 1751532351
transform 1 0 1568 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_18
timestamp 1751532351
transform 1 0 3360 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_34
timestamp 1751532423
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_37
timestamp 1751532246
transform 1 0 5488 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_41
timestamp 1751532423
transform 1 0 5936 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_100
timestamp 1751532246
transform 1 0 12544 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_104
timestamp 1751532423
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_107
timestamp 1751532351
transform 1 0 13328 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_123
timestamp 1751532246
transform 1 0 15120 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_147
timestamp 1751532423
transform 1 0 17808 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_177
timestamp 1751532351
transform 1 0 21168 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_259
timestamp 1751532246
transform 1 0 30352 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_263
timestamp 1751532440
transform 1 0 30800 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_297
timestamp 1751532440
transform 1 0 34608 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_311
timestamp 1751532440
transform 1 0 36176 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_335
timestamp 1751532246
transform 1 0 38864 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_339
timestamp 1751532423
transform 1 0 39312 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_379
timestamp 1751532246
transform 1 0 43792 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_383
timestamp 1751532423
transform 1 0 44240 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_2
timestamp 1751532351
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_18
timestamp 1751532351
transform 1 0 3360 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_34
timestamp 1751532351
transform 1 0 5152 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_50
timestamp 1751532312
transform 1 0 6944 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_58
timestamp 1751532246
transform 1 0 7840 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_62
timestamp 1751532440
transform 1 0 8288 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_169
timestamp 1751532351
transform 1 0 20272 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_185
timestamp 1751532351
transform 1 0 22064 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_201
timestamp 1751532440
transform 1 0 23856 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_216
timestamp 1751532423
transform 1 0 25536 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_242
timestamp 1751532351
transform 1 0 28448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_258
timestamp 1751532312
transform 1 0 30240 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_266
timestamp 1751532246
transform 1 0 31136 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_270
timestamp 1751532440
transform 1 0 31584 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_279
timestamp 1751532423
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_309
timestamp 1751532440
transform 1 0 35952 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_311
timestamp 1751532423
transform 1 0 36176 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_323
timestamp 1751532440
transform 1 0 37520 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_379
timestamp 1751532246
transform 1 0 43792 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_383
timestamp 1751532423
transform 1 0 44240 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_2
timestamp 1751532351
transform 1 0 1568 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_18
timestamp 1751532351
transform 1 0 3360 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_34
timestamp 1751532423
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_37
timestamp 1751532351
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_53
timestamp 1751532351
transform 1 0 7280 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_69
timestamp 1751532312
transform 1 0 9072 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_77
timestamp 1751532423
transform 1 0 9968 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_113
timestamp 1751532246
transform 1 0 14000 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_117
timestamp 1751532423
transform 1 0 14448 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_157
timestamp 1751532351
transform 1 0 18928 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_173
timestamp 1751532440
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_183
timestamp 1751532351
transform 1 0 21840 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_199
timestamp 1751532351
transform 1 0 23632 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_215
timestamp 1751532440
transform 1 0 25424 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_235
timestamp 1751532440
transform 1 0 27664 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_239
timestamp 1751532246
transform 1 0 28112 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_243
timestamp 1751532440
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_247
timestamp 1751532351
transform 1 0 29008 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_263
timestamp 1751532440
transform 1 0 30800 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_265
timestamp 1751532423
transform 1 0 31024 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_274
timestamp 1751532423
transform 1 0 32032 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_302
timestamp 1751532440
transform 1 0 35168 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_304
timestamp 1751532423
transform 1 0 35392 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_377
timestamp 1751532246
transform 1 0 43568 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_381
timestamp 1751532440
transform 1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_383
timestamp 1751532423
transform 1 0 44240 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_2
timestamp 1751532351
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_18
timestamp 1751532351
transform 1 0 3360 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_34
timestamp 1751532351
transform 1 0 5152 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_50
timestamp 1751532351
transform 1 0 6944 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_66
timestamp 1751532246
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_86
timestamp 1751532440
transform 1 0 10976 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_102
timestamp 1751532440
transform 1 0 12768 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_104
timestamp 1751532423
transform 1 0 12992 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_139
timestamp 1751532423
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_148
timestamp 1751532351
transform 1 0 17920 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_164
timestamp 1751532440
transform 1 0 19712 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_193
timestamp 1751532440
transform 1 0 22960 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_197
timestamp 1751532312
transform 1 0 23408 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_205
timestamp 1751532246
transform 1 0 24304 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_209
timestamp 1751532423
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_212
timestamp 1751532246
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_216
timestamp 1751532440
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_218
timestamp 1751532423
transform 1 0 25760 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_255
timestamp 1751532246
transform 1 0 29904 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_259
timestamp 1751532423
transform 1 0 30352 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_266
timestamp 1751532423
transform 1 0 31136 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_289
timestamp 1751532423
transform 1 0 33712 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_307
timestamp 1751532312
transform 1 0 35728 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_315
timestamp 1751532440
transform 1 0 36624 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_328
timestamp 1751532312
transform 1 0 38080 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_336
timestamp 1751532440
transform 1 0 38976 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_379
timestamp 1751532246
transform 1 0 43792 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_383
timestamp 1751532423
transform 1 0 44240 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_2
timestamp 1751532351
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_18
timestamp 1751532351
transform 1 0 3360 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_34
timestamp 1751532423
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_37
timestamp 1751532351
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_53
timestamp 1751532351
transform 1 0 7280 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_69
timestamp 1751532351
transform 1 0 9072 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_85
timestamp 1751532246
transform 1 0 10864 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_89
timestamp 1751532440
transform 1 0 11312 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_97
timestamp 1751532312
transform 1 0 12208 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_107
timestamp 1751532351
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_123
timestamp 1751532351
transform 1 0 15120 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_139
timestamp 1751532351
transform 1 0 16912 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_155
timestamp 1751532312
transform 1 0 18704 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_163
timestamp 1751532246
transform 1 0 19600 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_167
timestamp 1751532423
transform 1 0 20048 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_198
timestamp 1751532351
transform 1 0 23520 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_214
timestamp 1751532312
transform 1 0 25312 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_222
timestamp 1751532246
transform 1 0 26208 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_226
timestamp 1751532423
transform 1 0 26656 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_241
timestamp 1751532246
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_266
timestamp 1751532440
transform 1 0 31136 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_268
timestamp 1751532423
transform 1 0 31360 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_276
timestamp 1751532246
transform 1 0 32256 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_280
timestamp 1751532423
transform 1 0 32704 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_301
timestamp 1751532312
transform 1 0 35056 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_309
timestamp 1751532246
transform 1 0 35952 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_313
timestamp 1751532440
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_342
timestamp 1751532246
transform 1 0 39648 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_346
timestamp 1751532440
transform 1 0 40096 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_2
timestamp 1751532351
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_18
timestamp 1751532351
transform 1 0 3360 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_34
timestamp 1751532351
transform 1 0 5152 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_50
timestamp 1751532351
transform 1 0 6944 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_66
timestamp 1751532246
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_72
timestamp 1751532351
transform 1 0 9408 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_88
timestamp 1751532351
transform 1 0 11200 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_104
timestamp 1751532351
transform 1 0 12992 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_120
timestamp 1751532351
transform 1 0 14784 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_136
timestamp 1751532246
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_142
timestamp 1751532351
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_158
timestamp 1751532246
transform 1 0 19040 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_162
timestamp 1751532423
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_204
timestamp 1751532246
transform 1 0 24192 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_208
timestamp 1751532440
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_43_212
timestamp 1751532312
transform 1 0 25088 0 -1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_220
timestamp 1751532246
transform 1 0 25984 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_224
timestamp 1751532440
transform 1 0 26432 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_236
timestamp 1751532440
transform 1 0 27776 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_279
timestamp 1751532423
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_302
timestamp 1751532246
transform 1 0 35168 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_332
timestamp 1751532246
transform 1 0 38528 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_336
timestamp 1751532440
transform 1 0 38976 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_352
timestamp 1751532423
transform 1 0 40768 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_380
timestamp 1751532246
transform 1 0 43904 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_2
timestamp 1751532351
transform 1 0 1568 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_18
timestamp 1751532351
transform 1 0 3360 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_34
timestamp 1751532423
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_37
timestamp 1751532351
transform 1 0 5488 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_53
timestamp 1751532351
transform 1 0 7280 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_69
timestamp 1751532351
transform 1 0 9072 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_85
timestamp 1751532351
transform 1 0 10864 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_101
timestamp 1751532246
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_107
timestamp 1751532351
transform 1 0 13328 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_123
timestamp 1751532351
transform 1 0 15120 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_139
timestamp 1751532351
transform 1 0 16912 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_44_155
timestamp 1751532312
transform 1 0 18704 0 1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_163
timestamp 1751532246
transform 1 0 19600 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_167
timestamp 1751532423
transform 1 0 20048 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_177
timestamp 1751532246
transform 1 0 21168 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_181
timestamp 1751532423
transform 1 0 21616 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_219
timestamp 1751532423
transform 1 0 25872 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_243
timestamp 1751532440
transform 1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_44_254
timestamp 1751532312
transform 1 0 29792 0 1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_262
timestamp 1751532423
transform 1 0 30688 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_276
timestamp 1751532351
transform 1 0 32256 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_44_299
timestamp 1751532312
transform 1 0 34832 0 1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_307
timestamp 1751532246
transform 1 0 35728 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_44_323
timestamp 1751532312
transform 1 0 37520 0 1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_381
timestamp 1751532440
transform 1 0 44016 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_383
timestamp 1751532423
transform 1 0 44240 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_2
timestamp 1751532351
transform 1 0 1568 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_18
timestamp 1751532351
transform 1 0 3360 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_34
timestamp 1751532351
transform 1 0 5152 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_50
timestamp 1751532351
transform 1 0 6944 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_66
timestamp 1751532246
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_72
timestamp 1751532351
transform 1 0 9408 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_88
timestamp 1751532351
transform 1 0 11200 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_104
timestamp 1751532351
transform 1 0 12992 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_120
timestamp 1751532351
transform 1 0 14784 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_136
timestamp 1751532246
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_142
timestamp 1751532351
transform 1 0 17248 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_158
timestamp 1751532246
transform 1 0 19040 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_162
timestamp 1751532440
transform 1 0 19488 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_201
timestamp 1751532440
transform 1 0 23856 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_264
timestamp 1751532440
transform 1 0 30912 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_266
timestamp 1751532423
transform 1 0 31136 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_289
timestamp 1751532312
transform 1 0 33712 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_297
timestamp 1751532423
transform 1 0 34608 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_331
timestamp 1751532312
transform 1 0 38416 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_379
timestamp 1751532246
transform 1 0 43792 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_383
timestamp 1751532423
transform 1 0 44240 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_2
timestamp 1751532351
transform 1 0 1568 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_18
timestamp 1751532351
transform 1 0 3360 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_34
timestamp 1751532423
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_37
timestamp 1751532351
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_53
timestamp 1751532351
transform 1 0 7280 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_69
timestamp 1751532351
transform 1 0 9072 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_85
timestamp 1751532351
transform 1 0 10864 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_101
timestamp 1751532246
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_107
timestamp 1751532351
transform 1 0 13328 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_123
timestamp 1751532351
transform 1 0 15120 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_139
timestamp 1751532351
transform 1 0 16912 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_155
timestamp 1751532351
transform 1 0 18704 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_171
timestamp 1751532246
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_177
timestamp 1751532246
transform 1 0 21168 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_181
timestamp 1751532423
transform 1 0 21616 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_199
timestamp 1751532246
transform 1 0 23632 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_241
timestamp 1751532440
transform 1 0 28336 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_247
timestamp 1751532312
transform 1 0 29008 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_255
timestamp 1751532440
transform 1 0 29904 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_257
timestamp 1751532423
transform 1 0 30128 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_299
timestamp 1751532246
transform 1 0 34832 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_303
timestamp 1751532423
transform 1 0 35280 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_328
timestamp 1751532312
transform 1 0 38080 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_336
timestamp 1751532440
transform 1 0 38976 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_338
timestamp 1751532423
transform 1 0 39200 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_383
timestamp 1751532423
transform 1 0 44240 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_2
timestamp 1751532351
transform 1 0 1568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_18
timestamp 1751532351
transform 1 0 3360 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_34
timestamp 1751532351
transform 1 0 5152 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_50
timestamp 1751532351
transform 1 0 6944 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_66
timestamp 1751532246
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_72
timestamp 1751532351
transform 1 0 9408 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_88
timestamp 1751532351
transform 1 0 11200 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_104
timestamp 1751532351
transform 1 0 12992 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_120
timestamp 1751532351
transform 1 0 14784 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_136
timestamp 1751532246
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_142
timestamp 1751532351
transform 1 0 17248 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_47_158
timestamp 1751532312
transform 1 0 19040 0 -1 40768
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_166
timestamp 1751532246
transform 1 0 19936 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_170
timestamp 1751532440
transform 1 0 20384 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_172
timestamp 1751532423
transform 1 0 20608 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_246
timestamp 1751532440
transform 1 0 28896 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_250
timestamp 1751532440
transform 1 0 29344 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_252
timestamp 1751532423
transform 1 0 29568 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_296
timestamp 1751532246
transform 1 0 34496 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_300
timestamp 1751532423
transform 1 0 34944 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_335
timestamp 1751532440
transform 1 0 38864 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_337
timestamp 1751532423
transform 1 0 39088 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_379
timestamp 1751532246
transform 1 0 43792 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_383
timestamp 1751532423
transform 1 0 44240 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_2
timestamp 1751532351
transform 1 0 1568 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_18
timestamp 1751532351
transform 1 0 3360 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_34
timestamp 1751532423
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_37
timestamp 1751532351
transform 1 0 5488 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_53
timestamp 1751532351
transform 1 0 7280 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_69
timestamp 1751532351
transform 1 0 9072 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_85
timestamp 1751532351
transform 1 0 10864 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_101
timestamp 1751532246
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_107
timestamp 1751532351
transform 1 0 13328 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_123
timestamp 1751532351
transform 1 0 15120 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_139
timestamp 1751532351
transform 1 0 16912 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_155
timestamp 1751532351
transform 1 0 18704 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_171
timestamp 1751532246
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_48_177
timestamp 1751532312
transform 1 0 21168 0 1 40768
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_199
timestamp 1751532351
transform 1 0 23632 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_215
timestamp 1751532423
transform 1 0 25424 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_48_230
timestamp 1751532312
transform 1 0 27104 0 1 40768
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_238
timestamp 1751532246
transform 1 0 28000 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_242
timestamp 1751532440
transform 1 0 28448 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_244
timestamp 1751532423
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_48_247
timestamp 1751532312
transform 1 0 29008 0 1 40768
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_255
timestamp 1751532440
transform 1 0 29904 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_48_291
timestamp 1751532312
transform 1 0 33936 0 1 40768
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_299
timestamp 1751532440
transform 1 0 34832 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_301
timestamp 1751532423
transform 1 0 35056 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_330
timestamp 1751532351
transform 1 0 38304 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_346
timestamp 1751532440
transform 1 0 40096 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_2
timestamp 1751532351
transform 1 0 1568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_18
timestamp 1751532351
transform 1 0 3360 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_36
timestamp 1751532351
transform 1 0 5376 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_52
timestamp 1751532351
transform 1 0 7168 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_70
timestamp 1751532351
transform 1 0 9184 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_86
timestamp 1751532351
transform 1 0 10976 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_104
timestamp 1751532351
transform 1 0 12992 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_120
timestamp 1751532351
transform 1 0 14784 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_138
timestamp 1751532351
transform 1 0 16800 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_154
timestamp 1751532351
transform 1 0 18592 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_172
timestamp 1751532351
transform 1 0 20608 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_188
timestamp 1751532351
transform 1 0 22400 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_206
timestamp 1751532351
transform 1 0 24416 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_222
timestamp 1751532351
transform 1 0 26208 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_240
timestamp 1751532351
transform 1 0 28224 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_49_256
timestamp 1751532312
transform 1 0 30016 0 -1 42336
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_264
timestamp 1751532423
transform 1 0 30912 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_284
timestamp 1751532351
transform 1 0 33152 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_300
timestamp 1751532246
transform 1 0 34944 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_304
timestamp 1751532440
transform 1 0 35392 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_308
timestamp 1751532246
transform 1 0 35840 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_312
timestamp 1751532423
transform 1 0 36288 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_320
timestamp 1751532351
transform 1 0 37184 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_336
timestamp 1751532246
transform 1 0 38976 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_342
timestamp 1751532246
transform 1 0 39648 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_346
timestamp 1751532440
transform 1 0 40096 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_348
timestamp 1751532423
transform 1 0 40320 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_49_376
timestamp 1751532312
transform 1 0 43456 0 -1 42336
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input1
timestamp 1751534193
transform -1 0 44352 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input2
timestamp 1751534193
transform -1 0 44352 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input3
timestamp 1751534193
transform -1 0 44352 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input4
timestamp 1751534193
transform -1 0 44352 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input5
timestamp 1751534193
transform -1 0 44352 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output6
timestamp 1751661108
transform 1 0 41552 0 -1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output7
timestamp 1751661108
transform -1 0 44352 0 -1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output8
timestamp 1751661108
transform -1 0 44352 0 1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output9
timestamp 1751661108
transform 1 0 41552 0 1 40768
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output10
timestamp 1751661108
transform -1 0 43232 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Left_50 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532504
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Right_0
timestamp 1751532504
transform -1 0 44576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Left_51
timestamp 1751532504
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Right_1
timestamp 1751532504
transform -1 0 44576 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Left_52
timestamp 1751532504
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Right_2
timestamp 1751532504
transform -1 0 44576 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Left_53
timestamp 1751532504
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Right_3
timestamp 1751532504
transform -1 0 44576 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Left_54
timestamp 1751532504
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Right_4
timestamp 1751532504
transform -1 0 44576 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Left_55
timestamp 1751532504
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Right_5
timestamp 1751532504
transform -1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Left_56
timestamp 1751532504
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Right_6
timestamp 1751532504
transform -1 0 44576 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Left_57
timestamp 1751532504
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Right_7
timestamp 1751532504
transform -1 0 44576 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Left_58
timestamp 1751532504
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Right_8
timestamp 1751532504
transform -1 0 44576 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Left_59
timestamp 1751532504
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Right_9
timestamp 1751532504
transform -1 0 44576 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Left_60
timestamp 1751532504
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Right_10
timestamp 1751532504
transform -1 0 44576 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Left_61
timestamp 1751532504
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Right_11
timestamp 1751532504
transform -1 0 44576 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Left_62
timestamp 1751532504
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Right_12
timestamp 1751532504
transform -1 0 44576 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Left_63
timestamp 1751532504
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Right_13
timestamp 1751532504
transform -1 0 44576 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Left_64
timestamp 1751532504
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Right_14
timestamp 1751532504
transform -1 0 44576 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Left_65
timestamp 1751532504
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Right_15
timestamp 1751532504
transform -1 0 44576 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Left_66
timestamp 1751532504
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Right_16
timestamp 1751532504
transform -1 0 44576 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Left_67
timestamp 1751532504
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Right_17
timestamp 1751532504
transform -1 0 44576 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Left_68
timestamp 1751532504
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Right_18
timestamp 1751532504
transform -1 0 44576 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Left_69
timestamp 1751532504
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Right_19
timestamp 1751532504
transform -1 0 44576 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Left_70
timestamp 1751532504
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Right_20
timestamp 1751532504
transform -1 0 44576 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Left_71
timestamp 1751532504
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Right_21
timestamp 1751532504
transform -1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Left_72
timestamp 1751532504
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Right_22
timestamp 1751532504
transform -1 0 44576 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Left_73
timestamp 1751532504
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Right_23
timestamp 1751532504
transform -1 0 44576 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Left_74
timestamp 1751532504
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Right_24
timestamp 1751532504
transform -1 0 44576 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Left_75
timestamp 1751532504
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Right_25
timestamp 1751532504
transform -1 0 44576 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Left_76
timestamp 1751532504
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Right_26
timestamp 1751532504
transform -1 0 44576 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Left_77
timestamp 1751532504
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Right_27
timestamp 1751532504
transform -1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Left_78
timestamp 1751532504
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Right_28
timestamp 1751532504
transform -1 0 44576 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Left_79
timestamp 1751532504
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Right_29
timestamp 1751532504
transform -1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Left_80
timestamp 1751532504
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Right_30
timestamp 1751532504
transform -1 0 44576 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Left_81
timestamp 1751532504
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Right_31
timestamp 1751532504
transform -1 0 44576 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Left_82
timestamp 1751532504
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Right_32
timestamp 1751532504
transform -1 0 44576 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Left_83
timestamp 1751532504
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Right_33
timestamp 1751532504
transform -1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Left_84
timestamp 1751532504
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Right_34
timestamp 1751532504
transform -1 0 44576 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Left_85
timestamp 1751532504
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Right_35
timestamp 1751532504
transform -1 0 44576 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Left_86
timestamp 1751532504
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Right_36
timestamp 1751532504
transform -1 0 44576 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Left_87
timestamp 1751532504
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Right_37
timestamp 1751532504
transform -1 0 44576 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Left_88
timestamp 1751532504
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Right_38
timestamp 1751532504
transform -1 0 44576 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Left_89
timestamp 1751532504
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Right_39
timestamp 1751532504
transform -1 0 44576 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Left_90
timestamp 1751532504
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Right_40
timestamp 1751532504
transform -1 0 44576 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Left_91
timestamp 1751532504
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Right_41
timestamp 1751532504
transform -1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Left_92
timestamp 1751532504
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Right_42
timestamp 1751532504
transform -1 0 44576 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_43_Left_93
timestamp 1751532504
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_43_Right_43
timestamp 1751532504
transform -1 0 44576 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_44_Left_94
timestamp 1751532504
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_44_Right_44
timestamp 1751532504
transform -1 0 44576 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_45_Left_95
timestamp 1751532504
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_45_Right_45
timestamp 1751532504
transform -1 0 44576 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_46_Left_96
timestamp 1751532504
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_46_Right_46
timestamp 1751532504
transform -1 0 44576 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_47_Left_97
timestamp 1751532504
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_47_Right_47
timestamp 1751532504
transform -1 0 44576 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_48_Left_98
timestamp 1751532504
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_48_Right_48
timestamp 1751532504
transform -1 0 44576 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_49_Left_99
timestamp 1751532504
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_49_Right_49
timestamp 1751532504
transform -1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_100
timestamp 1751532504
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_101
timestamp 1751532504
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_102
timestamp 1751532504
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_103
timestamp 1751532504
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_104
timestamp 1751532504
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_105
timestamp 1751532504
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_106
timestamp 1751532504
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_107
timestamp 1751532504
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_108
timestamp 1751532504
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_109
timestamp 1751532504
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_110
timestamp 1751532504
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_111
timestamp 1751532504
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_112
timestamp 1751532504
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_113
timestamp 1751532504
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_114
timestamp 1751532504
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_115
timestamp 1751532504
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_116
timestamp 1751532504
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_117
timestamp 1751532504
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_118
timestamp 1751532504
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_119
timestamp 1751532504
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_120
timestamp 1751532504
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_121
timestamp 1751532504
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_122
timestamp 1751532504
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_123
timestamp 1751532504
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_124
timestamp 1751532504
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_125
timestamp 1751532504
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_126
timestamp 1751532504
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_127
timestamp 1751532504
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_128
timestamp 1751532504
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_129
timestamp 1751532504
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_130
timestamp 1751532504
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_131
timestamp 1751532504
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_132
timestamp 1751532504
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_133
timestamp 1751532504
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_134
timestamp 1751532504
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_135
timestamp 1751532504
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_136
timestamp 1751532504
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_137
timestamp 1751532504
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_138
timestamp 1751532504
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_139
timestamp 1751532504
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_140
timestamp 1751532504
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_141
timestamp 1751532504
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_142
timestamp 1751532504
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_143
timestamp 1751532504
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_144
timestamp 1751532504
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_145
timestamp 1751532504
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_146
timestamp 1751532504
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_147
timestamp 1751532504
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_148
timestamp 1751532504
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_149
timestamp 1751532504
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_150
timestamp 1751532504
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_151
timestamp 1751532504
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_152
timestamp 1751532504
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_153
timestamp 1751532504
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_154
timestamp 1751532504
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_155
timestamp 1751532504
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_156
timestamp 1751532504
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_157
timestamp 1751532504
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_158
timestamp 1751532504
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_159
timestamp 1751532504
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_160
timestamp 1751532504
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_161
timestamp 1751532504
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_162
timestamp 1751532504
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_163
timestamp 1751532504
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_164
timestamp 1751532504
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_165
timestamp 1751532504
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_166
timestamp 1751532504
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_167
timestamp 1751532504
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_168
timestamp 1751532504
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_169
timestamp 1751532504
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_170
timestamp 1751532504
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_171
timestamp 1751532504
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_172
timestamp 1751532504
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_173
timestamp 1751532504
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_174
timestamp 1751532504
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_175
timestamp 1751532504
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_176
timestamp 1751532504
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_177
timestamp 1751532504
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_178
timestamp 1751532504
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_179
timestamp 1751532504
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_180
timestamp 1751532504
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_181
timestamp 1751532504
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_182
timestamp 1751532504
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_183
timestamp 1751532504
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_184
timestamp 1751532504
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_185
timestamp 1751532504
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_186
timestamp 1751532504
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_187
timestamp 1751532504
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_188
timestamp 1751532504
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_189
timestamp 1751532504
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_190
timestamp 1751532504
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_191
timestamp 1751532504
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_192
timestamp 1751532504
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_193
timestamp 1751532504
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_194
timestamp 1751532504
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_195
timestamp 1751532504
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_196
timestamp 1751532504
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_197
timestamp 1751532504
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_198
timestamp 1751532504
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_199
timestamp 1751532504
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_200
timestamp 1751532504
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_201
timestamp 1751532504
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_202
timestamp 1751532504
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_203
timestamp 1751532504
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_204
timestamp 1751532504
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_205
timestamp 1751532504
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_206
timestamp 1751532504
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_207
timestamp 1751532504
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_208
timestamp 1751532504
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_209
timestamp 1751532504
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_210
timestamp 1751532504
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_211
timestamp 1751532504
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_212
timestamp 1751532504
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_213
timestamp 1751532504
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_214
timestamp 1751532504
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_215
timestamp 1751532504
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_216
timestamp 1751532504
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_217
timestamp 1751532504
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_218
timestamp 1751532504
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_219
timestamp 1751532504
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_220
timestamp 1751532504
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_221
timestamp 1751532504
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_222
timestamp 1751532504
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_223
timestamp 1751532504
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_224
timestamp 1751532504
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_225
timestamp 1751532504
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_226
timestamp 1751532504
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_227
timestamp 1751532504
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_228
timestamp 1751532504
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_229
timestamp 1751532504
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_230
timestamp 1751532504
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_231
timestamp 1751532504
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_232
timestamp 1751532504
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_233
timestamp 1751532504
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_234
timestamp 1751532504
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_235
timestamp 1751532504
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_236
timestamp 1751532504
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_237
timestamp 1751532504
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_238
timestamp 1751532504
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_239
timestamp 1751532504
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_240
timestamp 1751532504
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_241
timestamp 1751532504
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_242
timestamp 1751532504
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_243
timestamp 1751532504
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_244
timestamp 1751532504
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_245
timestamp 1751532504
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_246
timestamp 1751532504
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_247
timestamp 1751532504
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_248
timestamp 1751532504
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_249
timestamp 1751532504
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_250
timestamp 1751532504
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_251
timestamp 1751532504
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_252
timestamp 1751532504
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_253
timestamp 1751532504
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_254
timestamp 1751532504
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_255
timestamp 1751532504
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_256
timestamp 1751532504
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_257
timestamp 1751532504
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_258
timestamp 1751532504
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_259
timestamp 1751532504
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_260
timestamp 1751532504
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_261
timestamp 1751532504
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_262
timestamp 1751532504
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_263
timestamp 1751532504
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_264
timestamp 1751532504
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_265
timestamp 1751532504
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_266
timestamp 1751532504
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_267
timestamp 1751532504
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_268
timestamp 1751532504
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_269
timestamp 1751532504
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_270
timestamp 1751532504
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_271
timestamp 1751532504
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_272
timestamp 1751532504
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_273
timestamp 1751532504
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_274
timestamp 1751532504
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_275
timestamp 1751532504
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_276
timestamp 1751532504
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_277
timestamp 1751532504
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_278
timestamp 1751532504
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_279
timestamp 1751532504
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_280
timestamp 1751532504
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_281
timestamp 1751532504
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_282
timestamp 1751532504
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_283
timestamp 1751532504
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_284
timestamp 1751532504
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_285
timestamp 1751532504
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_286
timestamp 1751532504
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_287
timestamp 1751532504
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_288
timestamp 1751532504
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_289
timestamp 1751532504
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_290
timestamp 1751532504
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_291
timestamp 1751532504
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_292
timestamp 1751532504
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_293
timestamp 1751532504
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_294
timestamp 1751532504
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_295
timestamp 1751532504
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_296
timestamp 1751532504
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_297
timestamp 1751532504
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_298
timestamp 1751532504
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_299
timestamp 1751532504
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_300
timestamp 1751532504
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_301
timestamp 1751532504
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_302
timestamp 1751532504
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_303
timestamp 1751532504
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_304
timestamp 1751532504
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_305
timestamp 1751532504
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_306
timestamp 1751532504
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_307
timestamp 1751532504
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_308
timestamp 1751532504
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_309
timestamp 1751532504
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_310
timestamp 1751532504
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_311
timestamp 1751532504
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_312
timestamp 1751532504
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_313
timestamp 1751532504
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_314
timestamp 1751532504
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_315
timestamp 1751532504
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_316
timestamp 1751532504
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_317
timestamp 1751532504
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_318
timestamp 1751532504
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_319
timestamp 1751532504
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_320
timestamp 1751532504
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_321
timestamp 1751532504
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_322
timestamp 1751532504
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_323
timestamp 1751532504
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_324
timestamp 1751532504
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_325
timestamp 1751532504
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_326
timestamp 1751532504
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_327
timestamp 1751532504
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_328
timestamp 1751532504
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_329
timestamp 1751532504
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_330
timestamp 1751532504
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_331
timestamp 1751532504
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_332
timestamp 1751532504
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_333
timestamp 1751532504
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_334
timestamp 1751532504
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_335
timestamp 1751532504
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_336
timestamp 1751532504
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_337
timestamp 1751532504
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_338
timestamp 1751532504
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_339
timestamp 1751532504
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_340
timestamp 1751532504
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_341
timestamp 1751532504
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_342
timestamp 1751532504
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_343
timestamp 1751532504
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_344
timestamp 1751532504
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_345
timestamp 1751532504
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_346
timestamp 1751532504
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_347
timestamp 1751532504
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_348
timestamp 1751532504
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_349
timestamp 1751532504
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_350
timestamp 1751532504
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_351
timestamp 1751532504
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_352
timestamp 1751532504
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_353
timestamp 1751532504
transform 1 0 12768 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_354
timestamp 1751532504
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_355
timestamp 1751532504
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_356
timestamp 1751532504
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_357
timestamp 1751532504
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_358
timestamp 1751532504
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_359
timestamp 1751532504
transform 1 0 35616 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_360
timestamp 1751532504
transform 1 0 39424 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_361
timestamp 1751532504
transform 1 0 43232 0 -1 42336
box -86 -86 310 870
<< labels >>
flabel metal3 s 45200 2688 46000 2800 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 45200 9408 46000 9520 0 FreeSans 448 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal3 s 45200 12768 46000 12880 0 FreeSans 448 0 0 0 io_in[1]
port 2 nsew signal input
flabel metal3 s 45200 16128 46000 16240 0 FreeSans 448 0 0 0 io_in[2]
port 3 nsew signal input
flabel metal3 s 45200 19488 46000 19600 0 FreeSans 448 0 0 0 io_in[3]
port 4 nsew signal input
flabel metal3 s 45200 22848 46000 22960 0 FreeSans 448 0 0 0 io_in[4]
port 5 nsew signal input
flabel metal3 s 45200 26208 46000 26320 0 FreeSans 448 0 0 0 io_in[5]
port 6 nsew signal input
flabel metal3 s 45200 29568 46000 29680 0 FreeSans 448 0 0 0 io_out[0]
port 7 nsew signal output
flabel metal3 s 45200 32928 46000 33040 0 FreeSans 448 0 0 0 io_out[1]
port 8 nsew signal output
flabel metal3 s 45200 36288 46000 36400 0 FreeSans 448 0 0 0 io_out[2]
port 9 nsew signal output
flabel metal3 s 45200 39648 46000 39760 0 FreeSans 448 0 0 0 io_out[3]
port 10 nsew signal output
flabel metal3 s 45200 43008 46000 43120 0 FreeSans 448 0 0 0 io_out[4]
port 11 nsew signal output
flabel metal3 s 45200 6048 46000 6160 0 FreeSans 448 0 0 0 rst_n
port 12 nsew signal input
flabel metal4 s 4448 3076 4768 42396 0 FreeSans 1280 90 0 0 vdd
port 13 nsew power bidirectional
flabel metal4 s 35168 3076 35488 42396 0 FreeSans 1280 90 0 0 vdd
port 13 nsew power bidirectional
flabel metal4 s 19808 3076 20128 42396 0 FreeSans 1280 90 0 0 vss
port 14 nsew ground bidirectional
rlabel metal1 22960 41552 22960 41552 0 vdd
rlabel metal1 22960 42336 22960 42336 0 vss
rlabel metal2 24080 27944 24080 27944 0 CIRCUIT_2223.CLK
rlabel metal2 26488 18648 26488 18648 0 CIRCUIT_2223.GATES_1.input1\[0\]
rlabel metal2 25536 16184 25536 16184 0 CIRCUIT_2223.GATES_1.input1\[1\]
rlabel metal2 30240 15288 30240 15288 0 CIRCUIT_2223.GATES_1.input1\[2\]
rlabel metal3 28112 16072 28112 16072 0 CIRCUIT_2223.GATES_1.input1\[3\]
rlabel metal2 30856 28504 30856 28504 0 CIRCUIT_2223.GATES_2.input2
rlabel metal3 27496 23800 27496 23800 0 CIRCUIT_2223.GATES_3.input2
rlabel via2 25480 31738 25480 31738 0 CIRCUIT_2223.GATES_4.input1\[0\]
rlabel metal2 24248 31864 24248 31864 0 CIRCUIT_2223.GATES_4.input1\[1\]
rlabel metal3 24584 30184 24584 30184 0 CIRCUIT_2223.GATES_4.input1\[2\]
rlabel via1 27440 30166 27440 30166 0 CIRCUIT_2223.GATES_4.input1\[3\]
rlabel metal2 28504 29456 28504 29456 0 CIRCUIT_2223.GATES_5.input2
rlabel metal2 14056 10864 14056 10864 0 CIRCUIT_2223.MEMORY_18.s_currentState
rlabel metal2 10360 25312 10360 25312 0 CIRCUIT_2223.MEMORY_19.s_currentState
rlabel metal3 11144 27832 11144 27832 0 CIRCUIT_2223.MEMORY_20.s_currentState
rlabel metal2 13384 25424 13384 25424 0 CIRCUIT_2223.MEMORY_21.s_currentState
rlabel metal2 16632 27160 16632 27160 0 CIRCUIT_2223.MEMORY_22.s_currentState
rlabel metal2 19992 24864 19992 24864 0 CIRCUIT_2223.MEMORY_23.s_currentState
rlabel metal2 23912 26152 23912 26152 0 CIRCUIT_2223.MEMORY_24.s_currentState
rlabel metal2 15736 24072 15736 24072 0 CIRCUIT_2223.MEMORY_25.s_currentState
rlabel metal2 17024 25592 17024 25592 0 CIRCUIT_2223.MEMORY_26.s_currentState
rlabel metal2 42448 30184 42448 30184 0 CIRCUIT_2223.MEMORY_28.s_currentState
rlabel metal3 42784 31864 42784 31864 0 CIRCUIT_2223.MEMORY_29.s_currentState
rlabel metal2 25592 29120 25592 29120 0 CIRCUIT_2223.s_logisimNet48
rlabel metal2 9912 33656 9912 33656 0 CIRCUIT_2223.tone_generator_1.GATES_1.result
rlabel metal3 10024 32536 10024 32536 0 CIRCUIT_2223.tone_generator_1.GATES_2.result
rlabel metal2 11816 34328 11816 34328 0 CIRCUIT_2223.tone_generator_1.GATES_3.result
rlabel metal2 13776 34216 13776 34216 0 CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState
rlabel metal2 16016 35672 16016 35672 0 CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState
rlabel metal2 16408 33656 16408 33656 0 CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState
rlabel metal3 16520 33320 16520 33320 0 CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState
rlabel metal2 19992 33544 19992 33544 0 CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState
rlabel metal2 15400 31192 15400 31192 0 CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState
rlabel metal2 16240 29512 16240 29512 0 CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState
rlabel metal2 17864 30800 17864 30800 0 CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState
rlabel metal2 17808 28728 17808 28728 0 CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState
rlabel metal2 19656 31416 19656 31416 0 CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState
rlabel metal2 8344 32368 8344 32368 0 CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState
rlabel metal2 6440 32984 6440 32984 0 CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState
rlabel metal2 8848 33432 8848 33432 0 CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState
rlabel metal3 10808 33432 10808 33432 0 CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState
rlabel metal2 12264 32760 12264 32760 0 CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState
rlabel metal2 10360 35168 10360 35168 0 CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState
rlabel metal3 34813 5880 34813 5880 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2
rlabel metal2 32424 11592 32424 11592 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2
rlabel metal2 35784 13384 35784 13384 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2
rlabel metal2 35728 14364 35728 14364 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2
rlabel metal2 38715 7812 38715 7812 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2
rlabel metal2 39928 15456 39928 15456 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2
rlabel metal2 41664 13468 41664 13468 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2
rlabel metal2 41748 15288 41748 15288 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2
rlabel metal2 21896 25116 21896 25116 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result
rlabel metal2 43288 12320 43288 12320 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2
rlabel metal2 36120 4480 36120 4480 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2
rlabel metal2 39592 5712 39592 5712 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2
rlabel metal3 42224 6552 42224 6552 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState
rlabel metal3 42672 4200 42672 4200 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState
rlabel metal3 39760 4312 39760 4312 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState
rlabel metal2 40936 5992 40936 5992 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState
rlabel metal2 31752 10864 31752 10864 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState
rlabel metal2 34664 10640 34664 10640 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState
rlabel metal3 35896 12936 35896 12936 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState
rlabel metal2 39592 7672 39592 7672 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState
rlabel metal2 39592 9856 39592 9856 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState
rlabel metal3 41552 9688 41552 9688 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState
rlabel metal2 43848 8802 43848 8802 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState
rlabel metal2 21672 29792 21672 29792 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d
rlabel metal2 20328 29848 20328 29848 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState
rlabel metal2 29932 7504 29932 7504 0 CIRCUIT_2223.tone_generator_2_1.GATES_10.input2
rlabel metal2 26040 11592 26040 11592 0 CIRCUIT_2223.tone_generator_2_1.GATES_11.input2
rlabel metal2 24584 11928 24584 11928 0 CIRCUIT_2223.tone_generator_2_1.GATES_12.input2
rlabel metal2 25368 11144 25368 11144 0 CIRCUIT_2223.tone_generator_2_1.GATES_13.input2
rlabel metal2 21336 13888 21336 13888 0 CIRCUIT_2223.tone_generator_2_1.GATES_14.input2
rlabel metal2 24360 5152 24360 5152 0 CIRCUIT_2223.tone_generator_2_1.GATES_15.input2
rlabel metal2 26059 6524 26059 6524 0 CIRCUIT_2223.tone_generator_2_1.GATES_16.input2
rlabel metal3 25638 5880 25638 5880 0 CIRCUIT_2223.tone_generator_2_1.GATES_17.input2
rlabel metal3 24136 21504 24136 21504 0 CIRCUIT_2223.tone_generator_2_1.GATES_27.result
rlabel metal2 23632 15176 23632 15176 0 CIRCUIT_2223.tone_generator_2_1.GATES_7.input2
rlabel metal2 29624 5544 29624 5544 0 CIRCUIT_2223.tone_generator_2_1.GATES_8.input2
rlabel metal3 28914 6664 28914 6664 0 CIRCUIT_2223.tone_generator_2_1.GATES_9.input2
rlabel metal3 15848 5880 15848 5880 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState
rlabel metal2 18480 6552 18480 6552 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState
rlabel metal2 19208 7392 19208 7392 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState
rlabel metal2 21560 8568 21560 8568 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState
rlabel metal2 17864 10080 17864 10080 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState
rlabel metal3 19544 11480 19544 11480 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState
rlabel metal2 19320 10080 19320 10080 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState
rlabel metal2 18984 6272 18984 6272 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState
rlabel metal3 21560 5152 21560 5152 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState
rlabel metal2 22904 4424 22904 4424 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState
rlabel metal2 20664 5600 20664 5600 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState
rlabel metal2 28336 22988 28336 22988 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d
rlabel metal2 28168 23352 28168 23352 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState
rlabel metal3 36904 18424 36904 18424 0 CIRCUIT_2223.tone_generator_2_2.GATES_10.input2
rlabel metal2 35616 17948 35616 17948 0 CIRCUIT_2223.tone_generator_2_2.GATES_11.input2
rlabel metal2 37184 19292 37184 19292 0 CIRCUIT_2223.tone_generator_2_2.GATES_12.input2
rlabel metal2 39144 22960 39144 22960 0 CIRCUIT_2223.tone_generator_2_2.GATES_13.input2
rlabel metal2 42336 22232 42336 22232 0 CIRCUIT_2223.tone_generator_2_2.GATES_14.input2
rlabel metal2 40544 19292 40544 19292 0 CIRCUIT_2223.tone_generator_2_2.GATES_15.input2
rlabel metal2 43568 19320 43568 19320 0 CIRCUIT_2223.tone_generator_2_2.GATES_16.input2
rlabel metal2 43512 18536 43512 18536 0 CIRCUIT_2223.tone_generator_2_2.GATES_17.input2
rlabel metal3 30016 26040 30016 26040 0 CIRCUIT_2223.tone_generator_2_2.GATES_27.result
rlabel metal2 43848 21840 43848 21840 0 CIRCUIT_2223.tone_generator_2_2.GATES_7.input2
rlabel metal2 35672 21000 35672 21000 0 CIRCUIT_2223.tone_generator_2_2.GATES_8.input2
rlabel metal3 35504 20888 35504 20888 0 CIRCUIT_2223.tone_generator_2_2.GATES_9.input2
rlabel metal3 38360 24696 38360 24696 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState
rlabel metal2 33824 23128 33824 23128 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState
rlabel metal3 32928 23128 32928 23128 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState
rlabel metal3 35952 23912 35952 23912 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState
rlabel metal2 32592 26264 32592 26264 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState
rlabel metal2 36960 26712 36960 26712 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState
rlabel metal3 37576 26376 37576 26376 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState
rlabel metal2 40656 28504 40656 28504 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState
rlabel metal2 43736 28112 43736 28112 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState
rlabel metal2 44016 27720 44016 27720 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState
rlabel metal2 40432 26264 40432 26264 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState
rlabel metal3 29988 27160 29988 27160 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d
rlabel metal2 31640 27888 31640 27888 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState
rlabel metal2 22176 21028 22176 21028 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2
rlabel metal2 15344 20664 15344 20664 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2
rlabel metal3 17080 21392 17080 21392 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2
rlabel metal2 18256 18116 18256 18116 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2
rlabel metal2 18256 17108 18256 17108 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2
rlabel metal2 14036 13664 14036 13664 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2
rlabel metal2 14504 13216 14504 13216 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2
rlabel metal2 18256 15428 18256 15428 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2
rlabel metal2 21112 23212 21112 23212 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result
rlabel metal2 14372 14420 14372 14420 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2
rlabel metal2 22456 17192 22456 17192 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2
rlabel metal2 21784 19656 21784 19656 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2
rlabel metal3 13496 14672 13496 14672 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState
rlabel metal3 9408 17752 9408 17752 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState
rlabel metal2 12600 22288 12600 22288 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState
rlabel metal2 12824 22792 12824 22792 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState
rlabel metal2 8792 19656 8792 19656 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState
rlabel metal2 9688 22064 9688 22064 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState
rlabel metal2 9128 16912 9128 16912 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState
rlabel metal3 10472 16856 10472 16856 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState
rlabel metal2 7560 14224 7560 14224 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState
rlabel metal2 7784 14448 7784 14448 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState
rlabel metal2 8568 13664 8568 13664 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState
rlabel metal2 22064 24024 22064 24024 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d
rlabel metal3 23464 26264 23464 26264 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState
rlabel metal2 28896 32396 28896 32396 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock
rlabel metal3 28812 31864 28812 31864 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d
rlabel metal3 26460 31640 26460 31640 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState
rlabel metal2 24248 33544 24248 33544 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock
rlabel metal3 28728 32536 28728 32536 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState
rlabel metal2 25480 33768 25480 33768 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState
rlabel metal3 43428 9016 43428 9016 0 _0000_
rlabel metal3 40068 9800 40068 9800 0 _0001_
rlabel metal2 36988 8008 36988 8008 0 _0002_
rlabel metal2 35448 11088 35448 11088 0 _0003_
rlabel metal2 33544 9296 33544 9296 0 _0004_
rlabel metal2 31752 9856 31752 9856 0 _0005_
rlabel metal2 42616 3584 42616 3584 0 _0006_
rlabel metal2 39928 5152 39928 5152 0 _0007_
rlabel metal2 44072 5376 44072 5376 0 _0008_
rlabel metal2 44128 6664 44128 6664 0 _0009_
rlabel metal2 7896 15792 7896 15792 0 _0010_
rlabel metal2 8260 17080 8260 17080 0 _0011_
rlabel metal2 8400 19124 8400 19124 0 _0012_
rlabel metal2 10136 22792 10136 22792 0 _0013_
rlabel metal3 8876 21560 8876 21560 0 _0014_
rlabel metal2 9744 18732 9744 18732 0 _0015_
rlabel metal2 9408 16856 9408 16856 0 _0016_
rlabel metal2 12376 14392 12376 14392 0 _0017_
rlabel metal2 7392 13216 7392 13216 0 _0018_
rlabel metal2 28728 31640 28728 31640 0 _0019_
rlabel metal2 25564 32536 25564 32536 0 _0020_
rlabel metal2 23324 33320 23324 33320 0 _0021_
rlabel metal2 8064 13048 8064 13048 0 _0022_
rlabel metal2 17864 5376 17864 5376 0 _0023_
rlabel metal2 16352 6384 16352 6384 0 _0024_
rlabel metal2 16800 7952 16800 7952 0 _0025_
rlabel metal3 17612 9016 17612 9016 0 _0026_
rlabel metal2 16828 9240 16828 9240 0 _0027_
rlabel metal2 22148 10584 22148 10584 0 _0028_
rlabel metal2 19096 7896 19096 7896 0 _0029_
rlabel metal2 19656 5712 19656 5712 0 _0030_
rlabel metal2 22232 4592 22232 4592 0 _0031_
rlabel metal2 17976 4816 17976 4816 0 _0032_
rlabel metal2 40376 27832 40376 27832 0 _0033_
rlabel metal2 37240 28168 37240 28168 0 _0034_
rlabel metal3 33180 23352 33180 23352 0 _0035_
rlabel metal2 33152 23632 33152 23632 0 _0036_
rlabel metal2 33236 26488 33236 26488 0 _0037_
rlabel metal2 35112 26544 35112 26544 0 _0038_
rlabel metal3 37324 28616 37324 28616 0 _0039_
rlabel metal2 40908 27272 40908 27272 0 _0040_
rlabel metal2 41160 28728 41160 28728 0 _0041_
rlabel metal2 40740 22904 40740 22904 0 _0042_
rlabel metal2 38136 30968 38136 30968 0 _0043_
rlabel metal2 39704 30016 39704 30016 0 _0044_
rlabel metal2 14392 25536 14392 25536 0 _0045_
rlabel metal2 14056 24976 14056 24976 0 _0046_
rlabel metal3 17080 24696 17080 24696 0 _0047_
rlabel metal2 13552 25200 13552 25200 0 _0048_
rlabel metal2 11340 27608 11340 27608 0 _0049_
rlabel metal2 9940 27048 9940 27048 0 _0050_
rlabel metal2 11116 24136 11116 24136 0 _0051_
rlabel metal2 17472 25760 17472 25760 0 _0052_
rlabel via2 39592 39578 39592 39578 0 _0053_
rlabel metal2 36176 38808 36176 38808 0 _0054_
rlabel metal2 35896 40880 35896 40880 0 _0055_
rlabel metal2 30520 41048 30520 41048 0 _0056_
rlabel metal3 32144 41272 32144 41272 0 _0057_
rlabel via1 39816 39578 39816 39578 0 _0058_
rlabel metal3 40880 40264 40880 40264 0 _0059_
rlabel metal3 40432 39704 40432 39704 0 _0060_
rlabel metal2 42952 38472 42952 38472 0 _0061_
rlabel metal3 42392 37240 42392 37240 0 _0062_
rlabel metal3 40544 35560 40544 35560 0 _0063_
rlabel metal3 39564 32760 39564 32760 0 _0064_
rlabel metal2 20552 17136 20552 17136 0 _0065_
rlabel metal2 19880 18480 19880 18480 0 _0066_
rlabel metal2 19992 20104 19992 20104 0 _0067_
rlabel metal2 24920 38892 24920 38892 0 _0068_
rlabel metal2 26488 40992 26488 40992 0 _0069_
rlabel metal3 25200 40264 25200 40264 0 _0070_
rlabel metal2 23016 39032 23016 39032 0 _0071_
rlabel metal2 20552 38668 20552 38668 0 _0072_
rlabel metal2 20440 36848 20440 36848 0 _0073_
rlabel metal2 21448 35224 21448 35224 0 _0074_
rlabel metal2 22232 28112 22232 28112 0 _0075_
rlabel metal2 29960 36736 29960 36736 0 _0076_
rlabel metal2 31080 39312 31080 39312 0 _0077_
rlabel metal3 28560 35672 28560 35672 0 _0078_
rlabel metal2 39032 34272 39032 34272 0 _0079_
rlabel metal2 35728 30968 35728 30968 0 _0080_
rlabel metal2 35840 32536 35840 32536 0 _0081_
rlabel metal2 33096 34552 33096 34552 0 _0082_
rlabel metal3 40488 35000 40488 35000 0 _0083_
rlabel metal3 25144 18424 25144 18424 0 _0084_
rlabel metal3 23408 16184 23408 16184 0 _0085_
rlabel metal3 28952 13160 28952 13160 0 _0086_
rlabel metal3 29512 15176 29512 15176 0 _0087_
rlabel metal2 14840 34384 14840 34384 0 _0088_
rlabel metal3 18032 34888 18032 34888 0 _0089_
rlabel metal2 18088 34776 18088 34776 0 _0090_
rlabel metal2 13496 31248 13496 31248 0 _0091_
rlabel metal2 14280 29680 14280 29680 0 _0092_
rlabel metal2 16520 28224 16520 28224 0 _0093_
rlabel metal2 15960 30128 15960 30128 0 _0094_
rlabel metal2 17920 30296 17920 30296 0 _0095_
rlabel metal2 38024 14952 38024 14952 0 _0096_
rlabel metal3 42336 15176 42336 15176 0 _0097_
rlabel metal3 42840 12152 42840 12152 0 _0098_
rlabel metal3 40768 13048 40768 13048 0 _0099_
rlabel metal2 30520 12824 30520 12824 0 _0100_
rlabel metal3 35168 12376 35168 12376 0 _0101_
rlabel metal3 36232 15064 36232 15064 0 _0102_
rlabel metal2 39032 13272 39032 13272 0 _0103_
rlabel metal3 43344 7336 43344 7336 0 _0104_
rlabel metal2 39928 7896 39928 7896 0 _0105_
rlabel metal2 37352 6188 37352 6188 0 _0106_
rlabel metal2 36008 8232 36008 8232 0 _0107_
rlabel metal3 35112 11480 35112 11480 0 _0108_
rlabel metal2 32592 9912 32592 9912 0 _0109_
rlabel metal2 29848 11200 29848 11200 0 _0110_
rlabel metal2 41832 4704 41832 4704 0 _0111_
rlabel metal2 38808 4368 38808 4368 0 _0112_
rlabel metal2 43288 3920 43288 3920 0 _0113_
rlabel metal2 43288 5992 43288 5992 0 _0114_
rlabel metal2 20160 32760 20160 32760 0 _0115_
rlabel metal2 32088 21056 32088 21056 0 _0116_
rlabel metal2 33320 21504 33320 21504 0 _0117_
rlabel metal2 34328 18704 34328 18704 0 _0118_
rlabel metal2 8232 15624 8232 15624 0 _0119_
rlabel metal2 8344 18144 8344 18144 0 _0120_
rlabel metal2 12264 20720 12264 20720 0 _0121_
rlabel metal2 10920 22568 10920 22568 0 _0122_
rlabel metal2 8344 20328 8344 20328 0 _0123_
rlabel metal2 10248 21672 10248 21672 0 _0124_
rlabel metal2 10136 18536 10136 18536 0 _0125_
rlabel metal2 9016 15512 9016 15512 0 _0126_
rlabel metal3 10192 14616 10192 14616 0 _0127_
rlabel metal2 8232 12880 8232 12880 0 _0128_
rlabel metal2 9800 13160 9800 13160 0 _0129_
rlabel metal2 17640 20496 17640 20496 0 _0130_
rlabel metal2 16240 21560 16240 21560 0 _0131_
rlabel metal2 16240 16184 16240 16184 0 _0132_
rlabel metal2 16632 17360 16632 17360 0 _0133_
rlabel metal3 16912 12152 16912 12152 0 _0134_
rlabel metal2 16408 13272 16408 13272 0 _0135_
rlabel metal2 16632 14840 16632 14840 0 _0136_
rlabel metal3 18480 15176 18480 15176 0 _0137_
rlabel metal2 34552 3752 34552 3752 0 _0138_
rlabel metal2 36736 3752 36736 3752 0 _0139_
rlabel metal3 35056 5096 35056 5096 0 _0140_
rlabel metal2 17080 5712 17080 5712 0 _0141_
rlabel metal3 17024 5768 17024 5768 0 _0142_
rlabel metal2 17304 8456 17304 8456 0 _0143_
rlabel metal2 18760 7868 18760 7868 0 _0144_
rlabel metal3 16128 10472 16128 10472 0 _0145_
rlabel metal2 18760 11760 18760 11760 0 _0146_
rlabel metal2 21224 9576 21224 9576 0 _0147_
rlabel metal2 19432 6160 19432 6160 0 _0148_
rlabel metal3 19544 5768 19544 5768 0 _0149_
rlabel metal3 21952 4200 21952 4200 0 _0150_
rlabel metal2 18088 4648 18088 4648 0 _0151_
rlabel metal2 27944 11704 27944 11704 0 _0152_
rlabel metal3 23576 10808 23576 10808 0 _0153_
rlabel metal3 27888 10472 27888 10472 0 _0154_
rlabel metal3 23856 13608 23856 13608 0 _0155_
rlabel metal2 26824 4704 26824 4704 0 _0156_
rlabel metal2 22568 5432 22568 5432 0 _0157_
rlabel metal2 27048 5208 27048 5208 0 _0158_
rlabel metal2 22120 15064 22120 15064 0 _0159_
rlabel metal2 31528 6216 31528 6216 0 _0160_
rlabel metal2 31304 6160 31304 6160 0 _0161_
rlabel metal3 30520 8344 30520 8344 0 _0162_
rlabel metal2 37576 28560 37576 28560 0 _0163_
rlabel metal2 35896 28448 35896 28448 0 _0164_
rlabel metal2 33544 25704 33544 25704 0 _0165_
rlabel metal3 34832 24024 34832 24024 0 _0166_
rlabel metal3 31416 25592 31416 25592 0 _0167_
rlabel metal2 34440 27608 34440 27608 0 _0168_
rlabel metal3 36456 27496 36456 27496 0 _0169_
rlabel metal3 40040 28728 40040 28728 0 _0170_
rlabel metal3 43708 26936 43708 26936 0 _0171_
rlabel metal2 42000 27272 42000 27272 0 _0172_
rlabel metal2 41720 27048 41720 27048 0 _0173_
rlabel metal2 38696 18088 38696 18088 0 _0174_
rlabel metal2 38584 19656 38584 19656 0 _0175_
rlabel metal2 39760 21560 39760 21560 0 _0176_
rlabel metal2 40264 20160 40264 20160 0 _0177_
rlabel metal2 40208 17752 40208 17752 0 _0178_
rlabel metal3 42336 17080 42336 17080 0 _0179_
rlabel metal2 41608 19096 41608 19096 0 _0180_
rlabel metal2 42224 21000 42224 21000 0 _0181_
rlabel metal2 15176 25256 15176 25256 0 _0182_
rlabel metal2 14840 24304 14840 24304 0 _0183_
rlabel metal3 21280 25592 21280 25592 0 _0184_
rlabel metal2 18088 24304 18088 24304 0 _0185_
rlabel metal3 15120 27160 15120 27160 0 _0186_
rlabel metal2 11592 25984 11592 25984 0 _0187_
rlabel metal2 10752 27048 10752 27048 0 _0188_
rlabel metal2 11480 24640 11480 24640 0 _0189_
rlabel metal2 18256 25592 18256 25592 0 _0190_
rlabel metal2 28112 25704 28112 25704 0 _0191_
rlabel metal3 24920 24024 24920 24024 0 _0192_
rlabel metal2 26376 28336 26376 28336 0 _0193_
rlabel metal2 25536 27160 25536 27160 0 _0194_
rlabel metal3 22064 26488 22064 26488 0 _0195_
rlabel metal2 20104 26376 20104 26376 0 _0196_
rlabel metal3 18312 26264 18312 26264 0 _0197_
rlabel metal2 16184 23912 16184 23912 0 _0198_
rlabel metal3 30912 22344 30912 22344 0 _0199_
rlabel metal3 21224 22344 21224 22344 0 _0200_
rlabel metal2 30184 16968 30184 16968 0 _0201_
rlabel metal2 29848 16940 29848 16940 0 _0202_
rlabel metal2 29960 16912 29960 16912 0 _0203_
rlabel metal2 29512 15994 29512 15994 0 _0204_
rlabel metal3 30184 19992 30184 19992 0 _0205_
rlabel metal2 27608 17248 27608 17248 0 _0206_
rlabel metal3 28896 18312 28896 18312 0 _0207_
rlabel metal2 29512 20468 29512 20468 0 _0208_
rlabel metal2 21672 25340 21672 25340 0 _0209_
rlabel metal2 22680 23072 22680 23072 0 _0210_
rlabel metal2 41944 22848 41944 22848 0 _0211_
rlabel metal2 40936 24620 40936 24620 0 _0212_
rlabel metal2 40712 24472 40712 24472 0 _0213_
rlabel metal2 40376 24808 40376 24808 0 _0214_
rlabel metal2 38248 23968 38248 23968 0 _0215_
rlabel metal2 38584 22624 38584 22624 0 _0216_
rlabel metal2 38864 22316 38864 22316 0 _0217_
rlabel metal2 39256 22848 39256 22848 0 _0218_
rlabel metal2 38248 23072 38248 23072 0 _0219_
rlabel metal2 37800 23128 37800 23128 0 _0220_
rlabel metal3 37296 22568 37296 22568 0 _0221_
rlabel metal2 38696 22904 38696 22904 0 _0222_
rlabel metal3 40992 22568 40992 22568 0 _0223_
rlabel metal2 37576 23688 37576 23688 0 _0224_
rlabel metal2 30968 26208 30968 26208 0 _0225_
rlabel metal2 29960 21840 29960 21840 0 _0226_
rlabel metal2 29316 21672 29316 21672 0 _0227_
rlabel metal2 31080 23632 31080 23632 0 _0228_
rlabel metal2 36176 25704 36176 25704 0 _0229_
rlabel metal3 39984 28056 39984 28056 0 _0230_
rlabel metal2 32424 23744 32424 23744 0 _0231_
rlabel metal2 27496 16128 27496 16128 0 _0232_
rlabel metal2 25480 17752 25480 17752 0 _0233_
rlabel metal2 27832 19488 27832 19488 0 _0234_
rlabel metal2 26600 17080 26600 17080 0 _0235_
rlabel metal2 27384 20384 27384 20384 0 _0236_
rlabel metal2 25256 8400 25256 8400 0 _0237_
rlabel metal2 23464 8736 23464 8736 0 _0238_
rlabel metal2 23912 11032 23912 11032 0 _0239_
rlabel metal2 24696 10864 24696 10864 0 _0240_
rlabel metal2 24136 6608 24136 6608 0 _0241_
rlabel via2 24472 6650 24472 6650 0 _0242_
rlabel metal2 24584 6328 24584 6328 0 _0243_
rlabel metal2 25144 7952 25144 7952 0 _0244_
rlabel metal2 24248 7504 24248 7504 0 _0245_
rlabel metal2 26488 6104 26488 6104 0 _0246_
rlabel metal2 28392 6944 28392 6944 0 _0247_
rlabel metal2 27496 7448 27496 7448 0 _0248_
rlabel metal2 28840 6272 28840 6272 0 _0249_
rlabel metal2 25928 8456 25928 8456 0 _0250_
rlabel metal2 25704 17556 25704 17556 0 _0251_
rlabel metal2 24696 21056 24696 21056 0 _0252_
rlabel metal3 22829 21000 22829 21000 0 _0253_
rlabel metal2 19488 17416 19488 17416 0 _0254_
rlabel via2 21336 9786 21336 9786 0 _0255_
rlabel metal2 21112 3738 21112 3738 0 _0256_
rlabel metal2 20440 10010 20440 10010 0 _0257_
rlabel metal2 14616 18144 14616 18144 0 _0258_
rlabel metal2 14952 20356 14952 20356 0 _0259_
rlabel metal2 15288 19292 15288 19292 0 _0260_
rlabel metal2 15008 18312 15008 18312 0 _0261_
rlabel metal2 13776 12264 13776 12264 0 _0262_
rlabel metal2 14616 14840 14616 14840 0 _0263_
rlabel metal2 13944 15456 13944 15456 0 _0264_
rlabel metal2 14224 13832 14224 13832 0 _0265_
rlabel metal2 15400 18508 15400 18508 0 _0266_
rlabel metal2 12712 18536 12712 18536 0 _0267_
rlabel metal2 13832 19124 13832 19124 0 _0268_
rlabel metal2 14224 19208 14224 19208 0 _0269_
rlabel metal2 12824 16688 12824 16688 0 _0270_
rlabel metal2 15736 19264 15736 19264 0 _0271_
rlabel metal2 15624 20020 15624 20020 0 _0272_
rlabel metal2 27944 18508 27944 18508 0 _0273_
rlabel metal2 22232 17584 22232 17584 0 _0274_
rlabel metal2 24920 16968 24920 16968 0 _0275_
rlabel metal2 26824 18480 26824 18480 0 _0276_
rlabel metal2 22232 18200 22232 18200 0 _0277_
rlabel metal2 26152 16968 26152 16968 0 _0278_
rlabel metal2 21560 17360 21560 17360 0 _0279_
rlabel metal2 20888 23086 20888 23086 0 _0280_
rlabel metal2 19899 22568 19899 22568 0 _0281_
rlabel metal2 19656 22680 19656 22680 0 _0282_
rlabel metal2 8904 19893 8904 19893 0 _0283_
rlabel metal2 10248 15469 10248 15469 0 _0284_
rlabel metal2 14728 20229 14728 20229 0 _0285_
rlabel metal2 35448 6328 35448 6328 0 _0286_
rlabel metal2 37016 4928 37016 4928 0 _0287_
rlabel metal2 37688 6608 37688 6608 0 _0288_
rlabel metal2 37128 7224 37128 7224 0 _0289_
rlabel metal3 40488 10584 40488 10584 0 _0290_
rlabel metal2 39368 10435 39368 10435 0 _0291_
rlabel metal2 39144 11032 39144 11032 0 _0292_
rlabel metal3 36512 10584 36512 10584 0 _0293_
rlabel metal2 39592 10248 39592 10248 0 _0294_
rlabel metal2 42840 8960 42840 8960 0 _0295_
rlabel metal2 37828 7504 37828 7504 0 _0296_
rlabel metal2 39256 5544 39256 5544 0 _0297_
rlabel metal2 37016 7616 37016 7616 0 _0298_
rlabel metal2 37688 7280 37688 7280 0 _0299_
rlabel metal2 39480 9576 39480 9576 0 _0300_
rlabel metal2 28588 16296 28588 16296 0 _0301_
rlabel metal2 30296 19208 30296 19208 0 _0302_
rlabel metal3 31724 17640 31724 17640 0 _0303_
rlabel metal2 32312 17136 32312 17136 0 _0304_
rlabel metal2 32088 18536 32088 18536 0 _0305_
rlabel metal2 31528 15764 31528 15764 0 _0306_
rlabel metal3 32928 16856 32928 16856 0 _0307_
rlabel metal2 29064 21574 29064 21574 0 _0308_
rlabel metal2 30836 22456 30836 22456 0 _0309_
rlabel metal2 31024 22232 31024 22232 0 _0310_
rlabel via2 37576 8218 37576 8218 0 _0311_
rlabel metal2 41720 5949 41720 5949 0 _0312_
rlabel metal2 34104 8568 34104 8568 0 _0313_
rlabel metal2 10808 34216 10808 34216 0 _0314_
rlabel metal2 37016 40488 37016 40488 0 _0315_
rlabel metal2 33096 36288 33096 36288 0 _0316_
rlabel metal2 34272 37240 34272 37240 0 _0317_
rlabel metal2 35336 38724 35336 38724 0 _0318_
rlabel metal3 37240 37240 37240 37240 0 _0319_
rlabel metal2 41272 36666 41272 36666 0 _0320_
rlabel metal2 33656 41552 33656 41552 0 _0321_
rlabel metal2 37464 40412 37464 40412 0 _0322_
rlabel metal2 37688 39984 37688 39984 0 _0323_
rlabel metal2 37632 41160 37632 41160 0 _0324_
rlabel metal2 36008 40412 36008 40412 0 _0325_
rlabel metal2 33451 40460 33451 40460 0 _0326_
rlabel metal2 35728 41160 35728 41160 0 _0327_
rlabel metal2 31192 41048 31192 41048 0 _0328_
rlabel metal2 33432 41320 33432 41320 0 _0329_
rlabel metal2 35896 37520 35896 37520 0 _0330_
rlabel metal2 37240 37184 37240 37184 0 _0331_
rlabel metal2 39928 37128 39928 37128 0 _0332_
rlabel metal2 40320 40096 40320 40096 0 _0333_
rlabel metal2 39816 40712 39816 40712 0 _0334_
rlabel metal2 43400 38304 43400 38304 0 _0335_
rlabel metal2 42588 38024 42588 38024 0 _0336_
rlabel metal2 31080 35616 31080 35616 0 _0337_
rlabel metal2 34776 33936 34776 33936 0 _0338_
rlabel metal2 32312 37240 32312 37240 0 _0339_
rlabel via2 41048 36442 41048 36442 0 _0340_
rlabel metal2 39816 36008 39816 36008 0 _0341_
rlabel metal2 33404 39480 33404 39480 0 _0342_
rlabel metal2 33992 35616 33992 35616 0 _0343_
rlabel metal2 34608 32732 34608 32732 0 _0344_
rlabel metal2 24752 19824 24752 19824 0 _0345_
rlabel metal3 22017 17640 22017 17640 0 _0346_
rlabel metal2 22008 19264 22008 19264 0 _0347_
rlabel via1 22241 19432 22241 19432 0 _0348_
rlabel metal3 24780 20888 24780 20888 0 _0349_
rlabel metal2 20888 20832 20888 20832 0 _0350_
rlabel metal2 24136 37520 24136 37520 0 _0351_
rlabel metal2 23352 39144 23352 39144 0 _0352_
rlabel metal2 28392 39536 28392 39536 0 _0353_
rlabel metal2 26264 37576 26264 37576 0 _0354_
rlabel metal3 26740 38024 26740 38024 0 _0355_
rlabel metal2 26376 40600 26376 40600 0 _0356_
rlabel metal2 28672 40712 28672 40712 0 _0357_
rlabel metal2 24360 39256 24360 39256 0 _0358_
rlabel metal2 24668 38920 24668 38920 0 _0359_
rlabel metal2 24808 40712 24808 40712 0 _0360_
rlabel metal2 23968 40460 23968 40460 0 _0361_
rlabel metal2 22676 39517 22676 39517 0 _0362_
rlabel metal2 22848 39116 22848 39116 0 _0363_
rlabel metal3 21896 38024 21896 38024 0 _0364_
rlabel metal2 22008 39816 22008 39816 0 _0365_
rlabel metal3 21056 38696 21056 38696 0 _0366_
rlabel metal2 22904 37576 22904 37576 0 _0367_
rlabel metal2 23968 37464 23968 37464 0 _0368_
rlabel via1 20440 36448 20440 36448 0 _0369_
rlabel metal3 22400 36456 22400 36456 0 _0370_
rlabel metal2 22456 36344 22456 36344 0 _0371_
rlabel metal2 23016 36512 23016 36512 0 _0372_
rlabel metal2 21784 35112 21784 35112 0 _0373_
rlabel metal2 22904 27272 22904 27272 0 _0374_
rlabel metal3 21756 27272 21756 27272 0 _0375_
rlabel metal2 30856 36736 30856 36736 0 _0376_
rlabel metal3 30436 36456 30436 36456 0 _0377_
rlabel metal2 34216 38220 34216 38220 0 _0378_
rlabel metal3 32564 38808 32564 38808 0 _0379_
rlabel metal3 31724 37016 31724 37016 0 _0380_
rlabel metal2 31696 38808 31696 38808 0 _0381_
rlabel metal2 32088 38752 32088 38752 0 _0382_
rlabel metal2 26824 30576 26824 30576 0 _0383_
rlabel metal2 26152 30869 26152 30869 0 _0384_
rlabel metal2 26712 29792 26712 29792 0 _0385_
rlabel metal2 27720 31976 27720 31976 0 _0386_
rlabel metal2 26264 31192 26264 31192 0 _0387_
rlabel metal2 33768 36652 33768 36652 0 _0388_
rlabel metal2 33908 36456 33908 36456 0 _0389_
rlabel metal2 26376 36344 26376 36344 0 _0390_
rlabel metal2 29064 36120 29064 36120 0 _0391_
rlabel metal2 26600 33208 26600 33208 0 _0392_
rlabel metal2 24472 33600 24472 33600 0 _0393_
rlabel metal2 27776 33544 27776 33544 0 _0394_
rlabel metal2 35784 35000 35784 35000 0 _0395_
rlabel metal2 35952 35168 35952 35168 0 _0396_
rlabel metal2 38024 32760 38024 32760 0 _0397_
rlabel metal2 28616 33404 28616 33404 0 _0398_
rlabel metal3 31640 33320 31640 33320 0 _0399_
rlabel metal2 25564 30184 25564 30184 0 _0400_
rlabel metal2 31172 31444 31172 31444 0 _0401_
rlabel metal2 31528 33368 31528 33368 0 _0402_
rlabel metal2 32424 33740 32424 33740 0 _0403_
rlabel metal2 32010 32442 32010 32442 0 _0404_
rlabel metal2 34888 31808 34888 31808 0 _0405_
rlabel metal3 35336 31808 35336 31808 0 _0406_
rlabel metal2 34636 31976 34636 31976 0 _0407_
rlabel metal2 30184 30912 30184 30912 0 _0408_
rlabel metal2 30856 30688 30856 30688 0 _0409_
rlabel metal3 34888 30968 34888 30968 0 _0410_
rlabel metal2 34552 30800 34552 30800 0 _0411_
rlabel metal2 34440 31668 34440 31668 0 _0412_
rlabel metal2 35980 31640 35980 31640 0 _0413_
rlabel metal2 34776 32900 34776 32900 0 _0414_
rlabel metal3 34804 32648 34804 32648 0 _0415_
rlabel metal2 30352 31304 30352 31304 0 _0416_
rlabel metal3 31752 31752 31752 31752 0 _0417_
rlabel metal2 33432 31808 33432 31808 0 _0418_
rlabel metal3 32368 30184 32368 30184 0 _0419_
rlabel metal3 30324 24808 30324 24808 0 _0420_
rlabel metal3 33152 30408 33152 30408 0 _0421_
rlabel metal2 33208 30072 33208 30072 0 _0422_
rlabel metal2 31080 29092 31080 29092 0 _0423_
rlabel metal2 32424 29568 32424 29568 0 _0424_
rlabel metal3 33628 30968 33628 30968 0 _0425_
rlabel metal2 33880 33058 33880 33058 0 _0426_
rlabel via2 33544 34120 33544 34120 0 _0427_
rlabel metal3 33964 35672 33964 35672 0 _0428_
rlabel metal2 32536 35308 32536 35308 0 _0429_
rlabel metal2 40040 31654 40040 31654 0 _0430_
rlabel metal2 39816 32844 39816 32844 0 _0431_
rlabel metal2 39564 32648 39564 32648 0 _0432_
rlabel metal2 24696 16688 24696 16688 0 _0433_
rlabel metal2 25144 18368 25144 18368 0 _0434_
rlabel metal2 23623 16856 23623 16856 0 _0435_
rlabel metal2 29064 13160 29064 13160 0 _0436_
rlabel metal2 43176 13832 43176 13832 0 _0437_
rlabel metal3 29904 15288 29904 15288 0 _0438_
rlabel metal2 25144 26544 25144 26544 0 _0439_
rlabel metal2 17752 30632 17752 30632 0 _0440_
rlabel metal2 15176 35560 15176 35560 0 _0441_
rlabel metal2 19544 25508 19544 25508 0 _0442_
rlabel metal3 17556 33544 17556 33544 0 _0443_
rlabel metal2 17556 33544 17556 33544 0 _0444_
rlabel metal2 15064 32032 15064 32032 0 _0445_
rlabel metal2 13944 30352 13944 30352 0 _0446_
rlabel metal2 16968 27832 16968 27832 0 _0447_
rlabel metal2 17500 31080 17500 31080 0 _0448_
rlabel metal2 18116 29512 18116 29512 0 _0449_
rlabel metal2 41496 15680 41496 15680 0 _0450_
rlabel via1 38239 15960 38239 15960 0 _0451_
rlabel metal2 42410 14056 42410 14056 0 _0452_
rlabel metal3 42905 15064 42905 15064 0 _0453_
rlabel metal3 41711 13720 41711 13720 0 _0454_
rlabel metal2 40096 17080 40096 17080 0 _0455_
rlabel metal2 16520 19488 16520 19488 0 _0456_
rlabel metal2 34160 12936 34160 12936 0 _0457_
rlabel metal2 32070 13440 32070 13440 0 _0458_
rlabel metal2 42840 17976 42840 17976 0 _0459_
rlabel metal3 20300 20552 20300 20552 0 _0460_
rlabel metal2 36120 12320 36120 12320 0 _0461_
rlabel metal2 42616 19656 42616 19656 0 _0462_
rlabel metal2 18928 18200 18928 18200 0 _0463_
rlabel metal2 35224 15204 35224 15204 0 _0464_
rlabel metal2 39144 14056 39144 14056 0 _0465_
rlabel metal2 19768 32648 19768 32648 0 _0466_
rlabel metal2 35000 17696 35000 17696 0 _0467_
rlabel metal2 33190 20160 33190 20160 0 _0468_
rlabel metal2 34534 20384 34534 20384 0 _0469_
rlabel metal2 34151 17864 34151 17864 0 _0470_
rlabel metal2 19208 20440 19208 20440 0 _0471_
rlabel metal3 17033 19992 17033 19992 0 _0472_
rlabel via1 18303 21000 18303 21000 0 _0473_
rlabel metal2 17239 18424 17239 18424 0 _0474_
rlabel metal3 18368 16856 18368 16856 0 _0475_
rlabel metal2 17239 16856 17239 16856 0 _0476_
rlabel metal3 17472 15288 17472 15288 0 _0477_
rlabel via1 15745 15064 15745 15064 0 _0478_
rlabel metal2 15783 13720 15783 13720 0 _0479_
rlabel metal2 17239 15288 17239 15288 0 _0480_
rlabel metal2 19302 14784 19302 14784 0 _0481_
rlabel metal2 27384 12880 27384 12880 0 _0482_
rlabel metal2 34328 3752 34328 3752 0 _0483_
rlabel metal2 26040 8176 26040 8176 0 _0484_
rlabel metal2 36456 4200 36456 4200 0 _0485_
rlabel metal2 26264 7504 26264 7504 0 _0486_
rlabel metal2 35952 5096 35952 5096 0 _0487_
rlabel metal2 25312 17752 25312 17752 0 _0488_
rlabel metal2 27832 12488 27832 12488 0 _0489_
rlabel metal2 24808 11256 24808 11256 0 _0490_
rlabel metal2 28168 10920 28168 10920 0 _0491_
rlabel metal2 24192 13720 24192 13720 0 _0492_
rlabel metal3 25116 15512 25116 15512 0 _0493_
rlabel metal3 28849 3752 28849 3752 0 _0494_
rlabel metal2 23296 5880 23296 5880 0 _0495_
rlabel metal2 26824 6104 26824 6104 0 _0496_
rlabel metal2 22727 15288 22727 15288 0 _0497_
rlabel metal3 30576 7560 30576 7560 0 _0498_
rlabel metal2 30538 4648 30538 4648 0 _0499_
rlabel metal2 30585 6664 30585 6664 0 _0500_
rlabel metal2 29158 7728 29158 7728 0 _0501_
rlabel metal2 38808 20636 38808 20636 0 _0502_
rlabel metal2 36633 17640 36633 17640 0 _0503_
rlabel metal2 38089 19208 38089 19208 0 _0504_
rlabel via1 39377 20888 39377 20888 0 _0505_
rlabel metal2 39928 20328 39928 20328 0 _0506_
rlabel metal2 43176 18284 43176 18284 0 _0507_
rlabel metal3 40311 19432 40311 19432 0 _0508_
rlabel metal2 42616 17192 42616 17192 0 _0509_
rlabel via1 41487 16968 41487 16968 0 _0510_
rlabel metal2 42775 20776 42775 20776 0 _0511_
rlabel metal3 30240 20104 30240 20104 0 _0512_
rlabel metal2 28392 19908 28392 19908 0 _0513_
rlabel metal2 26656 26488 26656 26488 0 _0514_
rlabel metal2 26376 22098 26376 22098 0 _0515_
rlabel metal2 27048 25396 27048 25396 0 _0516_
rlabel via2 26824 28608 26824 28608 0 _0517_
rlabel metal3 28056 27272 28056 27272 0 _0518_
rlabel metal2 27496 25396 27496 25396 0 _0519_
rlabel metal2 25928 25284 25928 25284 0 _0520_
rlabel metal2 26152 25368 26152 25368 0 _0521_
rlabel metal2 24808 24976 24808 24976 0 _0522_
rlabel metal2 26376 25275 26376 25275 0 _0523_
rlabel metal2 26544 26264 26544 26264 0 _0524_
rlabel metal2 26264 27524 26264 27524 0 _0525_
rlabel metal2 27048 25592 27048 25592 0 _0526_
rlabel metal2 26600 27972 26600 27972 0 _0527_
rlabel metal2 25648 28616 25648 28616 0 _0528_
rlabel metal3 41090 2744 41090 2744 0 clk
rlabel metal3 24136 22568 24136 22568 0 clknet_0__0209_
rlabel metal3 25256 24472 25256 24472 0 clknet_0__0210_
rlabel metal3 36008 25368 36008 25368 0 clknet_0__0228_
rlabel metal2 41272 26781 41272 26781 0 clknet_0__0229_
rlabel metal3 41328 24920 41328 24920 0 clknet_0__0230_
rlabel metal2 39816 25354 39816 25354 0 clknet_0__0231_
rlabel metal2 21448 11984 21448 11984 0 clknet_0__0254_
rlabel metal2 17976 9898 17976 9898 0 clknet_0__0255_
rlabel metal3 23576 3528 23576 3528 0 clknet_0__0256_
rlabel metal2 21672 8988 21672 8988 0 clknet_0__0257_
rlabel metal2 15176 22610 15176 22610 0 clknet_0__0282_
rlabel metal2 9128 18634 9128 18634 0 clknet_0__0283_
rlabel metal3 12152 15512 12152 15512 0 clknet_0__0284_
rlabel metal2 13328 20216 13328 20216 0 clknet_0__0285_
rlabel metal3 36232 12152 36232 12152 0 clknet_0__0310_
rlabel metal3 40376 8232 40376 8232 0 clknet_0__0311_
rlabel metal2 40264 5837 40264 5837 0 clknet_0__0312_
rlabel metal2 40376 8722 40376 8722 0 clknet_0__0313_
rlabel metal2 28280 34173 28280 34173 0 clknet_0_clk
rlabel metal2 22288 22344 22288 22344 0 clknet_1_0__leaf__0209_
rlabel metal2 21224 23436 21224 23436 0 clknet_1_0__leaf__0210_
rlabel metal3 31808 23128 31808 23128 0 clknet_1_0__leaf__0228_
rlabel metal2 32200 26594 32200 26594 0 clknet_1_0__leaf__0229_
rlabel metal2 41272 29351 41272 29351 0 clknet_1_0__leaf__0230_
rlabel metal2 33768 28134 33768 28134 0 clknet_1_0__leaf__0231_
rlabel metal2 18984 9912 18984 9912 0 clknet_1_0__leaf__0254_
rlabel metal2 17528 5439 17528 5439 0 clknet_1_0__leaf__0255_
rlabel metal2 22568 4039 22568 4039 0 clknet_1_0__leaf__0256_
rlabel metal2 18536 7175 18536 7175 0 clknet_1_0__leaf__0257_
rlabel metal2 8512 21560 8512 21560 0 clknet_1_0__leaf__0282_
rlabel metal2 9072 14504 9072 14504 0 clknet_1_0__leaf__0283_
rlabel via2 8120 13727 8120 13727 0 clknet_1_0__leaf__0284_
rlabel via2 10248 18431 10248 18431 0 clknet_1_0__leaf__0285_
rlabel metal3 31472 9016 31472 9016 0 clknet_1_0__leaf__0310_
rlabel metal2 39816 10808 39816 10808 0 clknet_1_0__leaf__0311_
rlabel metal2 39368 5824 39368 5824 0 clknet_1_0__leaf__0312_
rlabel metal2 34944 10668 34944 10668 0 clknet_1_0__leaf__0313_
rlabel metal2 26488 21504 26488 21504 0 clknet_1_1__leaf__0209_
rlabel metal2 28728 23968 28728 23968 0 clknet_1_1__leaf__0210_
rlabel metal3 37296 25480 37296 25480 0 clknet_1_1__leaf__0228_
rlabel metal3 40936 27048 40936 27048 0 clknet_1_1__leaf__0229_
rlabel metal2 43512 23430 43512 23430 0 clknet_1_1__leaf__0230_
rlabel metal3 36736 25256 36736 25256 0 clknet_1_1__leaf__0231_
rlabel metal2 20328 13608 20328 13608 0 clknet_1_1__leaf__0254_
rlabel metal2 17024 9912 17024 9912 0 clknet_1_1__leaf__0255_
rlabel metal2 18536 5958 18536 5958 0 clknet_1_1__leaf__0256_
rlabel via1 18760 12159 18760 12159 0 clknet_1_1__leaf__0257_
rlabel metal2 16184 22848 16184 22848 0 clknet_1_1__leaf__0282_
rlabel metal3 9128 19432 9128 19432 0 clknet_1_1__leaf__0283_
rlabel metal3 8904 16464 8904 16464 0 clknet_1_1__leaf__0284_
rlabel metal2 9912 23206 9912 23206 0 clknet_1_1__leaf__0285_
rlabel metal2 39032 10024 39032 10024 0 clknet_1_1__leaf__0310_
rlabel via2 43848 7455 43848 7455 0 clknet_1_1__leaf__0311_
rlabel via1 43344 5081 43344 5081 0 clknet_1_1__leaf__0312_
rlabel metal2 36120 7750 36120 7750 0 clknet_1_1__leaf__0313_
rlabel metal2 28672 39760 28672 39760 0 clknet_2_0__leaf_clk
rlabel via2 20776 39592 20776 39592 0 clknet_2_1__leaf_clk
rlabel metal2 38920 33600 38920 33600 0 clknet_2_2__leaf_clk
rlabel metal3 35280 38808 35280 38808 0 clknet_2_3__leaf_clk
rlabel metal2 44296 9632 44296 9632 0 io_in[0]
rlabel metal2 44352 11368 44352 11368 0 io_in[1]
rlabel metal3 44758 16184 44758 16184 0 io_in[2]
rlabel metal3 42812 19992 42812 19992 0 io_in[3]
rlabel metal2 43064 21392 43064 21392 0 io_in[4]
rlabel metal2 44324 28392 44324 28392 0 io_in[5]
rlabel metal3 44338 29624 44338 29624 0 io_out[0]
rlabel metal2 43176 32704 43176 32704 0 io_out[1]
rlabel metal2 43176 36456 43176 36456 0 io_out[2]
rlabel metal2 43400 40320 43400 40320 0 io_out[3]
rlabel metal2 41720 42616 41720 42616 0 io_out[4]
rlabel metal3 31276 15400 31276 15400 0 net1
rlabel metal2 43064 40893 43064 40893 0 net10
rlabel metal2 21224 32144 21224 32144 0 net11
rlabel metal3 8904 33320 8904 33320 0 net12
rlabel metal2 13048 34496 13048 34496 0 net13
rlabel metal2 11872 36232 11872 36232 0 net14
rlabel metal2 13496 29288 13496 29288 0 net15
rlabel metal2 14784 31080 14784 31080 0 net16
rlabel metal2 13160 34664 13160 34664 0 net17
rlabel metal2 12936 34944 12936 34944 0 net18
rlabel metal2 14056 27272 14056 27272 0 net19
rlabel metal3 37856 11592 37856 11592 0 net2
rlabel metal2 20496 26600 20496 26600 0 net20
rlabel metal3 20944 26824 20944 26824 0 net21
rlabel metal3 15848 14504 15848 14504 0 net22
rlabel metal3 18704 14616 18704 14616 0 net23
rlabel metal2 21896 12936 21896 12936 0 net24
rlabel metal2 26040 4592 26040 4592 0 net25
rlabel metal2 26488 14840 26488 14840 0 net26
rlabel metal3 23968 15288 23968 15288 0 net27
rlabel metal2 15848 16856 15848 16856 0 net28
rlabel metal2 18984 19992 18984 19992 0 net29
rlabel metal2 43036 29960 43036 29960 0 net3
rlabel metal2 18424 21672 18424 21672 0 net30
rlabel metal2 23800 27720 23800 27720 0 net31
rlabel metal2 24864 21140 24864 21140 0 net32
rlabel metal2 24584 22848 24584 22848 0 net33
rlabel metal3 23968 19656 23968 19656 0 net34
rlabel metal2 31976 8176 31976 8176 0 net35
rlabel metal2 29176 8960 29176 8960 0 net36
rlabel metal2 40600 13720 40600 13720 0 net37
rlabel metal2 37128 15792 37128 15792 0 net38
rlabel metal2 36120 13832 36120 13832 0 net39
rlabel metal3 25340 19992 25340 19992 0 net4
rlabel metal3 33040 20776 33040 20776 0 net40
rlabel metal2 40936 19712 40936 19712 0 net41
rlabel metal3 40320 18424 40320 18424 0 net42
rlabel metal2 40152 19152 40152 19152 0 net43
rlabel metal2 31976 22232 31976 22232 0 net44
rlabel metal3 30744 20776 30744 20776 0 net45
rlabel metal2 24248 25172 24248 25172 0 net46
rlabel metal2 21224 25592 21224 25592 0 net47
rlabel via3 31388 20552 31388 20552 0 net5
rlabel metal2 41944 30085 41944 30085 0 net6
rlabel metal2 43848 32829 43848 32829 0 net7
rlabel metal2 43848 36162 43848 36162 0 net8
rlabel metal2 42840 37072 42840 37072 0 net9
rlabel metal2 44296 5264 44296 5264 0 rst_n
rlabel metal2 27272 39536 27272 39536 0 slow_clock\[0\]
rlabel metal2 27720 39116 27720 39116 0 slow_clock\[1\]
rlabel metal2 28000 40376 28000 40376 0 slow_clock\[2\]
rlabel metal2 23632 40376 23632 40376 0 slow_clock\[3\]
rlabel metal2 22456 39312 22456 39312 0 slow_clock\[4\]
rlabel metal3 22904 37240 22904 37240 0 slow_clock\[5\]
rlabel metal2 21504 36456 21504 36456 0 slow_clock\[6\]
rlabel metal3 37016 38024 37016 38024 0 spi_dac_i_2.counter\[0\]
rlabel metal2 38360 41048 38360 41048 0 spi_dac_i_2.counter\[1\]
rlabel via2 37128 41160 37128 41160 0 spi_dac_i_2.counter\[2\]
rlabel metal2 32424 41216 32424 41216 0 spi_dac_i_2.counter\[3\]
rlabel metal3 34160 39592 34160 39592 0 spi_dac_i_2.counter\[4\]
rlabel metal2 43512 33656 43512 33656 0 spi_dac_i_2.spi_clk
rlabel metal3 43512 35616 43512 35616 0 spi_dac_i_2.spi_dat
rlabel metal2 31640 37352 31640 37352 0 spi_dac_i_2.spi_dat_buff\[0\]
rlabel metal2 34160 35532 34160 35532 0 spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal3 41496 34776 41496 34776 0 spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 33656 38920 33656 38920 0 spi_dac_i_2.spi_dat_buff\[1\]
rlabel metal2 41384 40628 41384 40628 0 spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 40824 40852 40824 40852 0 spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal3 41328 38696 41328 38696 0 spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 42168 37716 42168 37716 0 spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal2 32984 36288 32984 36288 0 spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal3 37240 35000 37240 35000 0 spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 37912 32172 37912 32172 0 spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal2 37352 33586 37352 33586 0 spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal2 42280 33208 42280 33208 0 spi_dac_i_2.spi_le
<< properties >>
string FIXED_BBOX 0 0 46000 46000
<< end >>
